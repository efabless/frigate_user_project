magic
tech sky130A
magscale 1 2
timestamp 1740504979
<< viali >>
rect 2513 37281 2547 37315
rect 13553 37281 13587 37315
rect 34069 37281 34103 37315
rect 39589 37281 39623 37315
rect 3525 37213 3559 37247
rect 5917 37213 5951 37247
rect 7021 37213 7055 37247
rect 7849 37213 7883 37247
rect 8769 37213 8803 37247
rect 11345 37213 11379 37247
rect 12081 37213 12115 37247
rect 14565 37213 14599 37247
rect 15209 37213 15243 37247
rect 18705 37213 18739 37247
rect 19533 37213 19567 37247
rect 20913 37213 20947 37247
rect 21925 37213 21959 37247
rect 22753 37213 22787 37247
rect 26249 37213 26283 37247
rect 28273 37213 28307 37247
rect 29285 37213 29319 37247
rect 31769 37213 31803 37247
rect 32781 37213 32815 37247
rect 33793 37213 33827 37247
rect 36829 37213 36863 37247
rect 37565 37213 37599 37247
rect 39129 37213 39163 37247
rect 40969 37213 41003 37247
rect 41889 37213 41923 37247
rect 43361 37213 43395 37247
rect 46489 37213 46523 37247
rect 48513 37213 48547 37247
rect 52009 37213 52043 37247
rect 52929 37213 52963 37247
rect 53849 37213 53883 37247
rect 56241 37213 56275 37247
rect 58817 37213 58851 37247
rect 16129 37145 16163 37179
rect 23673 37145 23707 37179
rect 27169 37145 27203 37179
rect 44281 37145 44315 37179
rect 47409 37145 47443 37179
rect 49433 37145 49467 37179
rect 54769 37145 54803 37179
rect 57161 37145 57195 37179
rect 59737 37145 59771 37179
rect 7757 36873 7791 36907
rect 11897 36873 11931 36907
rect 15117 36873 15151 36907
rect 19073 36873 19107 36907
rect 22477 36873 22511 36907
rect 26157 36873 26191 36907
rect 33793 36873 33827 36907
rect 37013 36873 37047 36907
rect 40877 36873 40911 36907
rect 48237 36873 48271 36907
rect 51917 36873 51951 36907
rect 55597 36873 55631 36907
rect 4353 36805 4387 36839
rect 9873 36805 9907 36839
rect 17969 36805 18003 36839
rect 24593 36805 24627 36839
rect 5457 36737 5491 36771
rect 7573 36737 7607 36771
rect 10885 36737 10919 36771
rect 11805 36737 11839 36771
rect 12081 36737 12115 36771
rect 14933 36737 14967 36771
rect 18981 36737 19015 36771
rect 19257 36737 19291 36771
rect 22293 36737 22327 36771
rect 25789 36737 25823 36771
rect 25973 36737 26007 36771
rect 29653 36737 29687 36771
rect 29929 36737 29963 36771
rect 33517 36737 33551 36771
rect 33701 36737 33735 36771
rect 33977 36737 34011 36771
rect 35449 36737 35483 36771
rect 37197 36737 37231 36771
rect 40693 36737 40727 36771
rect 44373 36737 44407 36771
rect 44649 36737 44683 36771
rect 48053 36737 48087 36771
rect 50169 36737 50203 36771
rect 51733 36737 51767 36771
rect 55413 36737 55447 36771
rect 58449 36737 58483 36771
rect 59369 36737 59403 36771
rect 11621 36669 11655 36703
rect 30389 36669 30423 36703
rect 35909 36669 35943 36703
rect 45109 36669 45143 36703
rect 50629 36669 50663 36703
rect 59829 36669 59863 36703
rect 29837 36601 29871 36635
rect 44557 36601 44591 36635
rect 58633 36601 58667 36635
rect 28733 11781 28767 11815
rect 29101 11713 29135 11747
rect 29469 11713 29503 11747
rect 29653 11713 29687 11747
rect 29745 11713 29779 11747
rect 28549 11509 28583 11543
rect 29285 11509 29319 11543
rect 24225 11305 24259 11339
rect 28457 11305 28491 11339
rect 28825 11305 28859 11339
rect 22109 11237 22143 11271
rect 22293 11237 22327 11271
rect 22753 11237 22787 11271
rect 23489 11237 23523 11271
rect 27997 11237 28031 11271
rect 28319 11237 28353 11271
rect 23857 11169 23891 11203
rect 25421 11169 25455 11203
rect 25605 11169 25639 11203
rect 28549 11169 28583 11203
rect 29653 11169 29687 11203
rect 21925 11101 21959 11135
rect 22017 11101 22051 11135
rect 22477 11101 22511 11135
rect 23673 11101 23707 11135
rect 23949 11101 23983 11135
rect 24133 11101 24167 11135
rect 24409 11101 24443 11135
rect 24593 11101 24627 11135
rect 24685 11101 24719 11135
rect 24777 11101 24811 11135
rect 24961 11101 24995 11135
rect 25513 11101 25547 11135
rect 25697 11101 25731 11135
rect 26065 11101 26099 11135
rect 26249 11101 26283 11135
rect 26341 11101 26375 11135
rect 26525 11101 26559 11135
rect 26617 11101 26651 11135
rect 27077 11101 27111 11135
rect 27261 11101 27295 11135
rect 27353 11101 27387 11135
rect 28181 11101 28215 11135
rect 29372 11101 29406 11135
rect 29837 11101 29871 11135
rect 22201 11033 22235 11067
rect 22937 11033 22971 11067
rect 24869 11033 24903 11067
rect 29469 11033 29503 11067
rect 25881 10965 25915 10999
rect 21925 10761 21959 10795
rect 22201 10761 22235 10795
rect 27905 10761 27939 10795
rect 28917 10761 28951 10795
rect 30941 10761 30975 10795
rect 23397 10693 23431 10727
rect 31217 10693 31251 10727
rect 35081 10693 35115 10727
rect 20453 10625 20487 10659
rect 20729 10625 20763 10659
rect 21281 10625 21315 10659
rect 21741 10625 21775 10659
rect 22017 10625 22051 10659
rect 22109 10625 22143 10659
rect 22385 10625 22419 10659
rect 22937 10625 22971 10659
rect 23581 10625 23615 10659
rect 27353 10625 27387 10659
rect 27721 10625 27755 10659
rect 28825 10625 28859 10659
rect 30757 10625 30791 10659
rect 31033 10625 31067 10659
rect 33517 10625 33551 10659
rect 34897 10625 34931 10659
rect 35173 10625 35207 10659
rect 35265 10625 35299 10659
rect 24133 10557 24167 10591
rect 25053 10557 25087 10591
rect 25329 10557 25363 10591
rect 26249 10557 26283 10591
rect 26801 10557 26835 10591
rect 28457 10557 28491 10591
rect 29469 10557 29503 10591
rect 29653 10557 29687 10591
rect 33241 10557 33275 10591
rect 33333 10557 33367 10591
rect 33425 10557 33459 10591
rect 33701 10557 33735 10591
rect 20729 10489 20763 10523
rect 30573 10489 30607 10523
rect 21373 10421 21407 10455
rect 21557 10421 21591 10455
rect 22569 10421 22603 10455
rect 22753 10421 22787 10455
rect 23121 10421 23155 10455
rect 24501 10421 24535 10455
rect 25973 10421 26007 10455
rect 26065 10421 26099 10455
rect 27537 10421 27571 10455
rect 28641 10421 28675 10455
rect 30205 10421 30239 10455
rect 31493 10421 31527 10455
rect 33057 10421 33091 10455
rect 34253 10421 34287 10455
rect 35449 10421 35483 10455
rect 19809 10217 19843 10251
rect 19993 10217 20027 10251
rect 27537 10217 27571 10251
rect 28549 10217 28583 10251
rect 27629 10149 27663 10183
rect 21005 10081 21039 10115
rect 22661 10081 22695 10115
rect 25973 10081 26007 10115
rect 26709 10081 26743 10115
rect 27905 10081 27939 10115
rect 31125 10081 31159 10115
rect 31217 10081 31251 10115
rect 31953 10081 31987 10115
rect 33517 10081 33551 10115
rect 34805 10081 34839 10115
rect 19625 10013 19659 10047
rect 19717 10013 19751 10047
rect 20729 10013 20763 10047
rect 20913 10013 20947 10047
rect 21925 10013 21959 10047
rect 23489 10013 23523 10047
rect 24133 10013 24167 10047
rect 24593 10013 24627 10047
rect 25513 10013 25547 10047
rect 25697 10013 25731 10047
rect 26893 10013 26927 10047
rect 27813 10013 27847 10047
rect 29653 10013 29687 10047
rect 31861 10013 31895 10047
rect 32689 10013 32723 10047
rect 34069 10013 34103 10047
rect 35633 10013 35667 10047
rect 36737 10013 36771 10047
rect 22845 9945 22879 9979
rect 25881 9945 25915 9979
rect 34253 9945 34287 9979
rect 20545 9877 20579 9911
rect 21373 9877 21407 9911
rect 22109 9877 22143 9911
rect 23581 9877 23615 9911
rect 25145 9877 25179 9911
rect 25329 9877 25363 9911
rect 25605 9877 25639 9911
rect 26157 9877 26191 9911
rect 28641 9877 28675 9911
rect 29009 9877 29043 9911
rect 30297 9877 30331 9911
rect 30481 9877 30515 9911
rect 32597 9877 32631 9911
rect 33333 9877 33367 9911
rect 36277 9877 36311 9911
rect 37289 9877 37323 9911
rect 24133 9673 24167 9707
rect 28825 9673 28859 9707
rect 33241 9673 33275 9707
rect 21741 9605 21775 9639
rect 22569 9605 22603 9639
rect 24393 9605 24427 9639
rect 24593 9605 24627 9639
rect 26617 9605 26651 9639
rect 27905 9605 27939 9639
rect 32873 9605 32907 9639
rect 34437 9605 34471 9639
rect 18705 9537 18739 9571
rect 19165 9537 19199 9571
rect 19257 9537 19291 9571
rect 19435 9537 19469 9571
rect 19533 9537 19567 9571
rect 19717 9537 19751 9571
rect 22017 9537 22051 9571
rect 22753 9537 22787 9571
rect 22845 9537 22879 9571
rect 23029 9537 23063 9571
rect 25421 9537 25455 9571
rect 25973 9537 26007 9571
rect 28089 9537 28123 9571
rect 29561 9537 29595 9571
rect 29745 9537 29779 9571
rect 33057 9537 33091 9571
rect 33333 9537 33367 9571
rect 33425 9537 33459 9571
rect 35909 9537 35943 9571
rect 38761 9537 38795 9571
rect 19625 9469 19659 9503
rect 19809 9469 19843 9503
rect 20453 9469 20487 9503
rect 20545 9469 20579 9503
rect 21373 9469 21407 9503
rect 23489 9469 23523 9503
rect 25329 9469 25363 9503
rect 27169 9469 27203 9503
rect 29377 9469 29411 9503
rect 30021 9469 30055 9503
rect 30665 9469 30699 9503
rect 31309 9469 31343 9503
rect 32045 9469 32079 9503
rect 32229 9469 32263 9503
rect 33701 9469 33735 9503
rect 34253 9469 34287 9503
rect 34989 9469 35023 9503
rect 36553 9469 36587 9503
rect 37381 9469 37415 9503
rect 18889 9401 18923 9435
rect 21189 9401 21223 9435
rect 24225 9401 24259 9435
rect 24685 9401 24719 9435
rect 31493 9401 31527 9435
rect 36001 9401 36035 9435
rect 18981 9333 19015 9367
rect 19441 9333 19475 9367
rect 21649 9333 21683 9367
rect 23213 9333 23247 9367
rect 23305 9333 23339 9367
rect 24409 9333 24443 9367
rect 28733 9333 28767 9367
rect 29929 9333 29963 9367
rect 30757 9333 30791 9367
rect 33609 9333 33643 9367
rect 35265 9333 35299 9367
rect 36737 9333 36771 9367
rect 38209 9333 38243 9367
rect 11805 9129 11839 9163
rect 17233 9129 17267 9163
rect 17601 9129 17635 9163
rect 27813 9129 27847 9163
rect 28641 9129 28675 9163
rect 34345 9129 34379 9163
rect 31033 9061 31067 9095
rect 17325 8993 17359 9027
rect 19349 8993 19383 9027
rect 21005 8993 21039 9027
rect 22477 8993 22511 9027
rect 23581 8993 23615 9027
rect 26249 8993 26283 9027
rect 26985 8993 27019 9027
rect 28825 8993 28859 9027
rect 29377 8993 29411 9027
rect 31217 8993 31251 9027
rect 31585 8993 31619 9027
rect 32505 8993 32539 9027
rect 36185 8993 36219 9027
rect 38025 8993 38059 9027
rect 11897 8925 11931 8959
rect 17233 8925 17267 8959
rect 19165 8925 19199 8959
rect 19901 8925 19935 8959
rect 20177 8925 20211 8959
rect 20361 8925 20395 8959
rect 21741 8925 21775 8959
rect 24317 8925 24351 8959
rect 24501 8925 24535 8959
rect 25329 8925 25363 8959
rect 26341 8925 26375 8959
rect 27721 8925 27755 8959
rect 27997 8925 28031 8959
rect 29653 8925 29687 8959
rect 31309 8925 31343 8959
rect 32413 8925 32447 8959
rect 33149 8925 33183 8959
rect 33977 8925 34011 8959
rect 34897 8925 34931 8959
rect 36369 8925 36403 8959
rect 36921 8925 36955 8959
rect 38117 8925 38151 8959
rect 18061 8857 18095 8891
rect 20453 8857 20487 8891
rect 23029 8857 23063 8891
rect 25605 8857 25639 8891
rect 28089 8857 28123 8891
rect 28365 8857 28399 8891
rect 30849 8857 30883 8891
rect 31677 8857 31711 8891
rect 37381 8857 37415 8891
rect 18613 8789 18647 8823
rect 20269 8789 20303 8823
rect 21189 8789 21223 8823
rect 21925 8789 21959 8823
rect 23765 8789 23799 8823
rect 25145 8789 25179 8823
rect 27077 8789 27111 8823
rect 28273 8789 28307 8823
rect 28457 8789 28491 8823
rect 30297 8789 30331 8823
rect 31769 8789 31803 8823
rect 33333 8789 33367 8823
rect 34989 8789 35023 8823
rect 35633 8789 35667 8823
rect 38669 8789 38703 8823
rect 19257 8585 19291 8619
rect 23029 8585 23063 8619
rect 33241 8585 33275 8619
rect 33977 8585 34011 8619
rect 19717 8517 19751 8551
rect 26341 8517 26375 8551
rect 28917 8517 28951 8551
rect 31677 8517 31711 8551
rect 32873 8517 32907 8551
rect 35081 8517 35115 8551
rect 16037 8449 16071 8483
rect 17877 8449 17911 8483
rect 27077 8449 27111 8483
rect 27905 8449 27939 8483
rect 28089 8449 28123 8483
rect 31769 8449 31803 8483
rect 33057 8449 33091 8483
rect 33241 8449 33275 8483
rect 33517 8449 33551 8483
rect 33609 8449 33643 8483
rect 33793 8449 33827 8483
rect 36921 8449 36955 8483
rect 16773 8381 16807 8415
rect 18613 8381 18647 8415
rect 20269 8381 20303 8415
rect 20453 8381 20487 8415
rect 21741 8381 21775 8415
rect 21925 8381 21959 8415
rect 23581 8381 23615 8415
rect 24041 8381 24075 8415
rect 24317 8381 24351 8415
rect 26065 8381 26099 8415
rect 26985 8381 27019 8415
rect 28181 8381 28215 8415
rect 28825 8381 28859 8415
rect 29469 8381 29503 8415
rect 29653 8381 29687 8415
rect 29929 8381 29963 8415
rect 32229 8381 32263 8415
rect 34621 8381 34655 8415
rect 34805 8381 34839 8415
rect 36829 8381 36863 8415
rect 38761 8381 38795 8415
rect 39313 8381 39347 8415
rect 39957 8381 39991 8415
rect 40233 8381 40267 8415
rect 15485 8313 15519 8347
rect 17325 8313 17359 8347
rect 18521 8313 18555 8347
rect 19441 8313 19475 8347
rect 21097 8313 21131 8347
rect 21189 8313 21223 8347
rect 27721 8313 27755 8347
rect 27905 8313 27939 8347
rect 33701 8313 33735 8347
rect 38209 8313 38243 8347
rect 40877 8313 40911 8347
rect 22569 8245 22603 8279
rect 31953 8245 31987 8279
rect 34069 8245 34103 8279
rect 37565 8245 37599 8279
rect 16681 8041 16715 8075
rect 18153 8041 18187 8075
rect 19625 8041 19659 8075
rect 21097 8041 21131 8075
rect 26341 8041 26375 8075
rect 27077 8041 27111 8075
rect 30297 8041 30331 8075
rect 30481 8041 30515 8075
rect 34713 8041 34747 8075
rect 35633 8041 35667 8075
rect 37761 8041 37795 8075
rect 24409 7973 24443 8007
rect 28089 7973 28123 8007
rect 29561 7973 29595 8007
rect 31769 7973 31803 8007
rect 17509 7905 17543 7939
rect 18981 7905 19015 7939
rect 21741 7905 21775 7939
rect 22109 7905 22143 7939
rect 24133 7905 24167 7939
rect 26249 7905 26283 7939
rect 28825 7905 28859 7939
rect 28917 7905 28951 7939
rect 33885 7905 33919 7939
rect 34161 7905 34195 7939
rect 38669 7905 38703 7939
rect 40049 7905 40083 7939
rect 14841 7837 14875 7871
rect 15393 7837 15427 7871
rect 16313 7837 16347 7871
rect 17233 7837 17267 7871
rect 18797 7837 18831 7871
rect 20453 7837 20487 7871
rect 20637 7837 20671 7871
rect 20729 7837 20763 7871
rect 20821 7837 20855 7871
rect 21189 7837 21223 7871
rect 24225 7837 24259 7871
rect 24409 7837 24443 7871
rect 25053 7837 25087 7871
rect 26985 7837 27019 7871
rect 27629 7837 27663 7871
rect 27813 7837 27847 7871
rect 28089 7837 28123 7871
rect 29653 7837 29687 7871
rect 30665 7837 30699 7871
rect 30849 7837 30883 7871
rect 30941 7837 30975 7871
rect 31585 7837 31619 7871
rect 31769 7837 31803 7871
rect 31861 7837 31895 7871
rect 34253 7837 34287 7871
rect 34529 7837 34563 7871
rect 34805 7837 34839 7871
rect 35633 7837 35667 7871
rect 35817 7837 35851 7871
rect 38025 7837 38059 7871
rect 40325 7837 40359 7871
rect 40601 7837 40635 7871
rect 22385 7769 22419 7803
rect 24501 7769 24535 7803
rect 31033 7769 31067 7803
rect 32045 7769 32079 7803
rect 32137 7769 32171 7803
rect 36001 7769 36035 7803
rect 14657 7701 14691 7735
rect 15761 7701 15795 7735
rect 18245 7701 18279 7735
rect 19809 7701 19843 7735
rect 25605 7701 25639 7735
rect 27905 7701 27939 7735
rect 28181 7701 28215 7735
rect 34345 7701 34379 7735
rect 35449 7701 35483 7735
rect 38117 7701 38151 7735
rect 39405 7701 39439 7735
rect 40141 7701 40175 7735
rect 40509 7701 40543 7735
rect 17601 7497 17635 7531
rect 20361 7497 20395 7531
rect 23397 7497 23431 7531
rect 29561 7497 29595 7531
rect 32229 7497 32263 7531
rect 33977 7497 34011 7531
rect 34713 7497 34747 7531
rect 25329 7429 25363 7463
rect 27353 7429 27387 7463
rect 27445 7429 27479 7463
rect 27537 7429 27571 7463
rect 32137 7429 32171 7463
rect 12725 7361 12759 7395
rect 14289 7361 14323 7395
rect 15393 7361 15427 7395
rect 17785 7361 17819 7395
rect 17877 7361 17911 7395
rect 18153 7361 18187 7395
rect 18981 7361 19015 7395
rect 19625 7361 19659 7395
rect 21097 7361 21131 7395
rect 21189 7361 21223 7395
rect 21282 7361 21316 7395
rect 21465 7361 21499 7395
rect 21557 7361 21591 7395
rect 21654 7361 21688 7395
rect 27077 7361 27111 7395
rect 28273 7361 28307 7395
rect 29745 7361 29779 7395
rect 31861 7361 31895 7395
rect 31953 7361 31987 7395
rect 32505 7361 32539 7395
rect 33333 7361 33367 7395
rect 34069 7361 34103 7395
rect 34529 7361 34563 7395
rect 37105 7361 37139 7395
rect 37473 7361 37507 7395
rect 40601 7361 40635 7395
rect 41429 7361 41463 7395
rect 15117 7293 15151 7327
rect 16589 7293 16623 7327
rect 17417 7293 17451 7327
rect 18245 7293 18279 7327
rect 19809 7293 19843 7327
rect 20453 7293 20487 7327
rect 22017 7293 22051 7327
rect 22753 7293 22787 7327
rect 23673 7293 23707 7327
rect 23765 7293 23799 7327
rect 24133 7293 24167 7327
rect 24961 7293 24995 7327
rect 25053 7293 25087 7327
rect 28917 7293 28951 7327
rect 30021 7293 30055 7327
rect 31769 7293 31803 7327
rect 32064 7293 32098 7327
rect 32413 7293 32447 7327
rect 32781 7293 32815 7327
rect 32873 7293 32907 7327
rect 34345 7293 34379 7327
rect 34805 7293 34839 7327
rect 36461 7293 36495 7327
rect 36553 7293 36587 7327
rect 38025 7293 38059 7327
rect 38761 7293 38795 7327
rect 39773 7293 39807 7327
rect 40049 7293 40083 7327
rect 14473 7225 14507 7259
rect 16773 7225 16807 7259
rect 18889 7225 18923 7259
rect 27169 7225 27203 7259
rect 28825 7225 28859 7259
rect 35817 7225 35851 7259
rect 39129 7225 39163 7259
rect 12541 7157 12575 7191
rect 14565 7157 14599 7191
rect 15945 7157 15979 7191
rect 16037 7157 16071 7191
rect 18061 7157 18095 7191
rect 21833 7157 21867 7191
rect 22569 7157 22603 7191
rect 23489 7157 23523 7191
rect 24317 7157 24351 7191
rect 27721 7157 27755 7191
rect 34253 7157 34287 7191
rect 35449 7157 35483 7191
rect 38209 7157 38243 7191
rect 40785 7157 40819 7191
rect 20440 6953 20474 6987
rect 22477 6953 22511 6987
rect 24133 6953 24167 6987
rect 25881 6953 25915 6987
rect 31033 6953 31067 6987
rect 32505 6953 32539 6987
rect 34713 6953 34747 6987
rect 35909 6953 35943 6987
rect 22661 6885 22695 6919
rect 35449 6885 35483 6919
rect 12541 6817 12575 6851
rect 13277 6817 13311 6851
rect 15577 6817 15611 6851
rect 17785 6817 17819 6851
rect 22845 6817 22879 6851
rect 23397 6817 23431 6851
rect 23489 6817 23523 6851
rect 24869 6817 24903 6851
rect 26709 6817 26743 6851
rect 28733 6817 28767 6851
rect 29561 6817 29595 6851
rect 30205 6817 30239 6851
rect 30573 6817 30607 6851
rect 30665 6817 30699 6851
rect 30849 6817 30883 6851
rect 33333 6817 33367 6851
rect 33977 6817 34011 6851
rect 36461 6817 36495 6851
rect 37381 6817 37415 6851
rect 39405 6817 39439 6851
rect 40049 6817 40083 6851
rect 40785 6817 40819 6851
rect 42809 6817 42843 6851
rect 10609 6749 10643 6783
rect 11161 6749 11195 6783
rect 11805 6749 11839 6783
rect 12449 6749 12483 6783
rect 13093 6749 13127 6783
rect 14841 6749 14875 6783
rect 15669 6749 15703 6783
rect 16497 6749 16531 6783
rect 17049 6749 17083 6783
rect 17969 6749 18003 6783
rect 18705 6749 18739 6783
rect 19257 6749 19291 6783
rect 19901 6749 19935 6783
rect 20177 6749 20211 6783
rect 22201 6749 22235 6783
rect 24225 6749 24259 6783
rect 25329 6749 25363 6783
rect 25513 6749 25547 6783
rect 25697 6749 25731 6783
rect 26065 6749 26099 6783
rect 30757 6749 30791 6783
rect 31125 6749 31159 6783
rect 31769 6749 31803 6783
rect 31861 6749 31895 6783
rect 33149 6749 33183 6783
rect 34069 6749 34103 6783
rect 34805 6749 34839 6783
rect 34897 6749 34931 6783
rect 35173 6749 35207 6783
rect 35265 6727 35299 6761
rect 35817 6749 35851 6783
rect 36645 6749 36679 6783
rect 42165 6749 42199 6783
rect 11253 6681 11287 6715
rect 13921 6681 13955 6715
rect 16313 6681 16347 6715
rect 22293 6681 22327 6715
rect 25605 6681 25639 6715
rect 26617 6681 26651 6715
rect 26985 6681 27019 6715
rect 32597 6681 32631 6715
rect 35081 6681 35115 6715
rect 37289 6681 37323 6715
rect 37657 6681 37691 6715
rect 40233 6681 40267 6715
rect 40417 6681 40451 6715
rect 12265 6613 12299 6647
rect 14289 6613 14323 6647
rect 15117 6613 15151 6647
rect 17141 6613 17175 6647
rect 18521 6613 18555 6647
rect 19349 6613 19383 6647
rect 22503 6613 22537 6647
rect 28917 6613 28951 6647
rect 29653 6613 29687 6647
rect 35725 6613 35759 6647
rect 39497 6613 39531 6647
rect 40601 6613 40635 6647
rect 41429 6613 41463 6647
rect 41521 6613 41555 6647
rect 42257 6613 42291 6647
rect 13737 6409 13771 6443
rect 15945 6409 15979 6443
rect 16681 6409 16715 6443
rect 18429 6409 18463 6443
rect 21741 6409 21775 6443
rect 23765 6409 23799 6443
rect 25145 6409 25179 6443
rect 26893 6409 26927 6443
rect 27261 6409 27295 6443
rect 27353 6409 27387 6443
rect 28825 6409 28859 6443
rect 30297 6409 30331 6443
rect 36553 6409 36587 6443
rect 16773 6341 16807 6375
rect 18337 6341 18371 6375
rect 22201 6341 22235 6375
rect 22417 6341 22451 6375
rect 31861 6341 31895 6375
rect 32689 6341 32723 6375
rect 33333 6341 33367 6375
rect 35081 6341 35115 6375
rect 37381 6341 37415 6375
rect 42809 6341 42843 6375
rect 9689 6273 9723 6307
rect 10793 6273 10827 6307
rect 12173 6273 12207 6307
rect 12725 6273 12759 6307
rect 13921 6273 13955 6307
rect 14565 6273 14599 6307
rect 16129 6273 16163 6307
rect 17785 6273 17819 6307
rect 19901 6273 19935 6307
rect 20729 6273 20763 6307
rect 22753 6273 22787 6307
rect 25237 6273 25271 6307
rect 26525 6273 26559 6307
rect 28273 6273 28307 6307
rect 29745 6273 29779 6307
rect 30481 6273 30515 6307
rect 31769 6273 31803 6307
rect 32597 6273 32631 6307
rect 33057 6273 33091 6307
rect 35909 6273 35943 6307
rect 36093 6273 36127 6307
rect 36185 6273 36219 6307
rect 36277 6273 36311 6307
rect 37933 6273 37967 6307
rect 38209 6273 38243 6307
rect 41797 6273 41831 6307
rect 42717 6273 42751 6307
rect 42993 6273 43027 6307
rect 10333 6205 10367 6239
rect 11345 6205 11379 6239
rect 13185 6205 13219 6239
rect 15393 6205 15427 6239
rect 17325 6205 17359 6239
rect 18981 6205 19015 6239
rect 19165 6205 19199 6239
rect 19809 6205 19843 6239
rect 21833 6205 21867 6239
rect 22017 6205 22051 6239
rect 23121 6205 23155 6239
rect 24409 6205 24443 6239
rect 24501 6205 24535 6239
rect 25789 6205 25823 6239
rect 27537 6205 27571 6239
rect 29469 6205 29503 6239
rect 31125 6205 31159 6239
rect 32413 6205 32447 6239
rect 35725 6205 35759 6239
rect 37289 6205 37323 6239
rect 38485 6205 38519 6239
rect 40233 6205 40267 6239
rect 40601 6205 40635 6239
rect 41245 6205 41279 6239
rect 41981 6205 42015 6239
rect 20545 6137 20579 6171
rect 22937 6137 22971 6171
rect 28917 6137 28951 6171
rect 9505 6069 9539 6103
rect 9781 6069 9815 6103
rect 11621 6069 11655 6103
rect 12725 6069 12759 6103
rect 14473 6069 14507 6103
rect 15209 6069 15243 6103
rect 21281 6069 21315 6103
rect 21373 6069 21407 6103
rect 22385 6069 22419 6103
rect 22569 6069 22603 6103
rect 23673 6069 23707 6103
rect 25973 6069 26007 6103
rect 31033 6069 31067 6103
rect 35173 6069 35207 6103
rect 36645 6069 36679 6103
rect 41153 6069 41187 6103
rect 42625 6069 42659 6103
rect 43177 6069 43211 6103
rect 10149 5865 10183 5899
rect 11161 5865 11195 5899
rect 14105 5865 14139 5899
rect 14841 5865 14875 5899
rect 18521 5865 18555 5899
rect 19257 5865 19291 5899
rect 20545 5865 20579 5899
rect 20729 5865 20763 5899
rect 25145 5865 25179 5899
rect 34713 5865 34747 5899
rect 36829 5865 36863 5899
rect 41521 5865 41555 5899
rect 23673 5797 23707 5831
rect 24409 5797 24443 5831
rect 28181 5797 28215 5831
rect 32137 5797 32171 5831
rect 38853 5797 38887 5831
rect 42993 5797 43027 5831
rect 12817 5729 12851 5763
rect 16313 5729 16347 5763
rect 17049 5729 17083 5763
rect 19349 5729 19383 5763
rect 21649 5729 21683 5763
rect 22385 5729 22419 5763
rect 22937 5729 22971 5763
rect 23121 5729 23155 5763
rect 30297 5729 30331 5763
rect 31033 5729 31067 5763
rect 34069 5729 34103 5763
rect 39129 5729 39163 5763
rect 41337 5729 41371 5763
rect 43545 5729 43579 5763
rect 9597 5661 9631 5695
rect 9965 5661 9999 5695
rect 10517 5661 10551 5695
rect 11437 5661 11471 5695
rect 11529 5661 11563 5695
rect 11897 5661 11931 5695
rect 12541 5661 12575 5695
rect 13553 5661 13587 5695
rect 14197 5661 14231 5695
rect 15853 5661 15887 5695
rect 17141 5661 17175 5695
rect 17877 5661 17911 5695
rect 18613 5661 18647 5695
rect 20177 5661 20211 5695
rect 20913 5661 20947 5695
rect 23857 5661 23891 5695
rect 24501 5661 24535 5695
rect 25513 5661 25547 5695
rect 26157 5661 26191 5695
rect 29561 5661 29595 5695
rect 31493 5661 31527 5695
rect 31585 5661 31619 5695
rect 31861 5661 31895 5695
rect 31953 5661 31987 5695
rect 34161 5661 34195 5695
rect 34529 5661 34563 5695
rect 35449 5661 35483 5695
rect 35817 5661 35851 5695
rect 36001 5661 36035 5695
rect 36093 5661 36127 5695
rect 36185 5661 36219 5695
rect 36921 5661 36955 5695
rect 38945 5661 38979 5695
rect 39681 5661 39715 5695
rect 40325 5661 40359 5695
rect 42073 5661 42107 5695
rect 42901 5661 42935 5695
rect 43729 5661 43763 5695
rect 44741 5661 44775 5695
rect 46581 5661 46615 5695
rect 11805 5593 11839 5627
rect 13369 5593 13403 5627
rect 15301 5593 15335 5627
rect 26893 5593 26927 5627
rect 30849 5593 30883 5627
rect 31769 5593 31803 5627
rect 32321 5593 32355 5627
rect 34345 5593 34379 5627
rect 34437 5593 34471 5627
rect 45293 5593 45327 5627
rect 9045 5525 9079 5559
rect 11989 5525 12023 5559
rect 16037 5525 16071 5559
rect 16405 5525 16439 5559
rect 17785 5525 17819 5559
rect 19993 5525 20027 5559
rect 20545 5525 20579 5559
rect 21465 5525 21499 5559
rect 22201 5525 22235 5559
rect 26065 5525 26099 5559
rect 26801 5525 26835 5559
rect 28917 5525 28951 5559
rect 29653 5525 29687 5559
rect 30481 5525 30515 5559
rect 30941 5525 30975 5559
rect 34805 5525 34839 5559
rect 35633 5525 35667 5559
rect 38209 5525 38243 5559
rect 39773 5525 39807 5559
rect 40785 5525 40819 5559
rect 42257 5525 42291 5559
rect 44281 5525 44315 5559
rect 45937 5525 45971 5559
rect 8953 5321 8987 5355
rect 10793 5321 10827 5355
rect 11529 5321 11563 5355
rect 14473 5321 14507 5355
rect 15209 5321 15243 5355
rect 15945 5321 15979 5355
rect 18153 5321 18187 5355
rect 18889 5321 18923 5355
rect 20821 5321 20855 5355
rect 21741 5321 21775 5355
rect 24041 5321 24075 5355
rect 25053 5321 25087 5355
rect 26249 5321 26283 5355
rect 32781 5321 32815 5355
rect 37473 5321 37507 5355
rect 41797 5321 41831 5355
rect 42717 5321 42751 5355
rect 8585 5253 8619 5287
rect 13001 5253 13035 5287
rect 13737 5253 13771 5287
rect 19257 5253 19291 5287
rect 22569 5253 22603 5287
rect 22753 5253 22787 5287
rect 27905 5253 27939 5287
rect 28181 5253 28215 5287
rect 30849 5253 30883 5287
rect 44097 5253 44131 5287
rect 8033 5185 8067 5219
rect 9965 5185 9999 5219
rect 10241 5185 10275 5219
rect 10885 5185 10919 5219
rect 11621 5185 11655 5219
rect 12265 5185 12299 5219
rect 12633 5185 12667 5219
rect 16681 5185 16715 5219
rect 17601 5185 17635 5219
rect 17877 5185 17911 5219
rect 18981 5185 19015 5219
rect 21189 5185 21223 5219
rect 21649 5185 21683 5219
rect 21833 5185 21867 5219
rect 24961 5185 24995 5219
rect 25697 5185 25731 5219
rect 26433 5185 26467 5219
rect 28917 5185 28951 5219
rect 29653 5185 29687 5219
rect 30573 5185 30607 5219
rect 32873 5185 32907 5219
rect 34069 5185 34103 5219
rect 34253 5185 34287 5219
rect 34345 5185 34379 5219
rect 34437 5185 34471 5219
rect 34897 5185 34931 5219
rect 36185 5185 36219 5219
rect 37381 5185 37415 5219
rect 38853 5185 38887 5219
rect 39681 5185 39715 5219
rect 40509 5185 40543 5219
rect 41061 5185 41095 5219
rect 42625 5185 42659 5219
rect 42901 5185 42935 5219
rect 44833 5185 44867 5219
rect 46949 5185 46983 5219
rect 9505 5117 9539 5151
rect 13185 5117 13219 5151
rect 13829 5117 13863 5151
rect 14565 5117 14599 5151
rect 15301 5117 15335 5151
rect 16773 5117 16807 5151
rect 18245 5117 18279 5151
rect 20729 5117 20763 5151
rect 21281 5117 21315 5151
rect 21373 5117 21407 5151
rect 21925 5117 21959 5151
rect 25237 5117 25271 5151
rect 27077 5117 27111 5151
rect 27629 5117 27663 5151
rect 28825 5117 28859 5151
rect 29561 5117 29595 5151
rect 30297 5117 30331 5151
rect 32597 5117 32631 5151
rect 33885 5117 33919 5151
rect 35633 5117 35667 5151
rect 36921 5117 36955 5151
rect 37657 5117 37691 5151
rect 38301 5117 38335 5151
rect 39037 5117 39071 5151
rect 40325 5117 40359 5151
rect 41153 5117 41187 5151
rect 42441 5117 42475 5151
rect 44005 5117 44039 5151
rect 44741 5117 44775 5151
rect 45477 5117 45511 5151
rect 45569 5117 45603 5151
rect 77493 5117 77527 5151
rect 16037 5049 16071 5083
rect 17417 5049 17451 5083
rect 36277 5049 36311 5083
rect 37013 5049 37047 5083
rect 41889 5049 41923 5083
rect 43361 5049 43395 5083
rect 9873 4981 9907 5015
rect 17969 4981 18003 5015
rect 24593 4981 24627 5015
rect 25421 4981 25455 5015
rect 26985 4981 27019 5015
rect 33333 4981 33367 5015
rect 34713 4981 34747 5015
rect 35449 4981 35483 5015
rect 39589 4981 39623 5015
rect 43085 4981 43119 5015
rect 46213 4981 46247 5015
rect 46305 4981 46339 5015
rect 76941 4981 76975 5015
rect 8953 4777 8987 4811
rect 9689 4777 9723 4811
rect 11897 4777 11931 4811
rect 12633 4777 12667 4811
rect 13369 4777 13403 4811
rect 14841 4777 14875 4811
rect 17049 4777 17083 4811
rect 22937 4777 22971 4811
rect 27813 4777 27847 4811
rect 31401 4777 31435 4811
rect 36185 4777 36219 4811
rect 38098 4777 38132 4811
rect 44741 4777 44775 4811
rect 76941 4777 76975 4811
rect 17785 4709 17819 4743
rect 18521 4709 18555 4743
rect 19257 4709 19291 4743
rect 27077 4709 27111 4743
rect 29561 4709 29595 4743
rect 33333 4709 33367 4743
rect 40601 4709 40635 4743
rect 8401 4641 8435 4675
rect 9137 4641 9171 4675
rect 11345 4641 11379 4675
rect 12081 4641 12115 4675
rect 12817 4641 12851 4675
rect 15209 4641 15243 4675
rect 15393 4641 15427 4675
rect 16405 4641 16439 4675
rect 17233 4641 17267 4675
rect 17877 4641 17911 4675
rect 20729 4641 20763 4675
rect 21373 4641 21407 4675
rect 23581 4641 23615 4675
rect 24685 4641 24719 4675
rect 25513 4641 25547 4675
rect 28365 4641 28399 4675
rect 28457 4641 28491 4675
rect 28917 4641 28951 4675
rect 29745 4641 29779 4675
rect 30757 4641 30791 4675
rect 31861 4641 31895 4675
rect 32045 4641 32079 4675
rect 32965 4641 32999 4675
rect 33977 4641 34011 4675
rect 34897 4641 34931 4675
rect 36829 4641 36863 4675
rect 37473 4641 37507 4675
rect 39865 4641 39899 4675
rect 39957 4641 39991 4675
rect 41521 4641 41555 4675
rect 43453 4641 43487 4675
rect 45109 4641 45143 4675
rect 45661 4641 45695 4675
rect 46581 4641 46615 4675
rect 47317 4641 47351 4675
rect 48145 4641 48179 4675
rect 7389 4573 7423 4607
rect 7665 4573 7699 4607
rect 10609 4573 10643 4607
rect 13461 4573 13495 4607
rect 14197 4573 14231 4607
rect 15117 4573 15151 4607
rect 15301 4573 15335 4607
rect 15761 4573 15795 4607
rect 18705 4573 18739 4607
rect 19441 4573 19475 4607
rect 20361 4573 20395 4607
rect 20637 4573 20671 4607
rect 21465 4573 21499 4607
rect 22293 4573 22327 4607
rect 25145 4573 25179 4607
rect 25973 4573 26007 4607
rect 26525 4573 26559 4607
rect 27261 4573 27295 4607
rect 31309 4573 31343 4607
rect 34161 4573 34195 4607
rect 34713 4573 34747 4607
rect 37749 4573 37783 4607
rect 37841 4573 37875 4607
rect 41797 4573 41831 4607
rect 42073 4573 42107 4607
rect 42809 4573 42843 4607
rect 44005 4573 44039 4607
rect 44189 4573 44223 4607
rect 46765 4573 46799 4607
rect 48053 4573 48087 4607
rect 48881 4573 48915 4607
rect 77585 4573 77619 4607
rect 10057 4505 10091 4539
rect 10425 4505 10459 4539
rect 22845 4505 22879 4539
rect 23305 4505 23339 4539
rect 31769 4505 31803 4539
rect 32413 4505 32447 4539
rect 40877 4505 40911 4539
rect 47409 4505 47443 4539
rect 6837 4437 6871 4471
rect 8217 4437 8251 4471
rect 11161 4437 11195 4471
rect 14105 4437 14139 4471
rect 15577 4437 15611 4471
rect 16313 4437 16347 4471
rect 19993 4437 20027 4471
rect 22109 4437 22143 4471
rect 23397 4437 23431 4471
rect 27905 4437 27939 4471
rect 28273 4437 28307 4471
rect 30297 4437 30331 4471
rect 33241 4437 33275 4471
rect 35449 4437 35483 4471
rect 41613 4437 41647 4471
rect 42625 4437 42659 4471
rect 43361 4437 43395 4471
rect 45937 4437 45971 4471
rect 48789 4437 48823 4471
rect 49525 4437 49559 4471
rect 19901 4233 19935 4267
rect 26525 4233 26559 4267
rect 38209 4233 38243 4267
rect 40233 4233 40267 4267
rect 7481 4165 7515 4199
rect 19441 4165 19475 4199
rect 20453 4165 20487 4199
rect 20653 4165 20687 4199
rect 21281 4165 21315 4199
rect 27721 4165 27755 4199
rect 30297 4165 30331 4199
rect 52653 4165 52687 4199
rect 6745 4097 6779 4131
rect 7849 4097 7883 4131
rect 9321 4097 9355 4131
rect 10793 4097 10827 4131
rect 12449 4097 12483 4131
rect 12541 4097 12575 4131
rect 13369 4097 13403 4131
rect 14841 4097 14875 4131
rect 15025 4097 15059 4131
rect 17233 4097 17267 4131
rect 21373 4097 21407 4131
rect 22845 4097 22879 4131
rect 24317 4097 24351 4131
rect 26433 4097 26467 4131
rect 26709 4097 26743 4131
rect 28457 4097 28491 4131
rect 32689 4097 32723 4131
rect 33057 4097 33091 4131
rect 33241 4097 33275 4131
rect 33425 4097 33459 4131
rect 34069 4097 34103 4131
rect 36093 4097 36127 4131
rect 36185 4097 36219 4131
rect 36829 4097 36863 4131
rect 38209 4097 38243 4131
rect 38393 4097 38427 4131
rect 38669 4097 38703 4131
rect 42717 4097 42751 4131
rect 45661 4097 45695 4131
rect 47869 4097 47903 4131
rect 50537 4097 50571 4131
rect 74733 4097 74767 4131
rect 76205 4097 76239 4131
rect 8033 4029 8067 4063
rect 8769 4029 8803 4063
rect 9505 4029 9539 4063
rect 10241 4029 10275 4063
rect 10885 4029 10919 4063
rect 11529 4029 11563 4063
rect 11713 4029 11747 4063
rect 12725 4029 12759 4063
rect 14381 4029 14415 4063
rect 15209 4029 15243 4063
rect 15393 4029 15427 4063
rect 16957 4029 16991 4063
rect 19993 4029 20027 4063
rect 20177 4029 20211 4063
rect 21557 4029 21591 4063
rect 21741 4029 21775 4063
rect 22385 4029 22419 4063
rect 23673 4029 23707 4063
rect 24593 4029 24627 4063
rect 26341 4029 26375 4063
rect 27353 4029 27387 4063
rect 27574 4029 27608 4063
rect 29101 4029 29135 4063
rect 30389 4029 30423 4063
rect 30573 4029 30607 4063
rect 30849 4029 30883 4063
rect 32413 4029 32447 4063
rect 33977 4029 34011 4063
rect 35081 4029 35115 4063
rect 35909 4029 35943 4063
rect 37289 4029 37323 4063
rect 39037 4029 39071 4063
rect 41705 4029 41739 4063
rect 41981 4029 42015 4063
rect 42165 4029 42199 4063
rect 43453 4029 43487 4063
rect 44189 4029 44223 4063
rect 44833 4029 44867 4063
rect 44925 4029 44959 4063
rect 45569 4029 45603 4063
rect 46949 4029 46983 4063
rect 47133 4029 47167 4063
rect 48513 4029 48547 4063
rect 49065 4029 49099 4063
rect 49893 4029 49927 4063
rect 65533 4029 65567 4063
rect 67649 4029 67683 4063
rect 71513 4029 71547 4063
rect 75929 4029 75963 4063
rect 77033 4029 77067 4063
rect 10057 3961 10091 3995
rect 15945 3961 15979 3995
rect 18153 3961 18187 3995
rect 26709 3961 26743 3995
rect 27261 3961 27295 3995
rect 29929 3961 29963 3995
rect 48053 3961 48087 3995
rect 6561 3893 6595 3927
rect 8585 3893 8619 3927
rect 12265 3893 12299 3927
rect 19533 3893 19567 3927
rect 20637 3893 20671 3927
rect 20821 3893 20855 3927
rect 20913 3893 20947 3927
rect 27445 3893 27479 3927
rect 31401 3893 31435 3927
rect 33057 3893 33091 3927
rect 36553 3893 36587 3927
rect 44097 3893 44131 3927
rect 46305 3893 46339 3927
rect 46397 3893 46431 3927
rect 47777 3893 47811 3927
rect 49249 3893 49283 3927
rect 49985 3893 50019 3927
rect 52745 3893 52779 3927
rect 66177 3893 66211 3927
rect 68201 3893 68235 3927
rect 72065 3893 72099 3927
rect 4905 3689 4939 3723
rect 6009 3689 6043 3723
rect 10885 3689 10919 3723
rect 11897 3689 11931 3723
rect 14841 3689 14875 3723
rect 28457 3689 28491 3723
rect 28733 3689 28767 3723
rect 32137 3689 32171 3723
rect 34161 3689 34195 3723
rect 34253 3689 34287 3723
rect 34713 3689 34747 3723
rect 35817 3689 35851 3723
rect 44833 3689 44867 3723
rect 48881 3689 48915 3723
rect 67925 3689 67959 3723
rect 71697 3689 71731 3723
rect 77585 3689 77619 3723
rect 7481 3621 7515 3655
rect 10793 3621 10827 3655
rect 14105 3621 14139 3655
rect 19809 3621 19843 3655
rect 25605 3621 25639 3655
rect 31953 3621 31987 3655
rect 41613 3621 41647 3655
rect 5457 3553 5491 3587
rect 6837 3553 6871 3587
rect 9045 3553 9079 3587
rect 12265 3553 12299 3587
rect 13737 3553 13771 3587
rect 14289 3553 14323 3587
rect 15485 3553 15519 3587
rect 15669 3553 15703 3587
rect 17877 3553 17911 3587
rect 18705 3553 18739 3587
rect 20821 3553 20855 3587
rect 22845 3553 22879 3587
rect 26157 3553 26191 3587
rect 26341 3553 26375 3587
rect 29377 3553 29411 3587
rect 32413 3553 32447 3587
rect 34621 3553 34655 3587
rect 35265 3553 35299 3587
rect 36829 3553 36863 3587
rect 38669 3553 38703 3587
rect 39681 3553 39715 3587
rect 41337 3553 41371 3587
rect 41889 3553 41923 3587
rect 42257 3553 42291 3587
rect 42533 3553 42567 3587
rect 44005 3553 44039 3587
rect 44281 3553 44315 3587
rect 44373 3553 44407 3587
rect 46765 3553 46799 3587
rect 49985 3553 50019 3587
rect 72433 3553 72467 3587
rect 77033 3553 77067 3587
rect 4721 3485 4755 3519
rect 5089 3485 5123 3519
rect 6101 3485 6135 3519
rect 7665 3485 7699 3519
rect 8217 3485 8251 3519
rect 8401 3485 8435 3519
rect 9689 3485 9723 3519
rect 10241 3485 10275 3519
rect 11437 3485 11471 3519
rect 11713 3485 11747 3519
rect 11989 3485 12023 3519
rect 13921 3485 13955 3519
rect 15393 3485 15427 3519
rect 18153 3485 18187 3519
rect 18245 3485 18279 3519
rect 19993 3485 20027 3519
rect 20361 3485 20395 3519
rect 21925 3485 21959 3519
rect 25145 3485 25179 3519
rect 25329 3485 25363 3519
rect 26709 3485 26743 3519
rect 28641 3485 28675 3519
rect 29101 3485 29135 3519
rect 30481 3485 30515 3519
rect 34437 3485 34471 3519
rect 36369 3485 36403 3519
rect 37749 3485 37783 3519
rect 39221 3485 39255 3519
rect 41981 3485 42015 3519
rect 44465 3485 44499 3519
rect 45477 3485 45511 3519
rect 45937 3485 45971 3519
rect 46489 3485 46523 3519
rect 48329 3485 48363 3519
rect 49801 3485 49835 3519
rect 52285 3485 52319 3519
rect 52469 3485 52503 3519
rect 53665 3485 53699 3519
rect 54309 3485 54343 3519
rect 54401 3485 54435 3519
rect 57989 3485 58023 3519
rect 58173 3485 58207 3519
rect 61945 3485 61979 3519
rect 62129 3485 62163 3519
rect 65717 3485 65751 3519
rect 67189 3485 67223 3519
rect 67833 3485 67867 3519
rect 68477 3485 68511 3519
rect 69121 3485 69155 3519
rect 69765 3485 69799 3519
rect 69857 3485 69891 3519
rect 72249 3485 72283 3519
rect 75101 3485 75135 3519
rect 76665 3485 76699 3519
rect 8953 3417 8987 3451
rect 15945 3417 15979 3451
rect 25605 3417 25639 3451
rect 26065 3417 26099 3451
rect 26985 3417 27019 3451
rect 31401 3417 31435 3451
rect 32321 3417 32355 3451
rect 32689 3417 32723 3451
rect 35081 3417 35115 3451
rect 35725 3417 35759 3451
rect 49249 3417 49283 3451
rect 75469 3417 75503 3451
rect 5273 3349 5307 3383
rect 6745 3349 6779 3383
rect 10057 3349 10091 3383
rect 15025 3349 15059 3383
rect 16221 3349 16255 3383
rect 16405 3349 16439 3383
rect 20269 3349 20303 3383
rect 23857 3349 23891 3383
rect 25421 3349 25455 3383
rect 25697 3349 25731 3383
rect 26617 3349 26651 3383
rect 32121 3349 32155 3383
rect 35173 3349 35207 3383
rect 40785 3349 40819 3383
rect 41153 3349 41187 3383
rect 41245 3349 41279 3383
rect 44925 3349 44959 3383
rect 46121 3349 46155 3383
rect 50629 3349 50663 3383
rect 51733 3349 51767 3383
rect 53113 3349 53147 3383
rect 55045 3349 55079 3383
rect 57437 3349 57471 3383
rect 58817 3349 58851 3383
rect 61393 3349 61427 3383
rect 62773 3349 62807 3383
rect 65165 3349 65199 3383
rect 70501 3349 70535 3383
rect 73077 3349 73111 3383
rect 74549 3349 74583 3383
rect 4905 3145 4939 3179
rect 6377 3145 6411 3179
rect 8217 3145 8251 3179
rect 12541 3145 12575 3179
rect 20085 3145 20119 3179
rect 22963 3145 22997 3179
rect 27077 3145 27111 3179
rect 28089 3145 28123 3179
rect 28549 3145 28583 3179
rect 30481 3145 30515 3179
rect 32689 3145 32723 3179
rect 33425 3145 33459 3179
rect 33517 3145 33551 3179
rect 34069 3145 34103 3179
rect 34161 3145 34195 3179
rect 38393 3145 38427 3179
rect 40417 3145 40451 3179
rect 41337 3145 41371 3179
rect 43177 3145 43211 3179
rect 45385 3145 45419 3179
rect 45661 3145 45695 3179
rect 48053 3145 48087 3179
rect 50077 3145 50111 3179
rect 51273 3145 51307 3179
rect 52009 3145 52043 3179
rect 53665 3145 53699 3179
rect 57345 3145 57379 3179
rect 58081 3145 58115 3179
rect 60933 3145 60967 3179
rect 61669 3145 61703 3179
rect 64705 3145 64739 3179
rect 65441 3145 65475 3179
rect 67189 3145 67223 3179
rect 69121 3145 69155 3179
rect 74457 3145 74491 3179
rect 10793 3077 10827 3111
rect 13369 3077 13403 3111
rect 17417 3077 17451 3111
rect 18613 3077 18647 3111
rect 22017 3077 22051 3111
rect 22201 3077 22235 3111
rect 22385 3077 22419 3111
rect 22753 3077 22787 3111
rect 30021 3077 30055 3111
rect 31217 3077 31251 3111
rect 35633 3077 35667 3111
rect 37657 3077 37691 3111
rect 43821 3077 43855 3111
rect 4353 3009 4387 3043
rect 5089 3009 5123 3043
rect 6561 3009 6595 3043
rect 7113 3009 7147 3043
rect 8401 3009 8435 3043
rect 9045 3009 9079 3043
rect 9781 3009 9815 3043
rect 10517 3009 10551 3043
rect 12725 3009 12759 3043
rect 12909 3009 12943 3043
rect 13001 3009 13035 3043
rect 13093 3009 13127 3043
rect 14933 3009 14967 3043
rect 18337 3009 18371 3043
rect 20177 3009 20211 3043
rect 22293 3009 22327 3043
rect 22569 3009 22603 3043
rect 23213 3009 23247 3043
rect 25053 3009 25087 3043
rect 25329 3009 25363 3043
rect 27261 3009 27295 3043
rect 27353 3009 27387 3043
rect 27537 3009 27571 3043
rect 28181 3009 28215 3043
rect 28273 3009 28307 3043
rect 30297 3009 30331 3043
rect 30389 3009 30423 3043
rect 30665 3009 30699 3043
rect 33885 3009 33919 3043
rect 34069 3009 34103 3043
rect 35909 3009 35943 3043
rect 36093 3009 36127 3043
rect 37933 3009 37967 3043
rect 38209 3009 38243 3043
rect 38669 3009 38703 3043
rect 40969 3009 41003 3043
rect 41418 3009 41452 3043
rect 43545 3009 43579 3043
rect 43913 3009 43947 3043
rect 45569 3009 45603 3043
rect 45845 3009 45879 3043
rect 46121 3009 46155 3043
rect 47501 3009 47535 3043
rect 48329 3009 48363 3043
rect 49801 3009 49835 3043
rect 50629 3009 50663 3043
rect 51089 3009 51123 3043
rect 51457 3009 51491 3043
rect 52101 3009 52135 3043
rect 53849 3009 53883 3043
rect 54033 3009 54067 3043
rect 56057 3009 56091 3043
rect 57161 3009 57195 3043
rect 57437 3009 57471 3043
rect 60749 3009 60783 3043
rect 61117 3009 61151 3043
rect 61761 3009 61795 3043
rect 64521 3009 64555 3043
rect 64889 3009 64923 3043
rect 65533 3009 65567 3043
rect 67005 3009 67039 3043
rect 67649 3009 67683 3043
rect 69305 3009 69339 3043
rect 69489 3009 69523 3043
rect 71513 3009 71547 3043
rect 72985 3009 73019 3043
rect 74273 3009 74307 3043
rect 74549 3009 74583 3043
rect 76665 3009 76699 3043
rect 5825 2941 5859 2975
rect 7665 2941 7699 2975
rect 8953 2941 8987 2975
rect 12265 2941 12299 2975
rect 15209 2941 15243 2975
rect 16681 2941 16715 2975
rect 16865 2941 16899 2975
rect 17601 2941 17635 2975
rect 20453 2941 20487 2975
rect 23489 2941 23523 2975
rect 25605 2941 25639 2975
rect 27445 2941 27479 2975
rect 27905 2941 27939 2975
rect 30941 2941 30975 2975
rect 33609 2941 33643 2975
rect 38945 2941 38979 2975
rect 40693 2941 40727 2975
rect 40877 2941 40911 2975
rect 41705 2941 41739 2975
rect 43729 2941 43763 2975
rect 45109 2941 45143 2975
rect 46489 2941 46523 2975
rect 48789 2941 48823 2975
rect 52561 2941 52595 2975
rect 54493 2941 54527 2975
rect 62221 2941 62255 2975
rect 65993 2941 66027 2975
rect 68017 2941 68051 2975
rect 69949 2941 69983 2975
rect 71973 2941 72007 2975
rect 75469 2941 75503 2975
rect 77309 2941 77343 2975
rect 5641 2873 5675 2907
rect 9689 2873 9723 2907
rect 27721 2873 27755 2907
rect 33057 2873 33091 2907
rect 48145 2873 48179 2907
rect 75193 2873 75227 2907
rect 7481 2805 7515 2839
rect 10425 2805 10459 2839
rect 14841 2805 14875 2839
rect 18245 2805 18279 2839
rect 21925 2805 21959 2839
rect 22937 2805 22971 2839
rect 23121 2805 23155 2839
rect 24961 2805 24995 2839
rect 25237 2805 25271 2839
rect 28457 2805 28491 2839
rect 30849 2805 30883 2839
rect 36185 2805 36219 2839
rect 43361 2805 43395 2839
rect 43545 2805 43579 2839
rect 55505 2805 55539 2839
rect 59369 2805 59403 2839
rect 70961 2805 70995 2839
rect 76757 2805 76791 2839
rect 3801 2601 3835 2635
rect 4537 2601 4571 2635
rect 4905 2601 4939 2635
rect 6377 2601 6411 2635
rect 8217 2601 8251 2635
rect 10057 2601 10091 2635
rect 12449 2601 12483 2635
rect 15117 2601 15151 2635
rect 17601 2601 17635 2635
rect 21373 2601 21407 2635
rect 33977 2601 34011 2635
rect 41705 2601 41739 2635
rect 44833 2601 44867 2635
rect 49985 2601 50019 2635
rect 70869 2601 70903 2635
rect 74089 2601 74123 2635
rect 76849 2601 76883 2635
rect 11253 2533 11287 2567
rect 18521 2533 18555 2567
rect 23673 2533 23707 2567
rect 25513 2533 25547 2567
rect 30665 2533 30699 2567
rect 35817 2533 35851 2567
rect 36553 2533 36587 2567
rect 40969 2533 41003 2567
rect 48145 2533 48179 2567
rect 50721 2533 50755 2567
rect 3985 2465 4019 2499
rect 5825 2465 5859 2499
rect 6561 2465 6595 2499
rect 9689 2465 9723 2499
rect 11805 2465 11839 2499
rect 12909 2465 12943 2499
rect 13093 2465 13127 2499
rect 15669 2465 15703 2499
rect 15853 2465 15887 2499
rect 18153 2465 18187 2499
rect 19349 2465 19383 2499
rect 20729 2465 20763 2499
rect 22753 2465 22787 2499
rect 24409 2465 24443 2499
rect 25605 2465 25639 2499
rect 26249 2465 26283 2499
rect 26801 2465 26835 2499
rect 28273 2465 28307 2499
rect 29837 2465 29871 2499
rect 32229 2465 32263 2499
rect 33425 2465 33459 2499
rect 37565 2465 37599 2499
rect 39957 2465 39991 2499
rect 40601 2465 40635 2499
rect 41153 2465 41187 2499
rect 43821 2465 43855 2499
rect 45385 2465 45419 2499
rect 46397 2465 46431 2499
rect 47961 2465 47995 2499
rect 49433 2465 49467 2499
rect 52101 2465 52135 2499
rect 54033 2465 54067 2499
rect 58173 2465 58207 2499
rect 59277 2465 59311 2499
rect 61761 2465 61795 2499
rect 65533 2465 65567 2499
rect 67649 2465 67683 2499
rect 69489 2465 69523 2499
rect 72617 2465 72651 2499
rect 73169 2465 73203 2499
rect 73537 2465 73571 2499
rect 75745 2465 75779 2499
rect 77401 2465 77435 2499
rect 3617 2397 3651 2431
rect 4721 2397 4755 2431
rect 5089 2397 5123 2431
rect 7665 2397 7699 2431
rect 8401 2397 8435 2431
rect 9137 2397 9171 2431
rect 10333 2397 10367 2431
rect 10609 2397 10643 2431
rect 11621 2397 11655 2431
rect 12265 2397 12299 2431
rect 12817 2397 12851 2431
rect 13369 2397 13403 2431
rect 14657 2397 14691 2431
rect 16037 2397 16071 2431
rect 18613 2397 18647 2431
rect 20177 2397 20211 2431
rect 20453 2397 20487 2431
rect 21557 2397 21591 2431
rect 22385 2397 22419 2431
rect 22569 2397 22603 2431
rect 23489 2397 23523 2431
rect 24593 2397 24627 2431
rect 25329 2397 25363 2431
rect 26341 2397 26375 2431
rect 27905 2397 27939 2431
rect 30205 2397 30239 2431
rect 30849 2397 30883 2431
rect 32873 2397 32907 2431
rect 35265 2397 35299 2431
rect 35633 2397 35667 2431
rect 36001 2397 36035 2431
rect 37933 2397 37967 2431
rect 38301 2397 38335 2431
rect 38853 2397 38887 2431
rect 38945 2397 38979 2431
rect 39681 2397 39715 2431
rect 40785 2397 40819 2431
rect 41797 2397 41831 2431
rect 42993 2397 43027 2431
rect 43361 2397 43395 2431
rect 45201 2397 45235 2431
rect 45293 2397 45327 2431
rect 45937 2397 45971 2431
rect 48329 2397 48363 2431
rect 49893 2397 49927 2431
rect 50537 2397 50571 2431
rect 53021 2397 53055 2431
rect 55045 2397 55079 2431
rect 55505 2397 55539 2431
rect 58633 2397 58667 2431
rect 58817 2397 58851 2431
rect 62773 2397 62807 2431
rect 63233 2397 63267 2431
rect 66269 2397 66303 2431
rect 68293 2397 68327 2431
rect 70501 2397 70535 2431
rect 70685 2397 70719 2431
rect 73077 2397 73111 2431
rect 76205 2397 76239 2431
rect 5641 2329 5675 2363
rect 7481 2329 7515 2363
rect 11161 2329 11195 2363
rect 13645 2329 13679 2363
rect 17233 2329 17267 2363
rect 23765 2329 23799 2363
rect 28825 2329 28859 2363
rect 34253 2329 34287 2363
rect 7113 2261 7147 2295
rect 8953 2261 8987 2295
rect 11713 2261 11747 2295
rect 15209 2261 15243 2295
rect 15577 2261 15611 2295
rect 17969 2261 18003 2295
rect 18061 2261 18095 2295
rect 20361 2261 20395 2295
rect 20637 2261 20671 2295
rect 22109 2261 22143 2295
rect 22201 2261 22235 2295
rect 23397 2261 23431 2295
rect 25145 2261 25179 2295
rect 28089 2261 28123 2295
rect 31401 2261 31435 2295
rect 38301 2261 38335 2295
rect 47409 2261 47443 2295
<< metal1 >>
rect 2024 37562 77924 37584
rect 2024 37510 5134 37562
rect 5186 37510 5198 37562
rect 5250 37510 5262 37562
rect 5314 37510 5326 37562
rect 5378 37510 5390 37562
rect 5442 37510 35854 37562
rect 35906 37510 35918 37562
rect 35970 37510 35982 37562
rect 36034 37510 36046 37562
rect 36098 37510 36110 37562
rect 36162 37510 66574 37562
rect 66626 37510 66638 37562
rect 66690 37510 66702 37562
rect 66754 37510 66766 37562
rect 66818 37510 66830 37562
rect 66882 37510 77924 37562
rect 2024 37488 77924 37510
rect 2222 37272 2228 37324
rect 2280 37312 2286 37324
rect 2501 37315 2559 37321
rect 2501 37312 2513 37315
rect 2280 37284 2513 37312
rect 2280 37272 2286 37284
rect 2501 37281 2513 37284
rect 2547 37281 2559 37315
rect 2501 37275 2559 37281
rect 13262 37272 13268 37324
rect 13320 37312 13326 37324
rect 13541 37315 13599 37321
rect 13541 37312 13553 37315
rect 13320 37284 13553 37312
rect 13320 37272 13326 37284
rect 13541 37281 13553 37284
rect 13587 37281 13599 37315
rect 13541 37275 13599 37281
rect 33502 37272 33508 37324
rect 33560 37312 33566 37324
rect 34057 37315 34115 37321
rect 34057 37312 34069 37315
rect 33560 37284 34069 37312
rect 33560 37272 33566 37284
rect 34057 37281 34069 37284
rect 34103 37281 34115 37315
rect 34057 37275 34115 37281
rect 39022 37272 39028 37324
rect 39080 37312 39086 37324
rect 39577 37315 39635 37321
rect 39577 37312 39589 37315
rect 39080 37284 39589 37312
rect 39080 37272 39086 37284
rect 39577 37281 39589 37284
rect 39623 37281 39635 37315
rect 39577 37275 39635 37281
rect 3510 37204 3516 37256
rect 3568 37204 3574 37256
rect 5902 37204 5908 37256
rect 5960 37204 5966 37256
rect 7006 37204 7012 37256
rect 7064 37204 7070 37256
rect 7742 37204 7748 37256
rect 7800 37244 7806 37256
rect 7837 37247 7895 37253
rect 7837 37244 7849 37247
rect 7800 37216 7849 37244
rect 7800 37204 7806 37216
rect 7837 37213 7849 37216
rect 7883 37213 7895 37247
rect 7837 37207 7895 37213
rect 7926 37204 7932 37256
rect 7984 37244 7990 37256
rect 8757 37247 8815 37253
rect 8757 37244 8769 37247
rect 7984 37216 8769 37244
rect 7984 37204 7990 37216
rect 8757 37213 8769 37216
rect 8803 37213 8815 37247
rect 8757 37207 8815 37213
rect 11333 37247 11391 37253
rect 11333 37213 11345 37247
rect 11379 37244 11391 37247
rect 11422 37244 11428 37256
rect 11379 37216 11428 37244
rect 11379 37213 11391 37216
rect 11333 37207 11391 37213
rect 11422 37204 11428 37216
rect 11480 37204 11486 37256
rect 11882 37204 11888 37256
rect 11940 37244 11946 37256
rect 12069 37247 12127 37253
rect 12069 37244 12081 37247
rect 11940 37216 12081 37244
rect 11940 37204 11946 37216
rect 12069 37213 12081 37216
rect 12115 37213 12127 37247
rect 12069 37207 12127 37213
rect 14550 37204 14556 37256
rect 14608 37204 14614 37256
rect 15102 37204 15108 37256
rect 15160 37244 15166 37256
rect 15197 37247 15255 37253
rect 15197 37244 15209 37247
rect 15160 37216 15209 37244
rect 15160 37204 15166 37216
rect 15197 37213 15209 37216
rect 15243 37213 15255 37247
rect 15197 37207 15255 37213
rect 18690 37204 18696 37256
rect 18748 37204 18754 37256
rect 18782 37204 18788 37256
rect 18840 37244 18846 37256
rect 19521 37247 19579 37253
rect 19521 37244 19533 37247
rect 18840 37216 19533 37244
rect 18840 37204 18846 37216
rect 19521 37213 19533 37216
rect 19567 37213 19579 37247
rect 19521 37207 19579 37213
rect 20622 37204 20628 37256
rect 20680 37244 20686 37256
rect 20901 37247 20959 37253
rect 20901 37244 20913 37247
rect 20680 37216 20913 37244
rect 20680 37204 20686 37216
rect 20901 37213 20913 37216
rect 20947 37213 20959 37247
rect 20901 37207 20959 37213
rect 21910 37204 21916 37256
rect 21968 37204 21974 37256
rect 22462 37204 22468 37256
rect 22520 37244 22526 37256
rect 22741 37247 22799 37253
rect 22741 37244 22753 37247
rect 22520 37216 22753 37244
rect 22520 37204 22526 37216
rect 22741 37213 22753 37216
rect 22787 37213 22799 37247
rect 22741 37207 22799 37213
rect 26050 37204 26056 37256
rect 26108 37244 26114 37256
rect 26237 37247 26295 37253
rect 26237 37244 26249 37247
rect 26108 37216 26249 37244
rect 26108 37204 26114 37216
rect 26237 37213 26249 37216
rect 26283 37213 26295 37247
rect 26237 37207 26295 37213
rect 27982 37204 27988 37256
rect 28040 37244 28046 37256
rect 28261 37247 28319 37253
rect 28261 37244 28273 37247
rect 28040 37216 28273 37244
rect 28040 37204 28046 37216
rect 28261 37213 28273 37216
rect 28307 37213 28319 37247
rect 28261 37207 28319 37213
rect 29270 37204 29276 37256
rect 29328 37204 29334 37256
rect 31662 37204 31668 37256
rect 31720 37244 31726 37256
rect 31757 37247 31815 37253
rect 31757 37244 31769 37247
rect 31720 37216 31769 37244
rect 31720 37204 31726 37216
rect 31757 37213 31769 37216
rect 31803 37213 31815 37247
rect 31757 37207 31815 37213
rect 32766 37204 32772 37256
rect 32824 37204 32830 37256
rect 33778 37204 33784 37256
rect 33836 37204 33842 37256
rect 36817 37247 36875 37253
rect 36817 37213 36829 37247
rect 36863 37244 36875 37247
rect 36998 37244 37004 37256
rect 36863 37216 37004 37244
rect 36863 37213 36875 37216
rect 36817 37207 36875 37213
rect 36998 37204 37004 37216
rect 37056 37204 37062 37256
rect 37182 37204 37188 37256
rect 37240 37244 37246 37256
rect 37553 37247 37611 37253
rect 37553 37244 37565 37247
rect 37240 37216 37565 37244
rect 37240 37204 37246 37216
rect 37553 37213 37565 37216
rect 37599 37213 37611 37247
rect 37553 37207 37611 37213
rect 39114 37204 39120 37256
rect 39172 37204 39178 37256
rect 40862 37204 40868 37256
rect 40920 37244 40926 37256
rect 40957 37247 41015 37253
rect 40957 37244 40969 37247
rect 40920 37216 40969 37244
rect 40920 37204 40926 37216
rect 40957 37213 40969 37216
rect 41003 37213 41015 37247
rect 40957 37207 41015 37213
rect 41046 37204 41052 37256
rect 41104 37244 41110 37256
rect 41877 37247 41935 37253
rect 41877 37244 41889 37247
rect 41104 37216 41889 37244
rect 41104 37204 41110 37216
rect 41877 37213 41889 37216
rect 41923 37213 41935 37247
rect 41877 37207 41935 37213
rect 43346 37204 43352 37256
rect 43404 37204 43410 37256
rect 46474 37204 46480 37256
rect 46532 37204 46538 37256
rect 48222 37204 48228 37256
rect 48280 37244 48286 37256
rect 48501 37247 48559 37253
rect 48501 37244 48513 37247
rect 48280 37216 48513 37244
rect 48280 37204 48286 37216
rect 48501 37213 48513 37216
rect 48547 37213 48559 37247
rect 48501 37207 48559 37213
rect 51902 37204 51908 37256
rect 51960 37244 51966 37256
rect 51997 37247 52055 37253
rect 51997 37244 52009 37247
rect 51960 37216 52009 37244
rect 51960 37204 51966 37216
rect 51997 37213 52009 37216
rect 52043 37213 52055 37247
rect 51997 37207 52055 37213
rect 52086 37204 52092 37256
rect 52144 37244 52150 37256
rect 52917 37247 52975 37253
rect 52917 37244 52929 37247
rect 52144 37216 52929 37244
rect 52144 37204 52150 37216
rect 52917 37213 52929 37216
rect 52963 37213 52975 37247
rect 52917 37207 52975 37213
rect 53834 37204 53840 37256
rect 53892 37204 53898 37256
rect 55582 37204 55588 37256
rect 55640 37244 55646 37256
rect 56229 37247 56287 37253
rect 56229 37244 56241 37247
rect 55640 37216 56241 37244
rect 55640 37204 55646 37216
rect 56229 37213 56241 37216
rect 56275 37213 56287 37247
rect 56229 37207 56287 37213
rect 58802 37204 58808 37256
rect 58860 37204 58866 37256
rect 15010 37136 15016 37188
rect 15068 37176 15074 37188
rect 16117 37179 16175 37185
rect 16117 37176 16129 37179
rect 15068 37148 16129 37176
rect 15068 37136 15074 37148
rect 16117 37145 16129 37148
rect 16163 37145 16175 37179
rect 16117 37139 16175 37145
rect 22554 37136 22560 37188
rect 22612 37176 22618 37188
rect 23661 37179 23719 37185
rect 23661 37176 23673 37179
rect 22612 37148 23673 37176
rect 22612 37136 22618 37148
rect 23661 37145 23673 37148
rect 23707 37145 23719 37179
rect 23661 37139 23719 37145
rect 26142 37136 26148 37188
rect 26200 37176 26206 37188
rect 27157 37179 27215 37185
rect 27157 37176 27169 37179
rect 26200 37148 27169 37176
rect 26200 37136 26206 37148
rect 27157 37145 27169 37148
rect 27203 37145 27215 37179
rect 27157 37139 27215 37145
rect 42702 37136 42708 37188
rect 42760 37176 42766 37188
rect 44269 37179 44327 37185
rect 44269 37176 44281 37179
rect 42760 37148 44281 37176
rect 42760 37136 42766 37148
rect 44269 37145 44281 37148
rect 44315 37145 44327 37179
rect 44269 37139 44327 37145
rect 46382 37136 46388 37188
rect 46440 37176 46446 37188
rect 47397 37179 47455 37185
rect 47397 37176 47409 37179
rect 46440 37148 47409 37176
rect 46440 37136 46446 37148
rect 47397 37145 47409 37148
rect 47443 37145 47455 37179
rect 47397 37139 47455 37145
rect 48130 37136 48136 37188
rect 48188 37176 48194 37188
rect 49421 37179 49479 37185
rect 49421 37176 49433 37179
rect 48188 37148 49433 37176
rect 48188 37136 48194 37148
rect 49421 37145 49433 37148
rect 49467 37145 49479 37179
rect 49421 37139 49479 37145
rect 53742 37136 53748 37188
rect 53800 37176 53806 37188
rect 54757 37179 54815 37185
rect 54757 37176 54769 37179
rect 53800 37148 54769 37176
rect 53800 37136 53806 37148
rect 54757 37145 54769 37148
rect 54803 37145 54815 37179
rect 54757 37139 54815 37145
rect 55674 37136 55680 37188
rect 55732 37176 55738 37188
rect 57149 37179 57207 37185
rect 57149 37176 57161 37179
rect 55732 37148 57161 37176
rect 55732 37136 55738 37148
rect 57149 37145 57161 37148
rect 57195 37145 57207 37179
rect 57149 37139 57207 37145
rect 57422 37136 57428 37188
rect 57480 37176 57486 37188
rect 59725 37179 59783 37185
rect 59725 37176 59737 37179
rect 57480 37148 59737 37176
rect 57480 37136 57486 37148
rect 59725 37145 59737 37148
rect 59771 37145 59783 37179
rect 59725 37139 59783 37145
rect 2024 37018 77924 37040
rect 2024 36966 5794 37018
rect 5846 36966 5858 37018
rect 5910 36966 5922 37018
rect 5974 36966 5986 37018
rect 6038 36966 6050 37018
rect 6102 36966 36514 37018
rect 36566 36966 36578 37018
rect 36630 36966 36642 37018
rect 36694 36966 36706 37018
rect 36758 36966 36770 37018
rect 36822 36966 67234 37018
rect 67286 36966 67298 37018
rect 67350 36966 67362 37018
rect 67414 36966 67426 37018
rect 67478 36966 67490 37018
rect 67542 36966 77924 37018
rect 2024 36944 77924 36966
rect 7742 36864 7748 36916
rect 7800 36864 7806 36916
rect 11882 36864 11888 36916
rect 11940 36864 11946 36916
rect 15102 36864 15108 36916
rect 15160 36864 15166 36916
rect 18690 36864 18696 36916
rect 18748 36904 18754 36916
rect 19061 36907 19119 36913
rect 19061 36904 19073 36907
rect 18748 36876 19073 36904
rect 18748 36864 18754 36876
rect 19061 36873 19073 36876
rect 19107 36873 19119 36907
rect 19061 36867 19119 36873
rect 22462 36864 22468 36916
rect 22520 36864 22526 36916
rect 26050 36864 26056 36916
rect 26108 36904 26114 36916
rect 26145 36907 26203 36913
rect 26145 36904 26157 36907
rect 26108 36876 26157 36904
rect 26108 36864 26114 36876
rect 26145 36873 26157 36876
rect 26191 36873 26203 36907
rect 26145 36867 26203 36873
rect 29656 36876 30604 36904
rect 4062 36796 4068 36848
rect 4120 36836 4126 36848
rect 4341 36839 4399 36845
rect 4341 36836 4353 36839
rect 4120 36808 4353 36836
rect 4120 36796 4126 36808
rect 4341 36805 4353 36808
rect 4387 36805 4399 36839
rect 4341 36799 4399 36805
rect 9582 36796 9588 36848
rect 9640 36836 9646 36848
rect 9861 36839 9919 36845
rect 9861 36836 9873 36839
rect 9640 36808 9873 36836
rect 9640 36796 9646 36808
rect 9861 36805 9873 36808
rect 9907 36805 9919 36839
rect 9861 36799 9919 36805
rect 16942 36796 16948 36848
rect 17000 36836 17006 36848
rect 17957 36839 18015 36845
rect 17957 36836 17969 36839
rect 17000 36808 17969 36836
rect 17000 36796 17006 36808
rect 17957 36805 17969 36808
rect 18003 36805 18015 36839
rect 17957 36799 18015 36805
rect 24302 36796 24308 36848
rect 24360 36836 24366 36848
rect 24581 36839 24639 36845
rect 24581 36836 24593 36839
rect 24360 36808 24593 36836
rect 24360 36796 24366 36808
rect 24581 36805 24593 36808
rect 24627 36805 24639 36839
rect 24581 36799 24639 36805
rect 5445 36771 5503 36777
rect 5445 36737 5457 36771
rect 5491 36768 5503 36771
rect 7561 36771 7619 36777
rect 7561 36768 7573 36771
rect 5491 36740 7573 36768
rect 5491 36737 5503 36740
rect 5445 36731 5503 36737
rect 7561 36737 7573 36740
rect 7607 36737 7619 36771
rect 7561 36731 7619 36737
rect 7576 36700 7604 36731
rect 10870 36728 10876 36780
rect 10928 36728 10934 36780
rect 11790 36728 11796 36780
rect 11848 36728 11854 36780
rect 12069 36771 12127 36777
rect 12069 36737 12081 36771
rect 12115 36768 12127 36771
rect 14921 36771 14979 36777
rect 14921 36768 14933 36771
rect 12115 36740 14933 36768
rect 12115 36737 12127 36740
rect 12069 36731 12127 36737
rect 14921 36737 14933 36740
rect 14967 36737 14979 36771
rect 14921 36731 14979 36737
rect 11609 36703 11667 36709
rect 11609 36700 11621 36703
rect 7576 36672 11621 36700
rect 11609 36669 11621 36672
rect 11655 36700 11667 36703
rect 12084 36700 12112 36731
rect 11655 36672 12112 36700
rect 14936 36700 14964 36731
rect 18966 36728 18972 36780
rect 19024 36728 19030 36780
rect 19245 36771 19303 36777
rect 19245 36737 19257 36771
rect 19291 36768 19303 36771
rect 22281 36771 22339 36777
rect 22281 36768 22293 36771
rect 19291 36740 22293 36768
rect 19291 36737 19303 36740
rect 19245 36731 19303 36737
rect 22281 36737 22293 36740
rect 22327 36737 22339 36771
rect 22281 36731 22339 36737
rect 19260 36700 19288 36731
rect 14936 36672 19288 36700
rect 22296 36700 22324 36731
rect 25774 36728 25780 36780
rect 25832 36728 25838 36780
rect 29656 36777 29684 36876
rect 29822 36796 29828 36848
rect 29880 36836 29886 36848
rect 30576 36836 30604 36876
rect 33778 36864 33784 36916
rect 33836 36864 33842 36916
rect 33888 36876 36952 36904
rect 33888 36836 33916 36876
rect 36924 36836 36952 36876
rect 36998 36864 37004 36916
rect 37056 36864 37062 36916
rect 40862 36864 40868 36916
rect 40920 36864 40926 36916
rect 48222 36864 48228 36916
rect 48280 36864 48286 36916
rect 51902 36864 51908 36916
rect 51960 36864 51966 36916
rect 55582 36864 55588 36916
rect 55640 36864 55646 36916
rect 29880 36808 30420 36836
rect 30576 36808 33916 36836
rect 33980 36808 35894 36836
rect 36924 36808 55214 36836
rect 29880 36796 29886 36808
rect 25961 36771 26019 36777
rect 25961 36737 25973 36771
rect 26007 36768 26019 36771
rect 29641 36771 29699 36777
rect 29641 36768 29653 36771
rect 26007 36740 29653 36768
rect 26007 36737 26019 36740
rect 25961 36731 26019 36737
rect 29641 36737 29653 36740
rect 29687 36737 29699 36771
rect 29917 36771 29975 36777
rect 29917 36768 29929 36771
rect 29641 36731 29699 36737
rect 29840 36740 29929 36768
rect 25976 36700 26004 36731
rect 22296 36672 26004 36700
rect 11655 36669 11667 36672
rect 11609 36663 11667 36669
rect 11790 36592 11796 36644
rect 11848 36632 11854 36644
rect 29840 36641 29868 36740
rect 29917 36737 29929 36740
rect 29963 36737 29975 36771
rect 29917 36731 29975 36737
rect 30392 36709 30420 36808
rect 33980 36777 34008 36808
rect 33505 36771 33563 36777
rect 33505 36737 33517 36771
rect 33551 36737 33563 36771
rect 33505 36731 33563 36737
rect 33689 36771 33747 36777
rect 33689 36737 33701 36771
rect 33735 36768 33747 36771
rect 33965 36771 34023 36777
rect 33965 36768 33977 36771
rect 33735 36740 33977 36768
rect 33735 36737 33747 36740
rect 33689 36731 33747 36737
rect 33965 36737 33977 36740
rect 34011 36737 34023 36771
rect 33965 36731 34023 36737
rect 30377 36703 30435 36709
rect 30377 36669 30389 36703
rect 30423 36669 30435 36703
rect 30377 36663 30435 36669
rect 29825 36635 29883 36641
rect 11848 36604 26234 36632
rect 11848 36592 11854 36604
rect 26206 36564 26234 36604
rect 29825 36601 29837 36635
rect 29871 36601 29883 36635
rect 29825 36595 29883 36601
rect 33520 36564 33548 36731
rect 35434 36728 35440 36780
rect 35492 36728 35498 36780
rect 35866 36768 35894 36808
rect 37185 36771 37243 36777
rect 37185 36768 37197 36771
rect 35866 36740 37197 36768
rect 37185 36737 37197 36740
rect 37231 36768 37243 36771
rect 40681 36771 40739 36777
rect 40681 36768 40693 36771
rect 37231 36740 40693 36768
rect 37231 36737 37243 36740
rect 37185 36731 37243 36737
rect 40681 36737 40693 36740
rect 40727 36768 40739 36771
rect 44361 36771 44419 36777
rect 44361 36768 44373 36771
rect 40727 36740 44373 36768
rect 40727 36737 40739 36740
rect 40681 36731 40739 36737
rect 44361 36737 44373 36740
rect 44407 36737 44419 36771
rect 44637 36771 44695 36777
rect 44637 36768 44649 36771
rect 44361 36731 44419 36737
rect 44560 36740 44649 36768
rect 35342 36660 35348 36712
rect 35400 36700 35406 36712
rect 35897 36703 35955 36709
rect 35897 36700 35909 36703
rect 35400 36672 35909 36700
rect 35400 36660 35406 36672
rect 35897 36669 35909 36672
rect 35943 36669 35955 36703
rect 35897 36663 35955 36669
rect 26206 36536 33548 36564
rect 44376 36564 44404 36731
rect 44560 36641 44588 36740
rect 44637 36737 44649 36740
rect 44683 36737 44695 36771
rect 44637 36731 44695 36737
rect 48041 36771 48099 36777
rect 48041 36737 48053 36771
rect 48087 36737 48099 36771
rect 48041 36731 48099 36737
rect 44726 36660 44732 36712
rect 44784 36700 44790 36712
rect 45097 36703 45155 36709
rect 45097 36700 45109 36703
rect 44784 36672 45109 36700
rect 44784 36660 44790 36672
rect 45097 36669 45109 36672
rect 45143 36669 45155 36703
rect 45097 36663 45155 36669
rect 44545 36635 44603 36641
rect 44545 36601 44557 36635
rect 44591 36601 44603 36635
rect 48056 36632 48084 36731
rect 50154 36728 50160 36780
rect 50212 36728 50218 36780
rect 51721 36771 51779 36777
rect 51721 36737 51733 36771
rect 51767 36737 51779 36771
rect 55186 36768 55214 36808
rect 59262 36796 59268 36848
rect 59320 36836 59326 36848
rect 59320 36808 59860 36836
rect 59320 36796 59326 36808
rect 55401 36771 55459 36777
rect 55401 36768 55413 36771
rect 55186 36740 55413 36768
rect 51721 36731 51779 36737
rect 55401 36737 55413 36740
rect 55447 36768 55459 36771
rect 58437 36771 58495 36777
rect 58437 36768 58449 36771
rect 55447 36740 58449 36768
rect 55447 36737 55459 36740
rect 55401 36731 55459 36737
rect 58437 36737 58449 36740
rect 58483 36737 58495 36771
rect 58437 36731 58495 36737
rect 59357 36771 59415 36777
rect 59357 36737 59369 36771
rect 59403 36737 59415 36771
rect 59357 36731 59415 36737
rect 50062 36660 50068 36712
rect 50120 36700 50126 36712
rect 50617 36703 50675 36709
rect 50617 36700 50629 36703
rect 50120 36672 50629 36700
rect 50120 36660 50126 36672
rect 50617 36669 50629 36672
rect 50663 36669 50675 36703
rect 50617 36663 50675 36669
rect 51736 36632 51764 36731
rect 44545 36595 44603 36601
rect 45526 36604 51764 36632
rect 58621 36635 58679 36641
rect 45526 36564 45554 36604
rect 58621 36601 58633 36635
rect 58667 36632 58679 36635
rect 59372 36632 59400 36731
rect 59832 36709 59860 36808
rect 59817 36703 59875 36709
rect 59817 36669 59829 36703
rect 59863 36669 59875 36703
rect 59817 36663 59875 36669
rect 58667 36604 59400 36632
rect 58667 36601 58679 36604
rect 58621 36595 58679 36601
rect 44376 36536 45554 36564
rect 2024 36474 77924 36496
rect 2024 36422 5134 36474
rect 5186 36422 5198 36474
rect 5250 36422 5262 36474
rect 5314 36422 5326 36474
rect 5378 36422 5390 36474
rect 5442 36422 35854 36474
rect 35906 36422 35918 36474
rect 35970 36422 35982 36474
rect 36034 36422 36046 36474
rect 36098 36422 36110 36474
rect 36162 36422 66574 36474
rect 66626 36422 66638 36474
rect 66690 36422 66702 36474
rect 66754 36422 66766 36474
rect 66818 36422 66830 36474
rect 66882 36422 77924 36474
rect 2024 36400 77924 36422
rect 2024 35930 77924 35952
rect 2024 35878 5794 35930
rect 5846 35878 5858 35930
rect 5910 35878 5922 35930
rect 5974 35878 5986 35930
rect 6038 35878 6050 35930
rect 6102 35878 36514 35930
rect 36566 35878 36578 35930
rect 36630 35878 36642 35930
rect 36694 35878 36706 35930
rect 36758 35878 36770 35930
rect 36822 35878 67234 35930
rect 67286 35878 67298 35930
rect 67350 35878 67362 35930
rect 67414 35878 67426 35930
rect 67478 35878 67490 35930
rect 67542 35878 77924 35930
rect 2024 35856 77924 35878
rect 2024 35386 77924 35408
rect 2024 35334 5134 35386
rect 5186 35334 5198 35386
rect 5250 35334 5262 35386
rect 5314 35334 5326 35386
rect 5378 35334 5390 35386
rect 5442 35334 35854 35386
rect 35906 35334 35918 35386
rect 35970 35334 35982 35386
rect 36034 35334 36046 35386
rect 36098 35334 36110 35386
rect 36162 35334 66574 35386
rect 66626 35334 66638 35386
rect 66690 35334 66702 35386
rect 66754 35334 66766 35386
rect 66818 35334 66830 35386
rect 66882 35334 77924 35386
rect 2024 35312 77924 35334
rect 2024 34842 77924 34864
rect 2024 34790 5794 34842
rect 5846 34790 5858 34842
rect 5910 34790 5922 34842
rect 5974 34790 5986 34842
rect 6038 34790 6050 34842
rect 6102 34790 36514 34842
rect 36566 34790 36578 34842
rect 36630 34790 36642 34842
rect 36694 34790 36706 34842
rect 36758 34790 36770 34842
rect 36822 34790 67234 34842
rect 67286 34790 67298 34842
rect 67350 34790 67362 34842
rect 67414 34790 67426 34842
rect 67478 34790 67490 34842
rect 67542 34790 77924 34842
rect 2024 34768 77924 34790
rect 2024 34298 77924 34320
rect 2024 34246 5134 34298
rect 5186 34246 5198 34298
rect 5250 34246 5262 34298
rect 5314 34246 5326 34298
rect 5378 34246 5390 34298
rect 5442 34246 35854 34298
rect 35906 34246 35918 34298
rect 35970 34246 35982 34298
rect 36034 34246 36046 34298
rect 36098 34246 36110 34298
rect 36162 34246 66574 34298
rect 66626 34246 66638 34298
rect 66690 34246 66702 34298
rect 66754 34246 66766 34298
rect 66818 34246 66830 34298
rect 66882 34246 77924 34298
rect 2024 34224 77924 34246
rect 2024 33754 77924 33776
rect 2024 33702 5794 33754
rect 5846 33702 5858 33754
rect 5910 33702 5922 33754
rect 5974 33702 5986 33754
rect 6038 33702 6050 33754
rect 6102 33702 36514 33754
rect 36566 33702 36578 33754
rect 36630 33702 36642 33754
rect 36694 33702 36706 33754
rect 36758 33702 36770 33754
rect 36822 33702 67234 33754
rect 67286 33702 67298 33754
rect 67350 33702 67362 33754
rect 67414 33702 67426 33754
rect 67478 33702 67490 33754
rect 67542 33702 77924 33754
rect 2024 33680 77924 33702
rect 2024 33210 77924 33232
rect 2024 33158 5134 33210
rect 5186 33158 5198 33210
rect 5250 33158 5262 33210
rect 5314 33158 5326 33210
rect 5378 33158 5390 33210
rect 5442 33158 35854 33210
rect 35906 33158 35918 33210
rect 35970 33158 35982 33210
rect 36034 33158 36046 33210
rect 36098 33158 36110 33210
rect 36162 33158 66574 33210
rect 66626 33158 66638 33210
rect 66690 33158 66702 33210
rect 66754 33158 66766 33210
rect 66818 33158 66830 33210
rect 66882 33158 77924 33210
rect 2024 33136 77924 33158
rect 25774 33056 25780 33108
rect 25832 33096 25838 33108
rect 27338 33096 27344 33108
rect 25832 33068 27344 33096
rect 25832 33056 25838 33068
rect 27338 33056 27344 33068
rect 27396 33056 27402 33108
rect 2024 32666 77924 32688
rect 2024 32614 5794 32666
rect 5846 32614 5858 32666
rect 5910 32614 5922 32666
rect 5974 32614 5986 32666
rect 6038 32614 6050 32666
rect 6102 32614 36514 32666
rect 36566 32614 36578 32666
rect 36630 32614 36642 32666
rect 36694 32614 36706 32666
rect 36758 32614 36770 32666
rect 36822 32614 67234 32666
rect 67286 32614 67298 32666
rect 67350 32614 67362 32666
rect 67414 32614 67426 32666
rect 67478 32614 67490 32666
rect 67542 32614 77924 32666
rect 2024 32592 77924 32614
rect 26326 32376 26332 32428
rect 26384 32416 26390 32428
rect 43346 32416 43352 32428
rect 26384 32388 43352 32416
rect 26384 32376 26390 32388
rect 43346 32376 43352 32388
rect 43404 32376 43410 32428
rect 2024 32122 77924 32144
rect 2024 32070 5134 32122
rect 5186 32070 5198 32122
rect 5250 32070 5262 32122
rect 5314 32070 5326 32122
rect 5378 32070 5390 32122
rect 5442 32070 35854 32122
rect 35906 32070 35918 32122
rect 35970 32070 35982 32122
rect 36034 32070 36046 32122
rect 36098 32070 36110 32122
rect 36162 32070 66574 32122
rect 66626 32070 66638 32122
rect 66690 32070 66702 32122
rect 66754 32070 66766 32122
rect 66818 32070 66830 32122
rect 66882 32070 77924 32122
rect 2024 32048 77924 32070
rect 2024 31578 77924 31600
rect 2024 31526 5794 31578
rect 5846 31526 5858 31578
rect 5910 31526 5922 31578
rect 5974 31526 5986 31578
rect 6038 31526 6050 31578
rect 6102 31526 36514 31578
rect 36566 31526 36578 31578
rect 36630 31526 36642 31578
rect 36694 31526 36706 31578
rect 36758 31526 36770 31578
rect 36822 31526 67234 31578
rect 67286 31526 67298 31578
rect 67350 31526 67362 31578
rect 67414 31526 67426 31578
rect 67478 31526 67490 31578
rect 67542 31526 77924 31578
rect 2024 31504 77924 31526
rect 2024 31034 77924 31056
rect 2024 30982 5134 31034
rect 5186 30982 5198 31034
rect 5250 30982 5262 31034
rect 5314 30982 5326 31034
rect 5378 30982 5390 31034
rect 5442 30982 35854 31034
rect 35906 30982 35918 31034
rect 35970 30982 35982 31034
rect 36034 30982 36046 31034
rect 36098 30982 36110 31034
rect 36162 30982 66574 31034
rect 66626 30982 66638 31034
rect 66690 30982 66702 31034
rect 66754 30982 66766 31034
rect 66818 30982 66830 31034
rect 66882 30982 77924 31034
rect 2024 30960 77924 30982
rect 2024 30490 77924 30512
rect 2024 30438 5794 30490
rect 5846 30438 5858 30490
rect 5910 30438 5922 30490
rect 5974 30438 5986 30490
rect 6038 30438 6050 30490
rect 6102 30438 36514 30490
rect 36566 30438 36578 30490
rect 36630 30438 36642 30490
rect 36694 30438 36706 30490
rect 36758 30438 36770 30490
rect 36822 30438 67234 30490
rect 67286 30438 67298 30490
rect 67350 30438 67362 30490
rect 67414 30438 67426 30490
rect 67478 30438 67490 30490
rect 67542 30438 77924 30490
rect 2024 30416 77924 30438
rect 2024 29946 77924 29968
rect 2024 29894 5134 29946
rect 5186 29894 5198 29946
rect 5250 29894 5262 29946
rect 5314 29894 5326 29946
rect 5378 29894 5390 29946
rect 5442 29894 35854 29946
rect 35906 29894 35918 29946
rect 35970 29894 35982 29946
rect 36034 29894 36046 29946
rect 36098 29894 36110 29946
rect 36162 29894 66574 29946
rect 66626 29894 66638 29946
rect 66690 29894 66702 29946
rect 66754 29894 66766 29946
rect 66818 29894 66830 29946
rect 66882 29894 77924 29946
rect 2024 29872 77924 29894
rect 26050 29588 26056 29640
rect 26108 29628 26114 29640
rect 50154 29628 50160 29640
rect 26108 29600 50160 29628
rect 26108 29588 26114 29600
rect 50154 29588 50160 29600
rect 50212 29588 50218 29640
rect 2024 29402 77924 29424
rect 2024 29350 5794 29402
rect 5846 29350 5858 29402
rect 5910 29350 5922 29402
rect 5974 29350 5986 29402
rect 6038 29350 6050 29402
rect 6102 29350 36514 29402
rect 36566 29350 36578 29402
rect 36630 29350 36642 29402
rect 36694 29350 36706 29402
rect 36758 29350 36770 29402
rect 36822 29350 67234 29402
rect 67286 29350 67298 29402
rect 67350 29350 67362 29402
rect 67414 29350 67426 29402
rect 67478 29350 67490 29402
rect 67542 29350 77924 29402
rect 2024 29328 77924 29350
rect 2024 28858 77924 28880
rect 2024 28806 5134 28858
rect 5186 28806 5198 28858
rect 5250 28806 5262 28858
rect 5314 28806 5326 28858
rect 5378 28806 5390 28858
rect 5442 28806 35854 28858
rect 35906 28806 35918 28858
rect 35970 28806 35982 28858
rect 36034 28806 36046 28858
rect 36098 28806 36110 28858
rect 36162 28806 66574 28858
rect 66626 28806 66638 28858
rect 66690 28806 66702 28858
rect 66754 28806 66766 28858
rect 66818 28806 66830 28858
rect 66882 28806 77924 28858
rect 2024 28784 77924 28806
rect 2024 28314 77924 28336
rect 2024 28262 5794 28314
rect 5846 28262 5858 28314
rect 5910 28262 5922 28314
rect 5974 28262 5986 28314
rect 6038 28262 6050 28314
rect 6102 28262 36514 28314
rect 36566 28262 36578 28314
rect 36630 28262 36642 28314
rect 36694 28262 36706 28314
rect 36758 28262 36770 28314
rect 36822 28262 67234 28314
rect 67286 28262 67298 28314
rect 67350 28262 67362 28314
rect 67414 28262 67426 28314
rect 67478 28262 67490 28314
rect 67542 28262 77924 28314
rect 2024 28240 77924 28262
rect 2024 27770 77924 27792
rect 2024 27718 5134 27770
rect 5186 27718 5198 27770
rect 5250 27718 5262 27770
rect 5314 27718 5326 27770
rect 5378 27718 5390 27770
rect 5442 27718 35854 27770
rect 35906 27718 35918 27770
rect 35970 27718 35982 27770
rect 36034 27718 36046 27770
rect 36098 27718 36110 27770
rect 36162 27718 66574 27770
rect 66626 27718 66638 27770
rect 66690 27718 66702 27770
rect 66754 27718 66766 27770
rect 66818 27718 66830 27770
rect 66882 27718 77924 27770
rect 2024 27696 77924 27718
rect 2024 27226 77924 27248
rect 2024 27174 5794 27226
rect 5846 27174 5858 27226
rect 5910 27174 5922 27226
rect 5974 27174 5986 27226
rect 6038 27174 6050 27226
rect 6102 27174 36514 27226
rect 36566 27174 36578 27226
rect 36630 27174 36642 27226
rect 36694 27174 36706 27226
rect 36758 27174 36770 27226
rect 36822 27174 67234 27226
rect 67286 27174 67298 27226
rect 67350 27174 67362 27226
rect 67414 27174 67426 27226
rect 67478 27174 67490 27226
rect 67542 27174 77924 27226
rect 2024 27152 77924 27174
rect 25682 26868 25688 26920
rect 25740 26908 25746 26920
rect 53834 26908 53840 26920
rect 25740 26880 53840 26908
rect 25740 26868 25746 26880
rect 53834 26868 53840 26880
rect 53892 26868 53898 26920
rect 2024 26682 77924 26704
rect 2024 26630 5134 26682
rect 5186 26630 5198 26682
rect 5250 26630 5262 26682
rect 5314 26630 5326 26682
rect 5378 26630 5390 26682
rect 5442 26630 35854 26682
rect 35906 26630 35918 26682
rect 35970 26630 35982 26682
rect 36034 26630 36046 26682
rect 36098 26630 36110 26682
rect 36162 26630 66574 26682
rect 66626 26630 66638 26682
rect 66690 26630 66702 26682
rect 66754 26630 66766 26682
rect 66818 26630 66830 26682
rect 66882 26630 77924 26682
rect 2024 26608 77924 26630
rect 2024 26138 77924 26160
rect 2024 26086 5794 26138
rect 5846 26086 5858 26138
rect 5910 26086 5922 26138
rect 5974 26086 5986 26138
rect 6038 26086 6050 26138
rect 6102 26086 36514 26138
rect 36566 26086 36578 26138
rect 36630 26086 36642 26138
rect 36694 26086 36706 26138
rect 36758 26086 36770 26138
rect 36822 26086 67234 26138
rect 67286 26086 67298 26138
rect 67350 26086 67362 26138
rect 67414 26086 67426 26138
rect 67478 26086 67490 26138
rect 67542 26086 77924 26138
rect 2024 26064 77924 26086
rect 2024 25594 77924 25616
rect 2024 25542 5134 25594
rect 5186 25542 5198 25594
rect 5250 25542 5262 25594
rect 5314 25542 5326 25594
rect 5378 25542 5390 25594
rect 5442 25542 35854 25594
rect 35906 25542 35918 25594
rect 35970 25542 35982 25594
rect 36034 25542 36046 25594
rect 36098 25542 36110 25594
rect 36162 25542 66574 25594
rect 66626 25542 66638 25594
rect 66690 25542 66702 25594
rect 66754 25542 66766 25594
rect 66818 25542 66830 25594
rect 66882 25542 77924 25594
rect 2024 25520 77924 25542
rect 2024 25050 77924 25072
rect 2024 24998 5794 25050
rect 5846 24998 5858 25050
rect 5910 24998 5922 25050
rect 5974 24998 5986 25050
rect 6038 24998 6050 25050
rect 6102 24998 36514 25050
rect 36566 24998 36578 25050
rect 36630 24998 36642 25050
rect 36694 24998 36706 25050
rect 36758 24998 36770 25050
rect 36822 24998 67234 25050
rect 67286 24998 67298 25050
rect 67350 24998 67362 25050
rect 67414 24998 67426 25050
rect 67478 24998 67490 25050
rect 67542 24998 77924 25050
rect 2024 24976 77924 24998
rect 2024 24506 77924 24528
rect 2024 24454 5134 24506
rect 5186 24454 5198 24506
rect 5250 24454 5262 24506
rect 5314 24454 5326 24506
rect 5378 24454 5390 24506
rect 5442 24454 35854 24506
rect 35906 24454 35918 24506
rect 35970 24454 35982 24506
rect 36034 24454 36046 24506
rect 36098 24454 36110 24506
rect 36162 24454 66574 24506
rect 66626 24454 66638 24506
rect 66690 24454 66702 24506
rect 66754 24454 66766 24506
rect 66818 24454 66830 24506
rect 66882 24454 77924 24506
rect 2024 24432 77924 24454
rect 25498 24080 25504 24132
rect 25556 24120 25562 24132
rect 46474 24120 46480 24132
rect 25556 24092 46480 24120
rect 25556 24080 25562 24092
rect 46474 24080 46480 24092
rect 46532 24080 46538 24132
rect 2024 23962 77924 23984
rect 2024 23910 5794 23962
rect 5846 23910 5858 23962
rect 5910 23910 5922 23962
rect 5974 23910 5986 23962
rect 6038 23910 6050 23962
rect 6102 23910 36514 23962
rect 36566 23910 36578 23962
rect 36630 23910 36642 23962
rect 36694 23910 36706 23962
rect 36758 23910 36770 23962
rect 36822 23910 67234 23962
rect 67286 23910 67298 23962
rect 67350 23910 67362 23962
rect 67414 23910 67426 23962
rect 67478 23910 67490 23962
rect 67542 23910 77924 23962
rect 2024 23888 77924 23910
rect 2024 23418 77924 23440
rect 2024 23366 5134 23418
rect 5186 23366 5198 23418
rect 5250 23366 5262 23418
rect 5314 23366 5326 23418
rect 5378 23366 5390 23418
rect 5442 23366 35854 23418
rect 35906 23366 35918 23418
rect 35970 23366 35982 23418
rect 36034 23366 36046 23418
rect 36098 23366 36110 23418
rect 36162 23366 66574 23418
rect 66626 23366 66638 23418
rect 66690 23366 66702 23418
rect 66754 23366 66766 23418
rect 66818 23366 66830 23418
rect 66882 23366 77924 23418
rect 2024 23344 77924 23366
rect 2024 22874 77924 22896
rect 2024 22822 5794 22874
rect 5846 22822 5858 22874
rect 5910 22822 5922 22874
rect 5974 22822 5986 22874
rect 6038 22822 6050 22874
rect 6102 22822 36514 22874
rect 36566 22822 36578 22874
rect 36630 22822 36642 22874
rect 36694 22822 36706 22874
rect 36758 22822 36770 22874
rect 36822 22822 67234 22874
rect 67286 22822 67298 22874
rect 67350 22822 67362 22874
rect 67414 22822 67426 22874
rect 67478 22822 67490 22874
rect 67542 22822 77924 22874
rect 2024 22800 77924 22822
rect 2024 22330 77924 22352
rect 2024 22278 5134 22330
rect 5186 22278 5198 22330
rect 5250 22278 5262 22330
rect 5314 22278 5326 22330
rect 5378 22278 5390 22330
rect 5442 22278 35854 22330
rect 35906 22278 35918 22330
rect 35970 22278 35982 22330
rect 36034 22278 36046 22330
rect 36098 22278 36110 22330
rect 36162 22278 66574 22330
rect 66626 22278 66638 22330
rect 66690 22278 66702 22330
rect 66754 22278 66766 22330
rect 66818 22278 66830 22330
rect 66882 22278 77924 22330
rect 2024 22256 77924 22278
rect 2024 21786 77924 21808
rect 2024 21734 5794 21786
rect 5846 21734 5858 21786
rect 5910 21734 5922 21786
rect 5974 21734 5986 21786
rect 6038 21734 6050 21786
rect 6102 21734 36514 21786
rect 36566 21734 36578 21786
rect 36630 21734 36642 21786
rect 36694 21734 36706 21786
rect 36758 21734 36770 21786
rect 36822 21734 67234 21786
rect 67286 21734 67298 21786
rect 67350 21734 67362 21786
rect 67414 21734 67426 21786
rect 67478 21734 67490 21786
rect 67542 21734 77924 21786
rect 2024 21712 77924 21734
rect 2024 21242 77924 21264
rect 2024 21190 5134 21242
rect 5186 21190 5198 21242
rect 5250 21190 5262 21242
rect 5314 21190 5326 21242
rect 5378 21190 5390 21242
rect 5442 21190 35854 21242
rect 35906 21190 35918 21242
rect 35970 21190 35982 21242
rect 36034 21190 36046 21242
rect 36098 21190 36110 21242
rect 36162 21190 66574 21242
rect 66626 21190 66638 21242
rect 66690 21190 66702 21242
rect 66754 21190 66766 21242
rect 66818 21190 66830 21242
rect 66882 21190 77924 21242
rect 2024 21168 77924 21190
rect 2024 20698 77924 20720
rect 2024 20646 5794 20698
rect 5846 20646 5858 20698
rect 5910 20646 5922 20698
rect 5974 20646 5986 20698
rect 6038 20646 6050 20698
rect 6102 20646 36514 20698
rect 36566 20646 36578 20698
rect 36630 20646 36642 20698
rect 36694 20646 36706 20698
rect 36758 20646 36770 20698
rect 36822 20646 67234 20698
rect 67286 20646 67298 20698
rect 67350 20646 67362 20698
rect 67414 20646 67426 20698
rect 67478 20646 67490 20698
rect 67542 20646 77924 20698
rect 2024 20624 77924 20646
rect 2024 20154 77924 20176
rect 2024 20102 5134 20154
rect 5186 20102 5198 20154
rect 5250 20102 5262 20154
rect 5314 20102 5326 20154
rect 5378 20102 5390 20154
rect 5442 20102 35854 20154
rect 35906 20102 35918 20154
rect 35970 20102 35982 20154
rect 36034 20102 36046 20154
rect 36098 20102 36110 20154
rect 36162 20102 66574 20154
rect 66626 20102 66638 20154
rect 66690 20102 66702 20154
rect 66754 20102 66766 20154
rect 66818 20102 66830 20154
rect 66882 20102 77924 20154
rect 2024 20080 77924 20102
rect 2024 19610 77924 19632
rect 2024 19558 5794 19610
rect 5846 19558 5858 19610
rect 5910 19558 5922 19610
rect 5974 19558 5986 19610
rect 6038 19558 6050 19610
rect 6102 19558 36514 19610
rect 36566 19558 36578 19610
rect 36630 19558 36642 19610
rect 36694 19558 36706 19610
rect 36758 19558 36770 19610
rect 36822 19558 67234 19610
rect 67286 19558 67298 19610
rect 67350 19558 67362 19610
rect 67414 19558 67426 19610
rect 67478 19558 67490 19610
rect 67542 19558 77924 19610
rect 2024 19536 77924 19558
rect 2024 19066 77924 19088
rect 2024 19014 5134 19066
rect 5186 19014 5198 19066
rect 5250 19014 5262 19066
rect 5314 19014 5326 19066
rect 5378 19014 5390 19066
rect 5442 19014 35854 19066
rect 35906 19014 35918 19066
rect 35970 19014 35982 19066
rect 36034 19014 36046 19066
rect 36098 19014 36110 19066
rect 36162 19014 66574 19066
rect 66626 19014 66638 19066
rect 66690 19014 66702 19066
rect 66754 19014 66766 19066
rect 66818 19014 66830 19066
rect 66882 19014 77924 19066
rect 2024 18992 77924 19014
rect 2024 18522 77924 18544
rect 2024 18470 5794 18522
rect 5846 18470 5858 18522
rect 5910 18470 5922 18522
rect 5974 18470 5986 18522
rect 6038 18470 6050 18522
rect 6102 18470 36514 18522
rect 36566 18470 36578 18522
rect 36630 18470 36642 18522
rect 36694 18470 36706 18522
rect 36758 18470 36770 18522
rect 36822 18470 67234 18522
rect 67286 18470 67298 18522
rect 67350 18470 67362 18522
rect 67414 18470 67426 18522
rect 67478 18470 67490 18522
rect 67542 18470 77924 18522
rect 2024 18448 77924 18470
rect 2024 17978 77924 18000
rect 2024 17926 5134 17978
rect 5186 17926 5198 17978
rect 5250 17926 5262 17978
rect 5314 17926 5326 17978
rect 5378 17926 5390 17978
rect 5442 17926 35854 17978
rect 35906 17926 35918 17978
rect 35970 17926 35982 17978
rect 36034 17926 36046 17978
rect 36098 17926 36110 17978
rect 36162 17926 66574 17978
rect 66626 17926 66638 17978
rect 66690 17926 66702 17978
rect 66754 17926 66766 17978
rect 66818 17926 66830 17978
rect 66882 17926 77924 17978
rect 2024 17904 77924 17926
rect 29270 17824 29276 17876
rect 29328 17864 29334 17876
rect 31110 17864 31116 17876
rect 29328 17836 31116 17864
rect 29328 17824 29334 17836
rect 31110 17824 31116 17836
rect 31168 17824 31174 17876
rect 31662 17824 31668 17876
rect 31720 17864 31726 17876
rect 35434 17864 35440 17876
rect 31720 17836 35440 17864
rect 31720 17824 31726 17836
rect 35434 17824 35440 17836
rect 35492 17824 35498 17876
rect 2024 17434 77924 17456
rect 2024 17382 5794 17434
rect 5846 17382 5858 17434
rect 5910 17382 5922 17434
rect 5974 17382 5986 17434
rect 6038 17382 6050 17434
rect 6102 17382 36514 17434
rect 36566 17382 36578 17434
rect 36630 17382 36642 17434
rect 36694 17382 36706 17434
rect 36758 17382 36770 17434
rect 36822 17382 67234 17434
rect 67286 17382 67298 17434
rect 67350 17382 67362 17434
rect 67414 17382 67426 17434
rect 67478 17382 67490 17434
rect 67542 17382 77924 17434
rect 2024 17360 77924 17382
rect 2024 16890 77924 16912
rect 2024 16838 5134 16890
rect 5186 16838 5198 16890
rect 5250 16838 5262 16890
rect 5314 16838 5326 16890
rect 5378 16838 5390 16890
rect 5442 16838 35854 16890
rect 35906 16838 35918 16890
rect 35970 16838 35982 16890
rect 36034 16838 36046 16890
rect 36098 16838 36110 16890
rect 36162 16838 66574 16890
rect 66626 16838 66638 16890
rect 66690 16838 66702 16890
rect 66754 16838 66766 16890
rect 66818 16838 66830 16890
rect 66882 16838 77924 16890
rect 2024 16816 77924 16838
rect 2024 16346 77924 16368
rect 2024 16294 5794 16346
rect 5846 16294 5858 16346
rect 5910 16294 5922 16346
rect 5974 16294 5986 16346
rect 6038 16294 6050 16346
rect 6102 16294 36514 16346
rect 36566 16294 36578 16346
rect 36630 16294 36642 16346
rect 36694 16294 36706 16346
rect 36758 16294 36770 16346
rect 36822 16294 67234 16346
rect 67286 16294 67298 16346
rect 67350 16294 67362 16346
rect 67414 16294 67426 16346
rect 67478 16294 67490 16346
rect 67542 16294 77924 16346
rect 2024 16272 77924 16294
rect 2024 15802 77924 15824
rect 2024 15750 5134 15802
rect 5186 15750 5198 15802
rect 5250 15750 5262 15802
rect 5314 15750 5326 15802
rect 5378 15750 5390 15802
rect 5442 15750 35854 15802
rect 35906 15750 35918 15802
rect 35970 15750 35982 15802
rect 36034 15750 36046 15802
rect 36098 15750 36110 15802
rect 36162 15750 66574 15802
rect 66626 15750 66638 15802
rect 66690 15750 66702 15802
rect 66754 15750 66766 15802
rect 66818 15750 66830 15802
rect 66882 15750 77924 15802
rect 2024 15728 77924 15750
rect 2024 15258 77924 15280
rect 2024 15206 5794 15258
rect 5846 15206 5858 15258
rect 5910 15206 5922 15258
rect 5974 15206 5986 15258
rect 6038 15206 6050 15258
rect 6102 15206 36514 15258
rect 36566 15206 36578 15258
rect 36630 15206 36642 15258
rect 36694 15206 36706 15258
rect 36758 15206 36770 15258
rect 36822 15206 67234 15258
rect 67286 15206 67298 15258
rect 67350 15206 67362 15258
rect 67414 15206 67426 15258
rect 67478 15206 67490 15258
rect 67542 15206 77924 15258
rect 2024 15184 77924 15206
rect 2024 14714 77924 14736
rect 2024 14662 5134 14714
rect 5186 14662 5198 14714
rect 5250 14662 5262 14714
rect 5314 14662 5326 14714
rect 5378 14662 5390 14714
rect 5442 14662 35854 14714
rect 35906 14662 35918 14714
rect 35970 14662 35982 14714
rect 36034 14662 36046 14714
rect 36098 14662 36110 14714
rect 36162 14662 66574 14714
rect 66626 14662 66638 14714
rect 66690 14662 66702 14714
rect 66754 14662 66766 14714
rect 66818 14662 66830 14714
rect 66882 14662 77924 14714
rect 2024 14640 77924 14662
rect 25958 14424 25964 14476
rect 26016 14464 26022 14476
rect 58802 14464 58808 14476
rect 26016 14436 58808 14464
rect 26016 14424 26022 14436
rect 58802 14424 58808 14436
rect 58860 14424 58866 14476
rect 2024 14170 77924 14192
rect 2024 14118 5794 14170
rect 5846 14118 5858 14170
rect 5910 14118 5922 14170
rect 5974 14118 5986 14170
rect 6038 14118 6050 14170
rect 6102 14118 36514 14170
rect 36566 14118 36578 14170
rect 36630 14118 36642 14170
rect 36694 14118 36706 14170
rect 36758 14118 36770 14170
rect 36822 14118 67234 14170
rect 67286 14118 67298 14170
rect 67350 14118 67362 14170
rect 67414 14118 67426 14170
rect 67478 14118 67490 14170
rect 67542 14118 77924 14170
rect 2024 14096 77924 14118
rect 2024 13626 77924 13648
rect 2024 13574 5134 13626
rect 5186 13574 5198 13626
rect 5250 13574 5262 13626
rect 5314 13574 5326 13626
rect 5378 13574 5390 13626
rect 5442 13574 35854 13626
rect 35906 13574 35918 13626
rect 35970 13574 35982 13626
rect 36034 13574 36046 13626
rect 36098 13574 36110 13626
rect 36162 13574 66574 13626
rect 66626 13574 66638 13626
rect 66690 13574 66702 13626
rect 66754 13574 66766 13626
rect 66818 13574 66830 13626
rect 66882 13574 77924 13626
rect 2024 13552 77924 13574
rect 2024 13082 77924 13104
rect 2024 13030 5794 13082
rect 5846 13030 5858 13082
rect 5910 13030 5922 13082
rect 5974 13030 5986 13082
rect 6038 13030 6050 13082
rect 6102 13030 36514 13082
rect 36566 13030 36578 13082
rect 36630 13030 36642 13082
rect 36694 13030 36706 13082
rect 36758 13030 36770 13082
rect 36822 13030 67234 13082
rect 67286 13030 67298 13082
rect 67350 13030 67362 13082
rect 67414 13030 67426 13082
rect 67478 13030 67490 13082
rect 67542 13030 77924 13082
rect 2024 13008 77924 13030
rect 14182 12656 14188 12708
rect 14240 12696 14246 12708
rect 27890 12696 27896 12708
rect 14240 12668 27896 12696
rect 14240 12656 14246 12668
rect 27890 12656 27896 12668
rect 27948 12656 27954 12708
rect 17586 12588 17592 12640
rect 17644 12628 17650 12640
rect 38010 12628 38016 12640
rect 17644 12600 38016 12628
rect 17644 12588 17650 12600
rect 38010 12588 38016 12600
rect 38068 12588 38074 12640
rect 2024 12538 77924 12560
rect 2024 12486 5134 12538
rect 5186 12486 5198 12538
rect 5250 12486 5262 12538
rect 5314 12486 5326 12538
rect 5378 12486 5390 12538
rect 5442 12486 35854 12538
rect 35906 12486 35918 12538
rect 35970 12486 35982 12538
rect 36034 12486 36046 12538
rect 36098 12486 36110 12538
rect 36162 12486 66574 12538
rect 66626 12486 66638 12538
rect 66690 12486 66702 12538
rect 66754 12486 66766 12538
rect 66818 12486 66830 12538
rect 66882 12486 77924 12538
rect 2024 12464 77924 12486
rect 25682 12044 25688 12096
rect 25740 12084 25746 12096
rect 30834 12084 30840 12096
rect 25740 12056 30840 12084
rect 25740 12044 25746 12056
rect 30834 12044 30840 12056
rect 30892 12044 30898 12096
rect 2024 11994 77924 12016
rect 2024 11942 5794 11994
rect 5846 11942 5858 11994
rect 5910 11942 5922 11994
rect 5974 11942 5986 11994
rect 6038 11942 6050 11994
rect 6102 11942 36514 11994
rect 36566 11942 36578 11994
rect 36630 11942 36642 11994
rect 36694 11942 36706 11994
rect 36758 11942 36770 11994
rect 36822 11942 67234 11994
rect 67286 11942 67298 11994
rect 67350 11942 67362 11994
rect 67414 11942 67426 11994
rect 67478 11942 67490 11994
rect 67542 11942 77924 11994
rect 2024 11920 77924 11942
rect 23106 11840 23112 11892
rect 23164 11880 23170 11892
rect 25314 11880 25320 11892
rect 23164 11852 25320 11880
rect 23164 11840 23170 11852
rect 25314 11840 25320 11852
rect 25372 11840 25378 11892
rect 36354 11880 36360 11892
rect 29104 11852 36360 11880
rect 22186 11772 22192 11824
rect 22244 11812 22250 11824
rect 27062 11812 27068 11824
rect 22244 11784 27068 11812
rect 22244 11772 22250 11784
rect 27062 11772 27068 11784
rect 27120 11772 27126 11824
rect 28074 11772 28080 11824
rect 28132 11812 28138 11824
rect 28721 11815 28779 11821
rect 28721 11812 28733 11815
rect 28132 11784 28733 11812
rect 28132 11772 28138 11784
rect 28721 11781 28733 11784
rect 28767 11781 28779 11815
rect 28721 11775 28779 11781
rect 24302 11704 24308 11756
rect 24360 11744 24366 11756
rect 24762 11744 24768 11756
rect 24360 11716 24768 11744
rect 24360 11704 24366 11716
rect 24762 11704 24768 11716
rect 24820 11744 24826 11756
rect 26234 11744 26240 11756
rect 24820 11716 26240 11744
rect 24820 11704 24826 11716
rect 26234 11704 26240 11716
rect 26292 11704 26298 11756
rect 29104 11753 29132 11852
rect 36354 11840 36360 11852
rect 36412 11840 36418 11892
rect 30282 11812 30288 11824
rect 29472 11784 30288 11812
rect 29472 11753 29500 11784
rect 30282 11772 30288 11784
rect 30340 11772 30346 11824
rect 29089 11747 29147 11753
rect 29089 11744 29101 11747
rect 28552 11716 29101 11744
rect 19426 11636 19432 11688
rect 19484 11676 19490 11688
rect 23934 11676 23940 11688
rect 19484 11648 23940 11676
rect 19484 11636 19490 11648
rect 23934 11636 23940 11648
rect 23992 11676 23998 11688
rect 27246 11676 27252 11688
rect 23992 11648 27252 11676
rect 23992 11636 23998 11648
rect 27246 11636 27252 11648
rect 27304 11636 27310 11688
rect 21910 11568 21916 11620
rect 21968 11608 21974 11620
rect 24854 11608 24860 11620
rect 21968 11580 24860 11608
rect 21968 11568 21974 11580
rect 24854 11568 24860 11580
rect 24912 11608 24918 11620
rect 25958 11608 25964 11620
rect 24912 11580 25964 11608
rect 24912 11568 24918 11580
rect 25958 11568 25964 11580
rect 26016 11568 26022 11620
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 28552 11549 28580 11716
rect 29089 11713 29101 11716
rect 29135 11713 29147 11747
rect 29089 11707 29147 11713
rect 29457 11747 29515 11753
rect 29457 11713 29469 11747
rect 29503 11713 29515 11747
rect 29457 11707 29515 11713
rect 29638 11704 29644 11756
rect 29696 11704 29702 11756
rect 29733 11747 29791 11753
rect 29733 11713 29745 11747
rect 29779 11713 29791 11747
rect 29733 11707 29791 11713
rect 28902 11636 28908 11688
rect 28960 11676 28966 11688
rect 29748 11676 29776 11707
rect 28960 11648 29776 11676
rect 28960 11636 28966 11648
rect 28994 11568 29000 11620
rect 29052 11608 29058 11620
rect 38838 11608 38844 11620
rect 29052 11580 38844 11608
rect 29052 11568 29058 11580
rect 38838 11568 38844 11580
rect 38896 11568 38902 11620
rect 28537 11543 28595 11549
rect 28537 11540 28549 11543
rect 13044 11512 28549 11540
rect 13044 11500 13050 11512
rect 28537 11509 28549 11512
rect 28583 11509 28595 11543
rect 28537 11503 28595 11509
rect 29270 11500 29276 11552
rect 29328 11500 29334 11552
rect 2024 11450 77924 11472
rect 2024 11398 5134 11450
rect 5186 11398 5198 11450
rect 5250 11398 5262 11450
rect 5314 11398 5326 11450
rect 5378 11398 5390 11450
rect 5442 11398 35854 11450
rect 35906 11398 35918 11450
rect 35970 11398 35982 11450
rect 36034 11398 36046 11450
rect 36098 11398 36110 11450
rect 36162 11398 66574 11450
rect 66626 11398 66638 11450
rect 66690 11398 66702 11450
rect 66754 11398 66766 11450
rect 66818 11398 66830 11450
rect 66882 11398 77924 11450
rect 2024 11376 77924 11398
rect 20346 11296 20352 11348
rect 20404 11336 20410 11348
rect 24213 11339 24271 11345
rect 24213 11336 24225 11339
rect 20404 11308 24225 11336
rect 20404 11296 20410 11308
rect 24213 11305 24225 11308
rect 24259 11305 24271 11339
rect 24670 11336 24676 11348
rect 24213 11299 24271 11305
rect 24320 11308 24676 11336
rect 22094 11228 22100 11280
rect 22152 11228 22158 11280
rect 22281 11271 22339 11277
rect 22281 11268 22293 11271
rect 22204 11240 22293 11268
rect 16574 11160 16580 11212
rect 16632 11200 16638 11212
rect 22204 11200 22232 11240
rect 22281 11237 22293 11240
rect 22327 11237 22339 11271
rect 22281 11231 22339 11237
rect 22741 11271 22799 11277
rect 22741 11237 22753 11271
rect 22787 11268 22799 11271
rect 23382 11268 23388 11280
rect 22787 11240 23388 11268
rect 22787 11237 22799 11240
rect 22741 11231 22799 11237
rect 23382 11228 23388 11240
rect 23440 11228 23446 11280
rect 23474 11228 23480 11280
rect 23532 11228 23538 11280
rect 24320 11268 24348 11308
rect 24670 11296 24676 11308
rect 24728 11296 24734 11348
rect 26970 11336 26976 11348
rect 25424 11308 26976 11336
rect 23584 11240 24348 11268
rect 23584 11200 23612 11240
rect 16632 11172 22232 11200
rect 22388 11172 23612 11200
rect 23845 11203 23903 11209
rect 16632 11160 16638 11172
rect 20806 11092 20812 11144
rect 20864 11132 20870 11144
rect 21910 11132 21916 11144
rect 20864 11104 21916 11132
rect 20864 11092 20870 11104
rect 21910 11092 21916 11104
rect 21968 11092 21974 11144
rect 22005 11135 22063 11141
rect 22005 11101 22017 11135
rect 22051 11132 22063 11135
rect 22388 11132 22416 11172
rect 23845 11169 23857 11203
rect 23891 11200 23903 11203
rect 24486 11200 24492 11212
rect 23891 11172 24492 11200
rect 23891 11169 23903 11172
rect 23845 11163 23903 11169
rect 24486 11160 24492 11172
rect 24544 11160 24550 11212
rect 24854 11200 24860 11212
rect 24596 11172 24860 11200
rect 22051 11104 22416 11132
rect 22051 11101 22063 11104
rect 22005 11095 22063 11101
rect 22462 11092 22468 11144
rect 22520 11092 22526 11144
rect 22554 11092 22560 11144
rect 22612 11132 22618 11144
rect 23661 11135 23719 11141
rect 23661 11132 23673 11135
rect 22612 11104 23673 11132
rect 22612 11092 22618 11104
rect 23661 11101 23673 11104
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 23934 11092 23940 11144
rect 23992 11092 23998 11144
rect 24596 11141 24624 11172
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 25424 11209 25452 11308
rect 26970 11296 26976 11308
rect 27028 11296 27034 11348
rect 27430 11296 27436 11348
rect 27488 11336 27494 11348
rect 28445 11339 28503 11345
rect 28445 11336 28457 11339
rect 27488 11308 28457 11336
rect 27488 11296 27494 11308
rect 28445 11305 28457 11308
rect 28491 11305 28503 11339
rect 28445 11299 28503 11305
rect 28813 11339 28871 11345
rect 28813 11305 28825 11339
rect 28859 11336 28871 11339
rect 28994 11336 29000 11348
rect 28859 11308 29000 11336
rect 28859 11305 28871 11308
rect 28813 11299 28871 11305
rect 28994 11296 29000 11308
rect 29052 11296 29058 11348
rect 27982 11228 27988 11280
rect 28040 11268 28046 11280
rect 28307 11271 28365 11277
rect 28307 11268 28319 11271
rect 28040 11240 28319 11268
rect 28040 11228 28046 11240
rect 28307 11237 28319 11240
rect 28353 11237 28365 11271
rect 30374 11268 30380 11280
rect 28307 11231 28365 11237
rect 28460 11240 30380 11268
rect 25409 11203 25467 11209
rect 25409 11169 25421 11203
rect 25455 11169 25467 11203
rect 25409 11163 25467 11169
rect 25593 11203 25651 11209
rect 25593 11169 25605 11203
rect 25639 11200 25651 11203
rect 28460 11200 28488 11240
rect 30374 11228 30380 11240
rect 30432 11228 30438 11280
rect 25639 11172 28488 11200
rect 25639 11169 25651 11172
rect 25593 11163 25651 11169
rect 28534 11160 28540 11212
rect 28592 11160 28598 11212
rect 28718 11160 28724 11212
rect 28776 11200 28782 11212
rect 29641 11203 29699 11209
rect 29641 11200 29653 11203
rect 28776 11172 29653 11200
rect 28776 11160 28782 11172
rect 29641 11169 29653 11172
rect 29687 11169 29699 11203
rect 29641 11163 29699 11169
rect 24121 11135 24179 11141
rect 24121 11101 24133 11135
rect 24167 11132 24179 11135
rect 24397 11135 24455 11141
rect 24397 11132 24409 11135
rect 24167 11104 24409 11132
rect 24167 11101 24179 11104
rect 24121 11095 24179 11101
rect 24397 11101 24409 11104
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 20254 11024 20260 11076
rect 20312 11064 20318 11076
rect 22186 11064 22192 11076
rect 20312 11036 22192 11064
rect 20312 11024 20318 11036
rect 22186 11024 22192 11036
rect 22244 11024 22250 11076
rect 22925 11067 22983 11073
rect 22925 11033 22937 11067
rect 22971 11064 22983 11067
rect 24210 11064 24216 11076
rect 22971 11036 24216 11064
rect 22971 11033 22983 11036
rect 22925 11027 22983 11033
rect 24210 11024 24216 11036
rect 24268 11024 24274 11076
rect 24412 11064 24440 11095
rect 24670 11092 24676 11144
rect 24728 11092 24734 11144
rect 24762 11092 24768 11144
rect 24820 11092 24826 11144
rect 24946 11092 24952 11144
rect 25004 11092 25010 11144
rect 25314 11092 25320 11144
rect 25372 11132 25378 11144
rect 25501 11135 25559 11141
rect 25501 11132 25513 11135
rect 25372 11104 25513 11132
rect 25372 11092 25378 11104
rect 25501 11101 25513 11104
rect 25547 11101 25559 11135
rect 25501 11095 25559 11101
rect 25682 11092 25688 11144
rect 25740 11092 25746 11144
rect 25774 11092 25780 11144
rect 25832 11132 25838 11144
rect 26053 11135 26111 11141
rect 26053 11132 26065 11135
rect 25832 11104 26065 11132
rect 25832 11092 25838 11104
rect 26053 11101 26065 11104
rect 26099 11101 26111 11135
rect 26053 11095 26111 11101
rect 26234 11092 26240 11144
rect 26292 11092 26298 11144
rect 26326 11092 26332 11144
rect 26384 11092 26390 11144
rect 26513 11135 26571 11141
rect 26513 11101 26525 11135
rect 26559 11101 26571 11135
rect 26513 11095 26571 11101
rect 26605 11135 26663 11141
rect 26605 11101 26617 11135
rect 26651 11132 26663 11135
rect 26694 11132 26700 11144
rect 26651 11104 26700 11132
rect 26651 11101 26663 11104
rect 26605 11095 26663 11101
rect 24412 11036 24716 11064
rect 24688 11008 24716 11036
rect 24854 11024 24860 11076
rect 24912 11024 24918 11076
rect 26528 11064 26556 11095
rect 26694 11092 26700 11104
rect 26752 11092 26758 11144
rect 27062 11092 27068 11144
rect 27120 11092 27126 11144
rect 27246 11092 27252 11144
rect 27304 11092 27310 11144
rect 27338 11092 27344 11144
rect 27396 11092 27402 11144
rect 28166 11092 28172 11144
rect 28224 11092 28230 11144
rect 28258 11092 28264 11144
rect 28316 11132 28322 11144
rect 29360 11135 29418 11141
rect 29360 11132 29372 11135
rect 28316 11104 29372 11132
rect 28316 11092 28322 11104
rect 29360 11101 29372 11104
rect 29406 11101 29418 11135
rect 29360 11095 29418 11101
rect 29822 11092 29828 11144
rect 29880 11092 29886 11144
rect 29178 11064 29184 11076
rect 24964 11036 26556 11064
rect 26620 11036 29184 11064
rect 18230 10956 18236 11008
rect 18288 10996 18294 11008
rect 24578 10996 24584 11008
rect 18288 10968 24584 10996
rect 18288 10956 18294 10968
rect 24578 10956 24584 10968
rect 24636 10956 24642 11008
rect 24670 10956 24676 11008
rect 24728 10956 24734 11008
rect 24762 10956 24768 11008
rect 24820 10996 24826 11008
rect 24964 10996 24992 11036
rect 24820 10968 24992 10996
rect 25869 10999 25927 11005
rect 24820 10956 24826 10968
rect 25869 10965 25881 10999
rect 25915 10996 25927 10999
rect 26620 10996 26648 11036
rect 29178 11024 29184 11036
rect 29236 11024 29242 11076
rect 29457 11067 29515 11073
rect 29457 11033 29469 11067
rect 29503 11064 29515 11067
rect 32122 11064 32128 11076
rect 29503 11036 32128 11064
rect 29503 11033 29515 11036
rect 29457 11027 29515 11033
rect 32122 11024 32128 11036
rect 32180 11024 32186 11076
rect 25915 10968 26648 10996
rect 25915 10965 25927 10968
rect 25869 10959 25927 10965
rect 27154 10956 27160 11008
rect 27212 10996 27218 11008
rect 29638 10996 29644 11008
rect 27212 10968 29644 10996
rect 27212 10956 27218 10968
rect 29638 10956 29644 10968
rect 29696 10956 29702 11008
rect 2024 10906 77924 10928
rect 2024 10854 5794 10906
rect 5846 10854 5858 10906
rect 5910 10854 5922 10906
rect 5974 10854 5986 10906
rect 6038 10854 6050 10906
rect 6102 10854 36514 10906
rect 36566 10854 36578 10906
rect 36630 10854 36642 10906
rect 36694 10854 36706 10906
rect 36758 10854 36770 10906
rect 36822 10854 67234 10906
rect 67286 10854 67298 10906
rect 67350 10854 67362 10906
rect 67414 10854 67426 10906
rect 67478 10854 67490 10906
rect 67542 10854 77924 10906
rect 2024 10832 77924 10854
rect 20070 10752 20076 10804
rect 20128 10792 20134 10804
rect 20714 10792 20720 10804
rect 20128 10764 20720 10792
rect 20128 10752 20134 10764
rect 20714 10752 20720 10764
rect 20772 10792 20778 10804
rect 21913 10795 21971 10801
rect 20772 10764 21772 10792
rect 20772 10752 20778 10764
rect 17494 10684 17500 10736
rect 17552 10724 17558 10736
rect 21634 10724 21640 10736
rect 17552 10696 21640 10724
rect 17552 10684 17558 10696
rect 21634 10684 21640 10696
rect 21692 10684 21698 10736
rect 21744 10724 21772 10764
rect 21913 10761 21925 10795
rect 21959 10792 21971 10795
rect 22189 10795 22247 10801
rect 22189 10792 22201 10795
rect 21959 10764 22201 10792
rect 21959 10761 21971 10764
rect 21913 10755 21971 10761
rect 22189 10761 22201 10764
rect 22235 10792 22247 10795
rect 22235 10764 22692 10792
rect 22235 10761 22247 10764
rect 22189 10755 22247 10761
rect 22664 10724 22692 10764
rect 22738 10752 22744 10804
rect 22796 10792 22802 10804
rect 23014 10792 23020 10804
rect 22796 10764 23020 10792
rect 22796 10752 22802 10764
rect 23014 10752 23020 10764
rect 23072 10792 23078 10804
rect 27798 10792 27804 10804
rect 23072 10764 27804 10792
rect 23072 10752 23078 10764
rect 27798 10752 27804 10764
rect 27856 10752 27862 10804
rect 27890 10752 27896 10804
rect 27948 10752 27954 10804
rect 28166 10752 28172 10804
rect 28224 10792 28230 10804
rect 28905 10795 28963 10801
rect 28905 10792 28917 10795
rect 28224 10764 28917 10792
rect 28224 10752 28230 10764
rect 28905 10761 28917 10764
rect 28951 10761 28963 10795
rect 28905 10755 28963 10761
rect 29638 10752 29644 10804
rect 29696 10792 29702 10804
rect 30929 10795 30987 10801
rect 30929 10792 30941 10795
rect 29696 10764 30941 10792
rect 29696 10752 29702 10764
rect 30929 10761 30941 10764
rect 30975 10792 30987 10795
rect 30975 10764 31156 10792
rect 30975 10761 30987 10764
rect 30929 10755 30987 10761
rect 22830 10724 22836 10736
rect 21744 10696 22416 10724
rect 22664 10696 22836 10724
rect 19242 10616 19248 10668
rect 19300 10656 19306 10668
rect 20441 10659 20499 10665
rect 20441 10656 20453 10659
rect 19300 10628 20453 10656
rect 19300 10616 19306 10628
rect 20441 10625 20453 10628
rect 20487 10625 20499 10659
rect 20441 10619 20499 10625
rect 20714 10616 20720 10668
rect 20772 10616 20778 10668
rect 21266 10616 21272 10668
rect 21324 10616 21330 10668
rect 21744 10665 21772 10696
rect 21729 10659 21787 10665
rect 21729 10625 21741 10659
rect 21775 10625 21787 10659
rect 22005 10659 22063 10665
rect 22005 10654 22017 10659
rect 21729 10619 21787 10625
rect 21928 10626 22017 10654
rect 16666 10548 16672 10600
rect 16724 10588 16730 10600
rect 21928 10588 21956 10626
rect 22005 10625 22017 10626
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22097 10659 22155 10665
rect 22097 10625 22109 10659
rect 22143 10656 22155 10659
rect 22278 10656 22284 10668
rect 22143 10628 22284 10656
rect 22143 10625 22155 10628
rect 22097 10619 22155 10625
rect 22278 10616 22284 10628
rect 22336 10616 22342 10668
rect 22388 10665 22416 10696
rect 22830 10684 22836 10696
rect 22888 10724 22894 10736
rect 23290 10724 23296 10736
rect 22888 10696 23296 10724
rect 22888 10684 22894 10696
rect 23290 10684 23296 10696
rect 23348 10684 23354 10736
rect 23382 10684 23388 10736
rect 23440 10684 23446 10736
rect 27982 10684 27988 10736
rect 28040 10724 28046 10736
rect 28040 10696 31064 10724
rect 28040 10684 28046 10696
rect 22373 10659 22431 10665
rect 22373 10625 22385 10659
rect 22419 10656 22431 10659
rect 22738 10656 22744 10668
rect 22419 10628 22744 10656
rect 22419 10625 22431 10628
rect 22373 10619 22431 10625
rect 22738 10616 22744 10628
rect 22796 10616 22802 10668
rect 22925 10659 22983 10665
rect 22925 10625 22937 10659
rect 22971 10656 22983 10659
rect 23569 10659 23627 10665
rect 23569 10656 23581 10659
rect 22971 10628 23581 10656
rect 22971 10625 22983 10628
rect 22925 10619 22983 10625
rect 23569 10625 23581 10628
rect 23615 10625 23627 10659
rect 27341 10659 27399 10665
rect 27341 10656 27353 10659
rect 23569 10619 23627 10625
rect 24044 10628 27353 10656
rect 24044 10588 24072 10628
rect 27341 10625 27353 10628
rect 27387 10656 27399 10659
rect 27709 10659 27767 10665
rect 27709 10656 27721 10659
rect 27387 10628 27721 10656
rect 27387 10625 27399 10628
rect 27341 10619 27399 10625
rect 27709 10625 27721 10628
rect 27755 10625 27767 10659
rect 27709 10619 27767 10625
rect 27798 10616 27804 10668
rect 27856 10656 27862 10668
rect 27856 10628 28580 10656
rect 27856 10616 27862 10628
rect 16724 10560 21956 10588
rect 22066 10560 24072 10588
rect 16724 10548 16730 10560
rect 10502 10480 10508 10532
rect 10560 10520 10566 10532
rect 20717 10523 20775 10529
rect 20717 10520 20729 10523
rect 10560 10492 20729 10520
rect 10560 10480 10566 10492
rect 20717 10489 20729 10492
rect 20763 10489 20775 10523
rect 22066 10520 22094 10560
rect 24118 10548 24124 10600
rect 24176 10548 24182 10600
rect 24578 10548 24584 10600
rect 24636 10588 24642 10600
rect 25041 10591 25099 10597
rect 25041 10588 25053 10591
rect 24636 10560 25053 10588
rect 24636 10548 24642 10560
rect 25041 10557 25053 10560
rect 25087 10557 25099 10591
rect 25041 10551 25099 10557
rect 25130 10548 25136 10600
rect 25188 10588 25194 10600
rect 25317 10591 25375 10597
rect 25317 10588 25329 10591
rect 25188 10560 25329 10588
rect 25188 10548 25194 10560
rect 25317 10557 25329 10560
rect 25363 10557 25375 10591
rect 25317 10551 25375 10557
rect 25406 10548 25412 10600
rect 25464 10588 25470 10600
rect 26050 10588 26056 10600
rect 25464 10560 26056 10588
rect 25464 10548 25470 10560
rect 26050 10548 26056 10560
rect 26108 10548 26114 10600
rect 26234 10548 26240 10600
rect 26292 10548 26298 10600
rect 26602 10548 26608 10600
rect 26660 10588 26666 10600
rect 26789 10591 26847 10597
rect 26789 10588 26801 10591
rect 26660 10560 26801 10588
rect 26660 10548 26666 10560
rect 26789 10557 26801 10560
rect 26835 10557 26847 10591
rect 26789 10551 26847 10557
rect 26878 10548 26884 10600
rect 26936 10588 26942 10600
rect 28445 10591 28503 10597
rect 28445 10588 28457 10591
rect 26936 10560 28457 10588
rect 26936 10548 26942 10560
rect 28445 10557 28457 10560
rect 28491 10557 28503 10591
rect 28552 10588 28580 10628
rect 28810 10616 28816 10668
rect 28868 10616 28874 10668
rect 30282 10656 30288 10668
rect 28920 10628 30288 10656
rect 28920 10588 28948 10628
rect 30282 10616 30288 10628
rect 30340 10656 30346 10668
rect 31036 10665 31064 10696
rect 30745 10659 30803 10665
rect 30745 10656 30757 10659
rect 30340 10628 30757 10656
rect 30340 10616 30346 10628
rect 30745 10625 30757 10628
rect 30791 10625 30803 10659
rect 30745 10619 30803 10625
rect 31021 10659 31079 10665
rect 31021 10625 31033 10659
rect 31067 10625 31079 10659
rect 31128 10656 31156 10764
rect 31294 10752 31300 10804
rect 31352 10792 31358 10804
rect 31352 10764 35112 10792
rect 31352 10752 31358 10764
rect 31202 10684 31208 10736
rect 31260 10684 31266 10736
rect 34238 10724 34244 10736
rect 31726 10696 34244 10724
rect 31726 10656 31754 10696
rect 34238 10684 34244 10696
rect 34296 10684 34302 10736
rect 35084 10733 35112 10764
rect 35069 10727 35127 10733
rect 35069 10693 35081 10727
rect 35115 10693 35127 10727
rect 35069 10687 35127 10693
rect 31128 10628 31754 10656
rect 33505 10659 33563 10665
rect 31021 10619 31079 10625
rect 33505 10625 33517 10659
rect 33551 10656 33563 10659
rect 33870 10656 33876 10668
rect 33551 10628 33876 10656
rect 33551 10625 33563 10628
rect 33505 10619 33563 10625
rect 33870 10616 33876 10628
rect 33928 10616 33934 10668
rect 34882 10616 34888 10668
rect 34940 10616 34946 10668
rect 35158 10616 35164 10668
rect 35216 10616 35222 10668
rect 35253 10659 35311 10665
rect 35253 10625 35265 10659
rect 35299 10625 35311 10659
rect 35253 10619 35311 10625
rect 28552 10560 28948 10588
rect 28445 10551 28503 10557
rect 28994 10548 29000 10600
rect 29052 10588 29058 10600
rect 29457 10591 29515 10597
rect 29457 10588 29469 10591
rect 29052 10560 29469 10588
rect 29052 10548 29058 10560
rect 29457 10557 29469 10560
rect 29503 10557 29515 10591
rect 29457 10551 29515 10557
rect 29641 10591 29699 10597
rect 29641 10557 29653 10591
rect 29687 10588 29699 10591
rect 29730 10588 29736 10600
rect 29687 10560 29736 10588
rect 29687 10557 29699 10560
rect 29641 10551 29699 10557
rect 29730 10548 29736 10560
rect 29788 10548 29794 10600
rect 31478 10548 31484 10600
rect 31536 10588 31542 10600
rect 31536 10560 31754 10588
rect 31536 10548 31542 10560
rect 31726 10532 31754 10560
rect 33134 10548 33140 10600
rect 33192 10588 33198 10600
rect 33229 10591 33287 10597
rect 33229 10588 33241 10591
rect 33192 10560 33241 10588
rect 33192 10548 33198 10560
rect 33229 10557 33241 10560
rect 33275 10557 33287 10591
rect 33229 10551 33287 10557
rect 33318 10548 33324 10600
rect 33376 10548 33382 10600
rect 33413 10591 33471 10597
rect 33413 10557 33425 10591
rect 33459 10557 33471 10591
rect 33413 10551 33471 10557
rect 30561 10523 30619 10529
rect 30561 10520 30573 10523
rect 20717 10483 20775 10489
rect 20824 10492 22094 10520
rect 29104 10492 30573 10520
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 20824 10452 20852 10492
rect 14792 10424 20852 10452
rect 14792 10412 14798 10424
rect 21358 10412 21364 10464
rect 21416 10412 21422 10464
rect 21542 10412 21548 10464
rect 21600 10412 21606 10464
rect 22557 10455 22615 10461
rect 22557 10421 22569 10455
rect 22603 10452 22615 10455
rect 22646 10452 22652 10464
rect 22603 10424 22652 10452
rect 22603 10421 22615 10424
rect 22557 10415 22615 10421
rect 22646 10412 22652 10424
rect 22704 10412 22710 10464
rect 22738 10412 22744 10464
rect 22796 10412 22802 10464
rect 23106 10412 23112 10464
rect 23164 10412 23170 10464
rect 23198 10412 23204 10464
rect 23256 10452 23262 10464
rect 23842 10452 23848 10464
rect 23256 10424 23848 10452
rect 23256 10412 23262 10424
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 24489 10455 24547 10461
rect 24489 10421 24501 10455
rect 24535 10452 24547 10455
rect 24578 10452 24584 10464
rect 24535 10424 24584 10452
rect 24535 10421 24547 10424
rect 24489 10415 24547 10421
rect 24578 10412 24584 10424
rect 24636 10412 24642 10464
rect 24670 10412 24676 10464
rect 24728 10452 24734 10464
rect 25406 10452 25412 10464
rect 24728 10424 25412 10452
rect 24728 10412 24734 10424
rect 25406 10412 25412 10424
rect 25464 10412 25470 10464
rect 25958 10412 25964 10464
rect 26016 10412 26022 10464
rect 26050 10412 26056 10464
rect 26108 10452 26114 10464
rect 26602 10452 26608 10464
rect 26108 10424 26608 10452
rect 26108 10412 26114 10424
rect 26602 10412 26608 10424
rect 26660 10412 26666 10464
rect 27522 10412 27528 10464
rect 27580 10412 27586 10464
rect 28626 10412 28632 10464
rect 28684 10412 28690 10464
rect 28810 10412 28816 10464
rect 28868 10452 28874 10464
rect 29104 10452 29132 10492
rect 30561 10489 30573 10492
rect 30607 10489 30619 10523
rect 30561 10483 30619 10489
rect 31662 10480 31668 10532
rect 31720 10520 31754 10532
rect 33428 10520 33456 10551
rect 33594 10548 33600 10600
rect 33652 10588 33658 10600
rect 33689 10591 33747 10597
rect 33689 10588 33701 10591
rect 33652 10560 33701 10588
rect 33652 10548 33658 10560
rect 33689 10557 33701 10560
rect 33735 10557 33747 10591
rect 33888 10588 33916 10616
rect 35268 10588 35296 10619
rect 33888 10560 35296 10588
rect 33689 10551 33747 10557
rect 31720 10492 33456 10520
rect 31720 10480 31726 10492
rect 28868 10424 29132 10452
rect 28868 10412 28874 10424
rect 30190 10412 30196 10464
rect 30248 10412 30254 10464
rect 31481 10455 31539 10461
rect 31481 10421 31493 10455
rect 31527 10452 31539 10455
rect 32306 10452 32312 10464
rect 31527 10424 32312 10452
rect 31527 10421 31539 10424
rect 31481 10415 31539 10421
rect 32306 10412 32312 10424
rect 32364 10412 32370 10464
rect 32490 10412 32496 10464
rect 32548 10452 32554 10464
rect 33045 10455 33103 10461
rect 33045 10452 33057 10455
rect 32548 10424 33057 10452
rect 32548 10412 32554 10424
rect 33045 10421 33057 10424
rect 33091 10421 33103 10455
rect 33045 10415 33103 10421
rect 34241 10455 34299 10461
rect 34241 10421 34253 10455
rect 34287 10452 34299 10455
rect 34790 10452 34796 10464
rect 34287 10424 34796 10452
rect 34287 10421 34299 10424
rect 34241 10415 34299 10421
rect 34790 10412 34796 10424
rect 34848 10412 34854 10464
rect 35434 10412 35440 10464
rect 35492 10412 35498 10464
rect 2024 10362 77924 10384
rect 2024 10310 5134 10362
rect 5186 10310 5198 10362
rect 5250 10310 5262 10362
rect 5314 10310 5326 10362
rect 5378 10310 5390 10362
rect 5442 10310 35854 10362
rect 35906 10310 35918 10362
rect 35970 10310 35982 10362
rect 36034 10310 36046 10362
rect 36098 10310 36110 10362
rect 36162 10310 66574 10362
rect 66626 10310 66638 10362
rect 66690 10310 66702 10362
rect 66754 10310 66766 10362
rect 66818 10310 66830 10362
rect 66882 10310 77924 10362
rect 2024 10288 77924 10310
rect 19797 10251 19855 10257
rect 19797 10217 19809 10251
rect 19843 10248 19855 10251
rect 19886 10248 19892 10260
rect 19843 10220 19892 10248
rect 19843 10217 19855 10220
rect 19797 10211 19855 10217
rect 19886 10208 19892 10220
rect 19944 10208 19950 10260
rect 19978 10208 19984 10260
rect 20036 10208 20042 10260
rect 21450 10248 21456 10260
rect 21008 10220 21456 10248
rect 16850 10140 16856 10192
rect 16908 10180 16914 10192
rect 21008 10180 21036 10220
rect 21450 10208 21456 10220
rect 21508 10208 21514 10260
rect 23198 10248 23204 10260
rect 22112 10220 23204 10248
rect 22112 10180 22140 10220
rect 23198 10208 23204 10220
rect 23256 10208 23262 10260
rect 23290 10208 23296 10260
rect 23348 10248 23354 10260
rect 24670 10248 24676 10260
rect 23348 10220 24676 10248
rect 23348 10208 23354 10220
rect 24670 10208 24676 10220
rect 24728 10248 24734 10260
rect 27154 10248 27160 10260
rect 24728 10220 27160 10248
rect 24728 10208 24734 10220
rect 27154 10208 27160 10220
rect 27212 10208 27218 10260
rect 27430 10208 27436 10260
rect 27488 10248 27494 10260
rect 27525 10251 27583 10257
rect 27525 10248 27537 10251
rect 27488 10220 27537 10248
rect 27488 10208 27494 10220
rect 27525 10217 27537 10220
rect 27571 10217 27583 10251
rect 27525 10211 27583 10217
rect 28534 10208 28540 10260
rect 28592 10208 28598 10260
rect 30282 10208 30288 10260
rect 30340 10248 30346 10260
rect 34330 10248 34336 10260
rect 30340 10220 34336 10248
rect 30340 10208 30346 10220
rect 34330 10208 34336 10220
rect 34388 10208 34394 10260
rect 27617 10183 27675 10189
rect 27617 10180 27629 10183
rect 16908 10152 21036 10180
rect 21284 10152 22140 10180
rect 23308 10152 27629 10180
rect 16908 10140 16914 10152
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 20993 10115 21051 10121
rect 20993 10112 21005 10115
rect 20864 10084 21005 10112
rect 20864 10072 20870 10084
rect 20993 10081 21005 10084
rect 21039 10081 21051 10115
rect 20993 10075 21051 10081
rect 19426 10004 19432 10056
rect 19484 10044 19490 10056
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 19484 10016 19625 10044
rect 19484 10004 19490 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 19613 10007 19671 10013
rect 19702 10004 19708 10056
rect 19760 10004 19766 10056
rect 20717 10047 20775 10053
rect 20717 10013 20729 10047
rect 20763 10013 20775 10047
rect 20717 10007 20775 10013
rect 13722 9936 13728 9988
rect 13780 9976 13786 9988
rect 20732 9976 20760 10007
rect 20898 10004 20904 10056
rect 20956 10004 20962 10056
rect 21082 9976 21088 9988
rect 13780 9948 20668 9976
rect 20732 9948 21088 9976
rect 13780 9936 13786 9948
rect 20530 9868 20536 9920
rect 20588 9868 20594 9920
rect 20640 9908 20668 9948
rect 21082 9936 21088 9948
rect 21140 9936 21146 9988
rect 21284 9908 21312 10152
rect 21450 10072 21456 10124
rect 21508 10112 21514 10124
rect 21508 10084 22048 10112
rect 21508 10072 21514 10084
rect 21818 10004 21824 10056
rect 21876 10044 21882 10056
rect 21913 10047 21971 10053
rect 21913 10044 21925 10047
rect 21876 10016 21925 10044
rect 21876 10004 21882 10016
rect 21913 10013 21925 10016
rect 21959 10013 21971 10047
rect 22020 10044 22048 10084
rect 22646 10072 22652 10124
rect 22704 10072 22710 10124
rect 22738 10044 22744 10056
rect 22020 10016 22744 10044
rect 21913 10007 21971 10013
rect 22738 10004 22744 10016
rect 22796 10004 22802 10056
rect 22922 10004 22928 10056
rect 22980 10044 22986 10056
rect 23308 10044 23336 10152
rect 27617 10149 27629 10152
rect 27663 10149 27675 10183
rect 37182 10180 37188 10192
rect 27617 10143 27675 10149
rect 31128 10152 37188 10180
rect 23842 10072 23848 10124
rect 23900 10112 23906 10124
rect 31128 10121 31156 10152
rect 37182 10140 37188 10152
rect 37240 10140 37246 10192
rect 25961 10115 26019 10121
rect 25961 10112 25973 10115
rect 23900 10084 25973 10112
rect 23900 10072 23906 10084
rect 25961 10081 25973 10084
rect 26007 10112 26019 10115
rect 26697 10115 26755 10121
rect 26697 10112 26709 10115
rect 26007 10084 26709 10112
rect 26007 10081 26019 10084
rect 25961 10075 26019 10081
rect 26697 10081 26709 10084
rect 26743 10081 26755 10115
rect 27893 10115 27951 10121
rect 27893 10112 27905 10115
rect 26697 10075 26755 10081
rect 27356 10084 27905 10112
rect 27356 10056 27384 10084
rect 27893 10081 27905 10084
rect 27939 10081 27951 10115
rect 27893 10075 27951 10081
rect 31113 10115 31171 10121
rect 31113 10081 31125 10115
rect 31159 10081 31171 10115
rect 31113 10075 31171 10081
rect 31202 10072 31208 10124
rect 31260 10072 31266 10124
rect 31941 10115 31999 10121
rect 31941 10112 31953 10115
rect 31726 10084 31953 10112
rect 22980 10016 23336 10044
rect 22980 10004 22986 10016
rect 23474 10004 23480 10056
rect 23532 10004 23538 10056
rect 24118 10004 24124 10056
rect 24176 10004 24182 10056
rect 24581 10047 24639 10053
rect 24581 10013 24593 10047
rect 24627 10044 24639 10047
rect 25130 10044 25136 10056
rect 24627 10016 25136 10044
rect 24627 10013 24639 10016
rect 24581 10007 24639 10013
rect 25130 10004 25136 10016
rect 25188 10004 25194 10056
rect 25498 10004 25504 10056
rect 25556 10004 25562 10056
rect 25590 10004 25596 10056
rect 25648 10044 25654 10056
rect 25685 10047 25743 10053
rect 25685 10044 25697 10047
rect 25648 10016 25697 10044
rect 25648 10004 25654 10016
rect 25685 10013 25697 10016
rect 25731 10013 25743 10047
rect 26050 10044 26056 10056
rect 25685 10007 25743 10013
rect 25792 10016 26056 10044
rect 22002 9936 22008 9988
rect 22060 9976 22066 9988
rect 22833 9979 22891 9985
rect 22833 9976 22845 9979
rect 22060 9948 22845 9976
rect 22060 9936 22066 9948
rect 22833 9945 22845 9948
rect 22879 9945 22891 9979
rect 22833 9939 22891 9945
rect 23290 9936 23296 9988
rect 23348 9976 23354 9988
rect 25792 9976 25820 10016
rect 26050 10004 26056 10016
rect 26108 10004 26114 10056
rect 26602 10004 26608 10056
rect 26660 10044 26666 10056
rect 26881 10047 26939 10053
rect 26881 10044 26893 10047
rect 26660 10016 26893 10044
rect 26660 10004 26666 10016
rect 26881 10013 26893 10016
rect 26927 10013 26939 10047
rect 26881 10007 26939 10013
rect 27338 10004 27344 10056
rect 27396 10004 27402 10056
rect 27798 10004 27804 10056
rect 27856 10004 27862 10056
rect 29454 10004 29460 10056
rect 29512 10044 29518 10056
rect 29641 10047 29699 10053
rect 29641 10044 29653 10047
rect 29512 10016 29653 10044
rect 29512 10004 29518 10016
rect 29641 10013 29653 10016
rect 29687 10013 29699 10047
rect 29641 10007 29699 10013
rect 23348 9948 25820 9976
rect 23348 9936 23354 9948
rect 25866 9936 25872 9988
rect 25924 9936 25930 9988
rect 29546 9936 29552 9988
rect 29604 9976 29610 9988
rect 31726 9976 31754 10084
rect 31941 10081 31953 10084
rect 31987 10081 31999 10115
rect 31941 10075 31999 10081
rect 32950 10072 32956 10124
rect 33008 10112 33014 10124
rect 33505 10115 33563 10121
rect 33505 10112 33517 10115
rect 33008 10084 33517 10112
rect 33008 10072 33014 10084
rect 33505 10081 33517 10084
rect 33551 10081 33563 10115
rect 33505 10075 33563 10081
rect 34790 10072 34796 10124
rect 34848 10072 34854 10124
rect 31846 10004 31852 10056
rect 31904 10004 31910 10056
rect 32582 10004 32588 10056
rect 32640 10044 32646 10056
rect 32677 10047 32735 10053
rect 32677 10044 32689 10047
rect 32640 10016 32689 10044
rect 32640 10004 32646 10016
rect 32677 10013 32689 10016
rect 32723 10013 32735 10047
rect 32677 10007 32735 10013
rect 32858 10004 32864 10056
rect 32916 10044 32922 10056
rect 34057 10047 34115 10053
rect 34057 10044 34069 10047
rect 32916 10016 34069 10044
rect 32916 10004 32922 10016
rect 34057 10013 34069 10016
rect 34103 10013 34115 10047
rect 34057 10007 34115 10013
rect 35618 10004 35624 10056
rect 35676 10004 35682 10056
rect 36725 10047 36783 10053
rect 36725 10013 36737 10047
rect 36771 10044 36783 10047
rect 36906 10044 36912 10056
rect 36771 10016 36912 10044
rect 36771 10013 36783 10016
rect 36725 10007 36783 10013
rect 36906 10004 36912 10016
rect 36964 10004 36970 10056
rect 29604 9948 31754 9976
rect 29604 9936 29610 9948
rect 32398 9936 32404 9988
rect 32456 9976 32462 9988
rect 34241 9979 34299 9985
rect 34241 9976 34253 9979
rect 32456 9948 34253 9976
rect 32456 9936 32462 9948
rect 34241 9945 34253 9948
rect 34287 9945 34299 9979
rect 34241 9939 34299 9945
rect 20640 9880 21312 9908
rect 21358 9868 21364 9920
rect 21416 9868 21422 9920
rect 22094 9868 22100 9920
rect 22152 9868 22158 9920
rect 22370 9868 22376 9920
rect 22428 9908 22434 9920
rect 23106 9908 23112 9920
rect 22428 9880 23112 9908
rect 22428 9868 22434 9880
rect 23106 9868 23112 9880
rect 23164 9868 23170 9920
rect 23474 9868 23480 9920
rect 23532 9908 23538 9920
rect 23569 9911 23627 9917
rect 23569 9908 23581 9911
rect 23532 9880 23581 9908
rect 23532 9868 23538 9880
rect 23569 9877 23581 9880
rect 23615 9877 23627 9911
rect 23569 9871 23627 9877
rect 25038 9868 25044 9920
rect 25096 9908 25102 9920
rect 25133 9911 25191 9917
rect 25133 9908 25145 9911
rect 25096 9880 25145 9908
rect 25096 9868 25102 9880
rect 25133 9877 25145 9880
rect 25179 9877 25191 9911
rect 25133 9871 25191 9877
rect 25222 9868 25228 9920
rect 25280 9908 25286 9920
rect 25317 9911 25375 9917
rect 25317 9908 25329 9911
rect 25280 9880 25329 9908
rect 25280 9868 25286 9880
rect 25317 9877 25329 9880
rect 25363 9877 25375 9911
rect 25317 9871 25375 9877
rect 25406 9868 25412 9920
rect 25464 9908 25470 9920
rect 25593 9911 25651 9917
rect 25593 9908 25605 9911
rect 25464 9880 25605 9908
rect 25464 9868 25470 9880
rect 25593 9877 25605 9880
rect 25639 9908 25651 9911
rect 26050 9908 26056 9920
rect 25639 9880 26056 9908
rect 25639 9877 25651 9880
rect 25593 9871 25651 9877
rect 26050 9868 26056 9880
rect 26108 9868 26114 9920
rect 26142 9868 26148 9920
rect 26200 9868 26206 9920
rect 28626 9868 28632 9920
rect 28684 9868 28690 9920
rect 28994 9868 29000 9920
rect 29052 9868 29058 9920
rect 30006 9868 30012 9920
rect 30064 9908 30070 9920
rect 30285 9911 30343 9917
rect 30285 9908 30297 9911
rect 30064 9880 30297 9908
rect 30064 9868 30070 9880
rect 30285 9877 30297 9880
rect 30331 9877 30343 9911
rect 30285 9871 30343 9877
rect 30466 9868 30472 9920
rect 30524 9868 30530 9920
rect 32585 9911 32643 9917
rect 32585 9877 32597 9911
rect 32631 9908 32643 9911
rect 32674 9908 32680 9920
rect 32631 9880 32680 9908
rect 32631 9877 32643 9880
rect 32585 9871 32643 9877
rect 32674 9868 32680 9880
rect 32732 9868 32738 9920
rect 33321 9911 33379 9917
rect 33321 9877 33333 9911
rect 33367 9908 33379 9911
rect 33410 9908 33416 9920
rect 33367 9880 33416 9908
rect 33367 9877 33379 9880
rect 33321 9871 33379 9877
rect 33410 9868 33416 9880
rect 33468 9868 33474 9920
rect 36262 9868 36268 9920
rect 36320 9868 36326 9920
rect 37277 9911 37335 9917
rect 37277 9877 37289 9911
rect 37323 9908 37335 9911
rect 38746 9908 38752 9920
rect 37323 9880 38752 9908
rect 37323 9877 37335 9880
rect 37277 9871 37335 9877
rect 38746 9868 38752 9880
rect 38804 9868 38810 9920
rect 2024 9818 77924 9840
rect 2024 9766 5794 9818
rect 5846 9766 5858 9818
rect 5910 9766 5922 9818
rect 5974 9766 5986 9818
rect 6038 9766 6050 9818
rect 6102 9766 36514 9818
rect 36566 9766 36578 9818
rect 36630 9766 36642 9818
rect 36694 9766 36706 9818
rect 36758 9766 36770 9818
rect 36822 9766 67234 9818
rect 67286 9766 67298 9818
rect 67350 9766 67362 9818
rect 67414 9766 67426 9818
rect 67478 9766 67490 9818
rect 67542 9766 77924 9818
rect 2024 9744 77924 9766
rect 23566 9704 23572 9716
rect 18800 9676 19656 9704
rect 15562 9596 15568 9648
rect 15620 9636 15626 9648
rect 18800 9636 18828 9676
rect 19628 9674 19656 9676
rect 22480 9676 23572 9704
rect 15620 9608 18828 9636
rect 15620 9596 15626 9608
rect 18874 9596 18880 9648
rect 18932 9636 18938 9648
rect 19334 9636 19340 9648
rect 18932 9608 19340 9636
rect 18932 9596 18938 9608
rect 19334 9596 19340 9608
rect 19392 9596 19398 9648
rect 19628 9646 19748 9674
rect 18690 9528 18696 9580
rect 18748 9528 18754 9580
rect 19150 9528 19156 9580
rect 19208 9528 19214 9580
rect 19426 9577 19432 9614
rect 19245 9571 19303 9577
rect 19245 9537 19257 9571
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 19423 9562 19432 9577
rect 19484 9562 19490 9614
rect 19521 9571 19579 9577
rect 19423 9537 19435 9562
rect 19469 9537 19481 9562
rect 19423 9531 19481 9537
rect 19521 9537 19533 9571
rect 19567 9568 19579 9571
rect 19610 9568 19616 9614
rect 19567 9562 19616 9568
rect 19668 9562 19674 9614
rect 19720 9577 19748 9646
rect 21729 9639 21787 9645
rect 21729 9605 21741 9639
rect 21775 9636 21787 9639
rect 22480 9636 22508 9676
rect 23566 9664 23572 9676
rect 23624 9664 23630 9716
rect 24118 9664 24124 9716
rect 24176 9664 24182 9716
rect 24320 9676 24808 9704
rect 21775 9608 22508 9636
rect 21775 9605 21787 9608
rect 21729 9599 21787 9605
rect 22554 9596 22560 9648
rect 22612 9596 22618 9648
rect 24320 9636 24348 9676
rect 22756 9608 24348 9636
rect 24381 9639 24439 9645
rect 19705 9571 19763 9577
rect 19567 9540 19656 9562
rect 19567 9537 19579 9540
rect 19521 9531 19579 9537
rect 19705 9537 19717 9571
rect 19751 9568 19763 9571
rect 19751 9540 19932 9568
rect 19751 9537 19763 9540
rect 19705 9531 19763 9537
rect 19058 9460 19064 9512
rect 19116 9500 19122 9512
rect 19260 9500 19288 9531
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19116 9472 19625 9500
rect 19116 9460 19122 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 19797 9503 19855 9509
rect 19797 9469 19809 9503
rect 19843 9469 19855 9503
rect 19797 9463 19855 9469
rect 18877 9435 18935 9441
rect 18877 9401 18889 9435
rect 18923 9432 18935 9435
rect 19812 9432 19840 9463
rect 18923 9404 19840 9432
rect 19904 9432 19932 9540
rect 19978 9528 19984 9580
rect 20036 9568 20042 9580
rect 20036 9540 21956 9568
rect 20036 9528 20042 9540
rect 20441 9503 20499 9509
rect 20441 9469 20453 9503
rect 20487 9500 20499 9503
rect 20533 9503 20591 9509
rect 20533 9500 20545 9503
rect 20487 9472 20545 9500
rect 20487 9469 20499 9472
rect 20441 9463 20499 9469
rect 20533 9469 20545 9472
rect 20579 9469 20591 9503
rect 20533 9463 20591 9469
rect 21361 9503 21419 9509
rect 21361 9469 21373 9503
rect 21407 9500 21419 9503
rect 21818 9500 21824 9512
rect 21407 9472 21824 9500
rect 21407 9469 21419 9472
rect 21361 9463 21419 9469
rect 21818 9460 21824 9472
rect 21876 9460 21882 9512
rect 21928 9500 21956 9540
rect 22002 9528 22008 9580
rect 22060 9528 22066 9580
rect 22756 9577 22784 9608
rect 24381 9605 24393 9639
rect 24427 9636 24439 9639
rect 24486 9636 24492 9648
rect 24427 9608 24492 9636
rect 24427 9605 24439 9608
rect 24381 9599 24439 9605
rect 24486 9596 24492 9608
rect 24544 9596 24550 9648
rect 24581 9639 24639 9645
rect 24581 9605 24593 9639
rect 24627 9636 24639 9639
rect 24670 9636 24676 9648
rect 24627 9608 24676 9636
rect 24627 9605 24639 9608
rect 24581 9599 24639 9605
rect 24670 9596 24676 9608
rect 24728 9596 24734 9648
rect 24780 9636 24808 9676
rect 27798 9664 27804 9716
rect 27856 9704 27862 9716
rect 28813 9707 28871 9713
rect 28813 9704 28825 9707
rect 27856 9676 28825 9704
rect 27856 9664 27862 9676
rect 28813 9673 28825 9676
rect 28859 9673 28871 9707
rect 28813 9667 28871 9673
rect 33229 9707 33287 9713
rect 33229 9673 33241 9707
rect 33275 9704 33287 9707
rect 33318 9704 33324 9716
rect 33275 9676 33324 9704
rect 33275 9673 33287 9676
rect 33229 9667 33287 9673
rect 33318 9664 33324 9676
rect 33376 9664 33382 9716
rect 26510 9636 26516 9648
rect 24780 9608 26516 9636
rect 26510 9596 26516 9608
rect 26568 9596 26574 9648
rect 26605 9639 26663 9645
rect 26605 9605 26617 9639
rect 26651 9636 26663 9639
rect 26878 9636 26884 9648
rect 26651 9608 26884 9636
rect 26651 9605 26663 9608
rect 26605 9599 26663 9605
rect 26878 9596 26884 9608
rect 26936 9596 26942 9648
rect 27706 9596 27712 9648
rect 27764 9636 27770 9648
rect 27893 9639 27951 9645
rect 27893 9636 27905 9639
rect 27764 9608 27905 9636
rect 27764 9596 27770 9608
rect 27893 9605 27905 9608
rect 27939 9636 27951 9639
rect 27939 9608 28120 9636
rect 27939 9605 27951 9608
rect 27893 9599 27951 9605
rect 22741 9571 22799 9577
rect 22741 9537 22753 9571
rect 22787 9537 22799 9571
rect 22741 9531 22799 9537
rect 22830 9528 22836 9580
rect 22888 9528 22894 9580
rect 23014 9528 23020 9580
rect 23072 9528 23078 9580
rect 25409 9571 25467 9577
rect 25409 9568 25421 9571
rect 23216 9540 25421 9568
rect 23216 9500 23244 9540
rect 25409 9537 25421 9540
rect 25455 9537 25467 9571
rect 25409 9531 25467 9537
rect 25958 9528 25964 9580
rect 26016 9528 26022 9580
rect 28092 9577 28120 9608
rect 28534 9596 28540 9648
rect 28592 9636 28598 9648
rect 28592 9608 29776 9636
rect 28592 9596 28598 9608
rect 29748 9577 29776 9608
rect 30650 9596 30656 9648
rect 30708 9636 30714 9648
rect 31570 9636 31576 9648
rect 30708 9608 31576 9636
rect 30708 9596 30714 9608
rect 31570 9596 31576 9608
rect 31628 9596 31634 9648
rect 32858 9596 32864 9648
rect 32916 9596 32922 9648
rect 34425 9639 34483 9645
rect 34425 9636 34437 9639
rect 32968 9608 34437 9636
rect 28077 9571 28135 9577
rect 28077 9537 28089 9571
rect 28123 9537 28135 9571
rect 29549 9571 29607 9577
rect 29549 9568 29561 9571
rect 28077 9531 28135 9537
rect 28552 9540 29561 9568
rect 21928 9472 23244 9500
rect 23290 9460 23296 9512
rect 23348 9500 23354 9512
rect 23477 9503 23535 9509
rect 23477 9500 23489 9503
rect 23348 9472 23489 9500
rect 23348 9460 23354 9472
rect 23477 9469 23489 9472
rect 23523 9469 23535 9503
rect 25222 9500 25228 9512
rect 23477 9463 23535 9469
rect 24136 9472 25228 9500
rect 21177 9435 21235 9441
rect 19904 9404 21128 9432
rect 18923 9401 18935 9404
rect 18877 9395 18935 9401
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 18969 9367 19027 9373
rect 18969 9364 18981 9367
rect 13872 9336 18981 9364
rect 13872 9324 13878 9336
rect 18969 9333 18981 9336
rect 19015 9333 19027 9367
rect 18969 9327 19027 9333
rect 19429 9367 19487 9373
rect 19429 9333 19441 9367
rect 19475 9364 19487 9367
rect 20990 9364 20996 9376
rect 19475 9336 20996 9364
rect 19475 9333 19487 9336
rect 19429 9327 19487 9333
rect 20990 9324 20996 9336
rect 21048 9324 21054 9376
rect 21100 9364 21128 9404
rect 21177 9401 21189 9435
rect 21223 9432 21235 9435
rect 21726 9432 21732 9444
rect 21223 9404 21732 9432
rect 21223 9401 21235 9404
rect 21177 9395 21235 9401
rect 21726 9392 21732 9404
rect 21784 9392 21790 9444
rect 23106 9392 23112 9444
rect 23164 9432 23170 9444
rect 24136 9432 24164 9472
rect 25222 9460 25228 9472
rect 25280 9460 25286 9512
rect 25317 9503 25375 9509
rect 25317 9469 25329 9503
rect 25363 9500 25375 9503
rect 25498 9500 25504 9512
rect 25363 9472 25504 9500
rect 25363 9469 25375 9472
rect 25317 9463 25375 9469
rect 25498 9460 25504 9472
rect 25556 9460 25562 9512
rect 27154 9460 27160 9512
rect 27212 9460 27218 9512
rect 28552 9500 28580 9540
rect 29549 9537 29561 9540
rect 29595 9537 29607 9571
rect 29549 9531 29607 9537
rect 29733 9571 29791 9577
rect 29733 9537 29745 9571
rect 29779 9537 29791 9571
rect 32968 9568 32996 9608
rect 34425 9605 34437 9608
rect 34471 9605 34483 9639
rect 34425 9599 34483 9605
rect 29733 9531 29791 9537
rect 31588 9540 32996 9568
rect 31588 9512 31616 9540
rect 33042 9528 33048 9580
rect 33100 9528 33106 9580
rect 33226 9528 33232 9580
rect 33284 9568 33290 9580
rect 33321 9571 33379 9577
rect 33321 9568 33333 9571
rect 33284 9540 33333 9568
rect 33284 9528 33290 9540
rect 33321 9537 33333 9540
rect 33367 9537 33379 9571
rect 33321 9531 33379 9537
rect 33413 9571 33471 9577
rect 33413 9537 33425 9571
rect 33459 9568 33471 9571
rect 33502 9568 33508 9580
rect 33459 9540 33508 9568
rect 33459 9537 33471 9540
rect 33413 9531 33471 9537
rect 33502 9528 33508 9540
rect 33560 9528 33566 9580
rect 35897 9571 35955 9577
rect 35897 9537 35909 9571
rect 35943 9568 35955 9571
rect 36262 9568 36268 9580
rect 35943 9540 36268 9568
rect 35943 9537 35955 9540
rect 35897 9531 35955 9537
rect 36262 9528 36268 9540
rect 36320 9528 36326 9580
rect 38746 9528 38752 9580
rect 38804 9528 38810 9580
rect 28000 9472 28580 9500
rect 23164 9404 24164 9432
rect 23164 9392 23170 9404
rect 24210 9392 24216 9444
rect 24268 9392 24274 9444
rect 24670 9392 24676 9444
rect 24728 9392 24734 9444
rect 25240 9432 25268 9460
rect 28000 9432 28028 9472
rect 28442 9432 28448 9444
rect 25240 9404 28028 9432
rect 28092 9404 28448 9432
rect 21637 9367 21695 9373
rect 21637 9364 21649 9367
rect 21100 9336 21649 9364
rect 21637 9333 21649 9336
rect 21683 9333 21695 9367
rect 21637 9327 21695 9333
rect 23198 9324 23204 9376
rect 23256 9324 23262 9376
rect 23290 9324 23296 9376
rect 23348 9324 23354 9376
rect 23566 9324 23572 9376
rect 23624 9364 23630 9376
rect 23842 9364 23848 9376
rect 23624 9336 23848 9364
rect 23624 9324 23630 9336
rect 23842 9324 23848 9336
rect 23900 9364 23906 9376
rect 24397 9367 24455 9373
rect 24397 9364 24409 9367
rect 23900 9336 24409 9364
rect 23900 9324 23906 9336
rect 24397 9333 24409 9336
rect 24443 9333 24455 9367
rect 24397 9327 24455 9333
rect 25314 9324 25320 9376
rect 25372 9364 25378 9376
rect 28092 9364 28120 9404
rect 28442 9392 28448 9404
rect 28500 9392 28506 9444
rect 28552 9432 28580 9472
rect 28626 9460 28632 9512
rect 28684 9500 28690 9512
rect 29365 9503 29423 9509
rect 29365 9500 29377 9503
rect 28684 9472 29377 9500
rect 28684 9460 28690 9472
rect 29365 9469 29377 9472
rect 29411 9469 29423 9503
rect 29365 9463 29423 9469
rect 29638 9460 29644 9512
rect 29696 9500 29702 9512
rect 30009 9503 30067 9509
rect 30009 9500 30021 9503
rect 29696 9472 30021 9500
rect 29696 9460 29702 9472
rect 30009 9469 30021 9472
rect 30055 9469 30067 9503
rect 30009 9463 30067 9469
rect 30653 9503 30711 9509
rect 30653 9469 30665 9503
rect 30699 9500 30711 9503
rect 30926 9500 30932 9512
rect 30699 9472 30932 9500
rect 30699 9469 30711 9472
rect 30653 9463 30711 9469
rect 30926 9460 30932 9472
rect 30984 9460 30990 9512
rect 31294 9460 31300 9512
rect 31352 9460 31358 9512
rect 31570 9460 31576 9512
rect 31628 9460 31634 9512
rect 32030 9460 32036 9512
rect 32088 9460 32094 9512
rect 32214 9460 32220 9512
rect 32272 9460 32278 9512
rect 33689 9503 33747 9509
rect 33689 9500 33701 9503
rect 32416 9472 33701 9500
rect 28994 9432 29000 9444
rect 28552 9404 29000 9432
rect 28994 9392 29000 9404
rect 29052 9392 29058 9444
rect 29086 9392 29092 9444
rect 29144 9432 29150 9444
rect 31481 9435 31539 9441
rect 31481 9432 31493 9435
rect 29144 9404 31493 9432
rect 29144 9392 29150 9404
rect 31481 9401 31493 9404
rect 31527 9401 31539 9435
rect 31481 9395 31539 9401
rect 25372 9336 28120 9364
rect 25372 9324 25378 9336
rect 28350 9324 28356 9376
rect 28408 9364 28414 9376
rect 28721 9367 28779 9373
rect 28721 9364 28733 9367
rect 28408 9336 28733 9364
rect 28408 9324 28414 9336
rect 28721 9333 28733 9336
rect 28767 9333 28779 9367
rect 28721 9327 28779 9333
rect 29178 9324 29184 9376
rect 29236 9364 29242 9376
rect 29917 9367 29975 9373
rect 29917 9364 29929 9367
rect 29236 9336 29929 9364
rect 29236 9324 29242 9336
rect 29917 9333 29929 9336
rect 29963 9333 29975 9367
rect 29917 9327 29975 9333
rect 30742 9324 30748 9376
rect 30800 9324 30806 9376
rect 31386 9324 31392 9376
rect 31444 9364 31450 9376
rect 32416 9364 32444 9472
rect 33689 9469 33701 9472
rect 33735 9469 33747 9503
rect 33689 9463 33747 9469
rect 34241 9503 34299 9509
rect 34241 9469 34253 9503
rect 34287 9469 34299 9503
rect 34241 9463 34299 9469
rect 34256 9432 34284 9463
rect 34974 9460 34980 9512
rect 35032 9460 35038 9512
rect 36354 9460 36360 9512
rect 36412 9500 36418 9512
rect 36541 9503 36599 9509
rect 36541 9500 36553 9503
rect 36412 9472 36553 9500
rect 36412 9460 36418 9472
rect 36541 9469 36553 9472
rect 36587 9469 36599 9503
rect 36541 9463 36599 9469
rect 37369 9503 37427 9509
rect 37369 9469 37381 9503
rect 37415 9500 37427 9503
rect 37918 9500 37924 9512
rect 37415 9472 37924 9500
rect 37415 9469 37427 9472
rect 37369 9463 37427 9469
rect 37918 9460 37924 9472
rect 37976 9460 37982 9512
rect 33152 9404 34284 9432
rect 31444 9336 32444 9364
rect 31444 9324 31450 9336
rect 32766 9324 32772 9376
rect 32824 9364 32830 9376
rect 33152 9364 33180 9404
rect 35066 9392 35072 9444
rect 35124 9432 35130 9444
rect 35342 9432 35348 9444
rect 35124 9404 35348 9432
rect 35124 9392 35130 9404
rect 35342 9392 35348 9404
rect 35400 9392 35406 9444
rect 35989 9435 36047 9441
rect 35989 9401 36001 9435
rect 36035 9432 36047 9435
rect 37090 9432 37096 9444
rect 36035 9404 37096 9432
rect 36035 9401 36047 9404
rect 35989 9395 36047 9401
rect 37090 9392 37096 9404
rect 37148 9392 37154 9444
rect 32824 9336 33180 9364
rect 33597 9367 33655 9373
rect 32824 9324 32830 9336
rect 33597 9333 33609 9367
rect 33643 9364 33655 9367
rect 34146 9364 34152 9376
rect 33643 9336 34152 9364
rect 33643 9333 33655 9336
rect 33597 9327 33655 9333
rect 34146 9324 34152 9336
rect 34204 9324 34210 9376
rect 35250 9324 35256 9376
rect 35308 9324 35314 9376
rect 36725 9367 36783 9373
rect 36725 9333 36737 9367
rect 36771 9364 36783 9367
rect 36998 9364 37004 9376
rect 36771 9336 37004 9364
rect 36771 9333 36783 9336
rect 36725 9327 36783 9333
rect 36998 9324 37004 9336
rect 37056 9324 37062 9376
rect 38194 9324 38200 9376
rect 38252 9324 38258 9376
rect 2024 9274 77924 9296
rect 2024 9222 5134 9274
rect 5186 9222 5198 9274
rect 5250 9222 5262 9274
rect 5314 9222 5326 9274
rect 5378 9222 5390 9274
rect 5442 9222 35854 9274
rect 35906 9222 35918 9274
rect 35970 9222 35982 9274
rect 36034 9222 36046 9274
rect 36098 9222 36110 9274
rect 36162 9222 66574 9274
rect 66626 9222 66638 9274
rect 66690 9222 66702 9274
rect 66754 9222 66766 9274
rect 66818 9222 66830 9274
rect 66882 9222 77924 9274
rect 2024 9200 77924 9222
rect 11790 9120 11796 9172
rect 11848 9120 11854 9172
rect 15930 9120 15936 9172
rect 15988 9160 15994 9172
rect 17221 9163 17279 9169
rect 17221 9160 17233 9163
rect 15988 9132 17233 9160
rect 15988 9120 15994 9132
rect 17221 9129 17233 9132
rect 17267 9129 17279 9163
rect 17221 9123 17279 9129
rect 17586 9120 17592 9172
rect 17644 9120 17650 9172
rect 17678 9120 17684 9172
rect 17736 9160 17742 9172
rect 17736 9132 21864 9160
rect 17736 9120 17742 9132
rect 18966 9052 18972 9104
rect 19024 9092 19030 9104
rect 19024 9064 21036 9092
rect 19024 9052 19030 9064
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 17313 9027 17371 9033
rect 17313 9024 17325 9027
rect 10928 8996 17325 9024
rect 10928 8984 10934 8996
rect 17313 8993 17325 8996
rect 17359 8993 17371 9027
rect 17313 8987 17371 8993
rect 17770 8984 17776 9036
rect 17828 9024 17834 9036
rect 21008 9033 21036 9064
rect 19337 9027 19395 9033
rect 19337 9024 19349 9027
rect 17828 8996 19349 9024
rect 17828 8984 17834 8996
rect 19337 8993 19349 8996
rect 19383 8993 19395 9027
rect 20993 9027 21051 9033
rect 19337 8987 19395 8993
rect 19444 8996 20484 9024
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 10008 8928 11897 8956
rect 10008 8916 10014 8928
rect 11885 8925 11897 8928
rect 11931 8925 11943 8959
rect 11885 8919 11943 8925
rect 17221 8959 17279 8965
rect 17221 8925 17233 8959
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 17236 8820 17264 8919
rect 17954 8916 17960 8968
rect 18012 8956 18018 8968
rect 19153 8959 19211 8965
rect 19153 8956 19165 8959
rect 18012 8928 19165 8956
rect 18012 8916 18018 8928
rect 19153 8925 19165 8928
rect 19199 8925 19211 8959
rect 19153 8919 19211 8925
rect 18046 8848 18052 8900
rect 18104 8848 18110 8900
rect 18138 8848 18144 8900
rect 18196 8888 18202 8900
rect 19444 8888 19472 8996
rect 19886 8916 19892 8968
rect 19944 8916 19950 8968
rect 20165 8959 20223 8965
rect 20165 8925 20177 8959
rect 20211 8925 20223 8959
rect 20165 8919 20223 8925
rect 18196 8860 19472 8888
rect 18196 8848 18202 8860
rect 19610 8848 19616 8900
rect 19668 8888 19674 8900
rect 20180 8888 20208 8919
rect 20254 8916 20260 8968
rect 20312 8956 20318 8968
rect 20349 8959 20407 8965
rect 20349 8956 20361 8959
rect 20312 8928 20361 8956
rect 20312 8916 20318 8928
rect 20349 8925 20361 8928
rect 20395 8925 20407 8959
rect 20456 8956 20484 8996
rect 20993 8993 21005 9027
rect 21039 8993 21051 9027
rect 20993 8987 21051 8993
rect 21729 8959 21787 8965
rect 21729 8956 21741 8959
rect 20456 8928 21741 8956
rect 20349 8919 20407 8925
rect 21729 8925 21741 8928
rect 21775 8925 21787 8959
rect 21836 8956 21864 9132
rect 23198 9120 23204 9172
rect 23256 9160 23262 9172
rect 23256 9132 25544 9160
rect 23256 9120 23262 9132
rect 21910 9052 21916 9104
rect 21968 9092 21974 9104
rect 23290 9092 23296 9104
rect 21968 9064 23296 9092
rect 21968 9052 21974 9064
rect 23290 9052 23296 9064
rect 23348 9052 23354 9104
rect 23400 9064 25452 9092
rect 22094 8984 22100 9036
rect 22152 9024 22158 9036
rect 22465 9027 22523 9033
rect 22465 9024 22477 9027
rect 22152 8996 22477 9024
rect 22152 8984 22158 8996
rect 22465 8993 22477 8996
rect 22511 8993 22523 9027
rect 22465 8987 22523 8993
rect 22922 8984 22928 9036
rect 22980 9024 22986 9036
rect 23400 9024 23428 9064
rect 22980 8996 23428 9024
rect 22980 8984 22986 8996
rect 23566 8984 23572 9036
rect 23624 8984 23630 9036
rect 21836 8928 23888 8956
rect 21729 8919 21787 8925
rect 19668 8860 20392 8888
rect 19668 8848 19674 8860
rect 18414 8820 18420 8832
rect 17236 8792 18420 8820
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 18598 8780 18604 8832
rect 18656 8780 18662 8832
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 20162 8820 20168 8832
rect 19576 8792 20168 8820
rect 19576 8780 19582 8792
rect 20162 8780 20168 8792
rect 20220 8780 20226 8832
rect 20254 8780 20260 8832
rect 20312 8780 20318 8832
rect 20364 8820 20392 8860
rect 20438 8848 20444 8900
rect 20496 8848 20502 8900
rect 20806 8888 20812 8900
rect 20656 8860 20812 8888
rect 20656 8820 20684 8860
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 21542 8848 21548 8900
rect 21600 8888 21606 8900
rect 23017 8891 23075 8897
rect 23017 8888 23029 8891
rect 21600 8860 23029 8888
rect 21600 8848 21606 8860
rect 23017 8857 23029 8860
rect 23063 8857 23075 8891
rect 23860 8888 23888 8928
rect 24302 8916 24308 8968
rect 24360 8916 24366 8968
rect 24486 8916 24492 8968
rect 24544 8916 24550 8968
rect 25130 8916 25136 8968
rect 25188 8956 25194 8968
rect 25317 8959 25375 8965
rect 25317 8956 25329 8959
rect 25188 8928 25329 8956
rect 25188 8916 25194 8928
rect 25317 8925 25329 8928
rect 25363 8925 25375 8959
rect 25424 8956 25452 9064
rect 25516 9024 25544 9132
rect 25682 9120 25688 9172
rect 25740 9160 25746 9172
rect 27801 9163 27859 9169
rect 27801 9160 27813 9163
rect 25740 9132 27813 9160
rect 25740 9120 25746 9132
rect 27801 9129 27813 9132
rect 27847 9129 27859 9163
rect 27801 9123 27859 9129
rect 28629 9163 28687 9169
rect 28629 9129 28641 9163
rect 28675 9160 28687 9163
rect 32858 9160 32864 9172
rect 28675 9132 32864 9160
rect 28675 9129 28687 9132
rect 28629 9123 28687 9129
rect 32858 9120 32864 9132
rect 32916 9160 32922 9172
rect 33134 9160 33140 9172
rect 32916 9132 33140 9160
rect 32916 9120 32922 9132
rect 33134 9120 33140 9132
rect 33192 9160 33198 9172
rect 33502 9160 33508 9172
rect 33192 9132 33508 9160
rect 33192 9120 33198 9132
rect 33502 9120 33508 9132
rect 33560 9120 33566 9172
rect 34333 9163 34391 9169
rect 34333 9129 34345 9163
rect 34379 9160 34391 9163
rect 35618 9160 35624 9172
rect 34379 9132 35624 9160
rect 34379 9129 34391 9132
rect 34333 9123 34391 9129
rect 35618 9120 35624 9132
rect 35676 9120 35682 9172
rect 25958 9052 25964 9104
rect 26016 9092 26022 9104
rect 31021 9095 31079 9101
rect 31021 9092 31033 9095
rect 26016 9064 31033 9092
rect 26016 9052 26022 9064
rect 31021 9061 31033 9064
rect 31067 9061 31079 9095
rect 31938 9092 31944 9104
rect 31021 9055 31079 9061
rect 31128 9064 31944 9092
rect 26237 9027 26295 9033
rect 26237 9024 26249 9027
rect 25516 8996 26249 9024
rect 26237 8993 26249 8996
rect 26283 8993 26295 9027
rect 26237 8987 26295 8993
rect 26973 9027 27031 9033
rect 26973 8993 26985 9027
rect 27019 9024 27031 9027
rect 27522 9024 27528 9036
rect 27019 8996 27528 9024
rect 27019 8993 27031 8996
rect 26973 8987 27031 8993
rect 27522 8984 27528 8996
rect 27580 8984 27586 9036
rect 28442 8984 28448 9036
rect 28500 9024 28506 9036
rect 28813 9027 28871 9033
rect 28813 9024 28825 9027
rect 28500 8996 28825 9024
rect 28500 8984 28506 8996
rect 28813 8993 28825 8996
rect 28859 8993 28871 9027
rect 28813 8987 28871 8993
rect 29270 8984 29276 9036
rect 29328 9024 29334 9036
rect 29365 9027 29423 9033
rect 29365 9024 29377 9027
rect 29328 8996 29377 9024
rect 29328 8984 29334 8996
rect 29365 8993 29377 8996
rect 29411 8993 29423 9027
rect 30466 9024 30472 9036
rect 29365 8987 29423 8993
rect 29472 8996 30472 9024
rect 26329 8959 26387 8965
rect 26329 8956 26341 8959
rect 25424 8928 26341 8956
rect 25317 8919 25375 8925
rect 26329 8925 26341 8928
rect 26375 8925 26387 8959
rect 26329 8919 26387 8925
rect 27706 8916 27712 8968
rect 27764 8916 27770 8968
rect 27985 8959 28043 8965
rect 27985 8925 27997 8959
rect 28031 8956 28043 8959
rect 29472 8956 29500 8996
rect 30466 8984 30472 8996
rect 30524 8984 30530 9036
rect 28031 8928 29500 8956
rect 28031 8925 28043 8928
rect 27985 8919 28043 8925
rect 29638 8916 29644 8968
rect 29696 8916 29702 8968
rect 31128 8956 31156 9064
rect 31938 9052 31944 9064
rect 31996 9052 32002 9104
rect 36078 9052 36084 9104
rect 36136 9092 36142 9104
rect 36446 9092 36452 9104
rect 36136 9064 36452 9092
rect 36136 9052 36142 9064
rect 36446 9052 36452 9064
rect 36504 9052 36510 9104
rect 31205 9027 31263 9033
rect 31205 8993 31217 9027
rect 31251 9024 31263 9027
rect 31573 9027 31631 9033
rect 31251 8996 31524 9024
rect 31251 8993 31263 8996
rect 31205 8987 31263 8993
rect 31297 8959 31355 8965
rect 31297 8956 31309 8959
rect 30484 8928 31309 8956
rect 30484 8900 30512 8928
rect 31297 8925 31309 8928
rect 31343 8925 31355 8959
rect 31496 8956 31524 8996
rect 31573 8993 31585 9027
rect 31619 9024 31631 9027
rect 32493 9027 32551 9033
rect 32493 9024 32505 9027
rect 31619 8996 32505 9024
rect 31619 8993 31631 8996
rect 31573 8987 31631 8993
rect 32493 8993 32505 8996
rect 32539 8993 32551 9027
rect 32493 8987 32551 8993
rect 34054 8984 34060 9036
rect 34112 9024 34118 9036
rect 34112 8996 35204 9024
rect 34112 8984 34118 8996
rect 31846 8956 31852 8968
rect 31496 8928 31852 8956
rect 31297 8919 31355 8925
rect 31846 8916 31852 8928
rect 31904 8916 31910 8968
rect 32398 8916 32404 8968
rect 32456 8916 32462 8968
rect 33134 8916 33140 8968
rect 33192 8916 33198 8968
rect 33965 8959 34023 8965
rect 33965 8925 33977 8959
rect 34011 8956 34023 8959
rect 34514 8956 34520 8968
rect 34011 8928 34520 8956
rect 34011 8925 34023 8928
rect 33965 8919 34023 8925
rect 34514 8916 34520 8928
rect 34572 8916 34578 8968
rect 34885 8959 34943 8965
rect 34885 8925 34897 8959
rect 34931 8956 34943 8959
rect 35066 8956 35072 8968
rect 34931 8928 35072 8956
rect 34931 8925 34943 8928
rect 34885 8919 34943 8925
rect 35066 8916 35072 8928
rect 35124 8916 35130 8968
rect 35176 8956 35204 8996
rect 35434 8984 35440 9036
rect 35492 9024 35498 9036
rect 36173 9027 36231 9033
rect 36173 9024 36185 9027
rect 35492 8996 36185 9024
rect 35492 8984 35498 8996
rect 36173 8993 36185 8996
rect 36219 8993 36231 9027
rect 36173 8987 36231 8993
rect 38013 9027 38071 9033
rect 38013 8993 38025 9027
rect 38059 9024 38071 9027
rect 38286 9024 38292 9036
rect 38059 8996 38292 9024
rect 38059 8993 38071 8996
rect 38013 8987 38071 8993
rect 38286 8984 38292 8996
rect 38344 8984 38350 9036
rect 36357 8959 36415 8965
rect 36357 8956 36369 8959
rect 35176 8928 36369 8956
rect 36357 8925 36369 8928
rect 36403 8925 36415 8959
rect 36357 8919 36415 8925
rect 36909 8959 36967 8965
rect 36909 8925 36921 8959
rect 36955 8925 36967 8959
rect 36909 8919 36967 8925
rect 25593 8891 25651 8897
rect 25593 8888 25605 8891
rect 23860 8860 25605 8888
rect 23017 8851 23075 8857
rect 25593 8857 25605 8860
rect 25639 8857 25651 8891
rect 25593 8851 25651 8857
rect 27430 8848 27436 8900
rect 27488 8888 27494 8900
rect 28077 8891 28135 8897
rect 28077 8888 28089 8891
rect 27488 8860 28089 8888
rect 27488 8848 27494 8860
rect 28077 8857 28089 8860
rect 28123 8857 28135 8891
rect 28077 8851 28135 8857
rect 28353 8891 28411 8897
rect 28353 8857 28365 8891
rect 28399 8888 28411 8891
rect 28994 8888 29000 8900
rect 28399 8860 29000 8888
rect 28399 8857 28411 8860
rect 28353 8851 28411 8857
rect 28994 8848 29000 8860
rect 29052 8848 29058 8900
rect 30466 8848 30472 8900
rect 30524 8848 30530 8900
rect 30837 8891 30895 8897
rect 30837 8857 30849 8891
rect 30883 8888 30895 8891
rect 31110 8888 31116 8900
rect 30883 8860 31116 8888
rect 30883 8857 30895 8860
rect 30837 8851 30895 8857
rect 31110 8848 31116 8860
rect 31168 8848 31174 8900
rect 31662 8848 31668 8900
rect 31720 8888 31726 8900
rect 31720 8860 33456 8888
rect 31720 8848 31726 8860
rect 20364 8792 20684 8820
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 21177 8823 21235 8829
rect 21177 8820 21189 8823
rect 20772 8792 21189 8820
rect 20772 8780 20778 8792
rect 21177 8789 21189 8792
rect 21223 8789 21235 8823
rect 21177 8783 21235 8789
rect 21450 8780 21456 8832
rect 21508 8820 21514 8832
rect 21913 8823 21971 8829
rect 21913 8820 21925 8823
rect 21508 8792 21925 8820
rect 21508 8780 21514 8792
rect 21913 8789 21925 8792
rect 21959 8789 21971 8823
rect 21913 8783 21971 8789
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 23753 8823 23811 8829
rect 23753 8820 23765 8823
rect 23532 8792 23765 8820
rect 23532 8780 23538 8792
rect 23753 8789 23765 8792
rect 23799 8789 23811 8823
rect 23753 8783 23811 8789
rect 25038 8780 25044 8832
rect 25096 8820 25102 8832
rect 25133 8823 25191 8829
rect 25133 8820 25145 8823
rect 25096 8792 25145 8820
rect 25096 8780 25102 8792
rect 25133 8789 25145 8792
rect 25179 8789 25191 8823
rect 25133 8783 25191 8789
rect 25222 8780 25228 8832
rect 25280 8820 25286 8832
rect 27065 8823 27123 8829
rect 27065 8820 27077 8823
rect 25280 8792 27077 8820
rect 25280 8780 25286 8792
rect 27065 8789 27077 8792
rect 27111 8789 27123 8823
rect 27065 8783 27123 8789
rect 27246 8780 27252 8832
rect 27304 8820 27310 8832
rect 28261 8823 28319 8829
rect 28261 8820 28273 8823
rect 27304 8792 28273 8820
rect 27304 8780 27310 8792
rect 28261 8789 28273 8792
rect 28307 8789 28319 8823
rect 28261 8783 28319 8789
rect 28442 8780 28448 8832
rect 28500 8780 28506 8832
rect 29362 8780 29368 8832
rect 29420 8820 29426 8832
rect 30285 8823 30343 8829
rect 30285 8820 30297 8823
rect 29420 8792 30297 8820
rect 29420 8780 29426 8792
rect 30285 8789 30297 8792
rect 30331 8789 30343 8823
rect 30285 8783 30343 8789
rect 31754 8780 31760 8832
rect 31812 8780 31818 8832
rect 31938 8780 31944 8832
rect 31996 8820 32002 8832
rect 32398 8820 32404 8832
rect 31996 8792 32404 8820
rect 31996 8780 32002 8792
rect 32398 8780 32404 8792
rect 32456 8780 32462 8832
rect 33318 8780 33324 8832
rect 33376 8780 33382 8832
rect 33428 8820 33456 8860
rect 33502 8848 33508 8900
rect 33560 8888 33566 8900
rect 36262 8888 36268 8900
rect 33560 8860 36268 8888
rect 33560 8848 33566 8860
rect 36262 8848 36268 8860
rect 36320 8848 36326 8900
rect 33870 8820 33876 8832
rect 33428 8792 33876 8820
rect 33870 8780 33876 8792
rect 33928 8780 33934 8832
rect 34514 8780 34520 8832
rect 34572 8820 34578 8832
rect 34977 8823 35035 8829
rect 34977 8820 34989 8823
rect 34572 8792 34989 8820
rect 34572 8780 34578 8792
rect 34977 8789 34989 8792
rect 35023 8789 35035 8823
rect 34977 8783 35035 8789
rect 35066 8780 35072 8832
rect 35124 8820 35130 8832
rect 35621 8823 35679 8829
rect 35621 8820 35633 8823
rect 35124 8792 35633 8820
rect 35124 8780 35130 8792
rect 35621 8789 35633 8792
rect 35667 8789 35679 8823
rect 35621 8783 35679 8789
rect 35710 8780 35716 8832
rect 35768 8820 35774 8832
rect 36924 8820 36952 8919
rect 37458 8916 37464 8968
rect 37516 8956 37522 8968
rect 38105 8959 38163 8965
rect 38105 8956 38117 8959
rect 37516 8928 38117 8956
rect 37516 8916 37522 8928
rect 38105 8925 38117 8928
rect 38151 8925 38163 8959
rect 38105 8919 38163 8925
rect 37366 8848 37372 8900
rect 37424 8848 37430 8900
rect 35768 8792 36952 8820
rect 35768 8780 35774 8792
rect 38654 8780 38660 8832
rect 38712 8780 38718 8832
rect 2024 8730 77924 8752
rect 2024 8678 5794 8730
rect 5846 8678 5858 8730
rect 5910 8678 5922 8730
rect 5974 8678 5986 8730
rect 6038 8678 6050 8730
rect 6102 8678 36514 8730
rect 36566 8678 36578 8730
rect 36630 8678 36642 8730
rect 36694 8678 36706 8730
rect 36758 8678 36770 8730
rect 36822 8678 67234 8730
rect 67286 8678 67298 8730
rect 67350 8678 67362 8730
rect 67414 8678 67426 8730
rect 67478 8678 67490 8730
rect 67542 8678 77924 8730
rect 2024 8656 77924 8678
rect 15102 8576 15108 8628
rect 15160 8616 15166 8628
rect 18138 8616 18144 8628
rect 15160 8588 18144 8616
rect 15160 8576 15166 8588
rect 18138 8576 18144 8588
rect 18196 8576 18202 8628
rect 19242 8576 19248 8628
rect 19300 8576 19306 8628
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 23017 8619 23075 8625
rect 23017 8616 23029 8619
rect 19484 8588 19932 8616
rect 19484 8576 19490 8588
rect 19904 8560 19932 8588
rect 19996 8588 23029 8616
rect 13906 8508 13912 8560
rect 13964 8548 13970 8560
rect 19705 8551 19763 8557
rect 19705 8548 19717 8551
rect 13964 8520 19717 8548
rect 13964 8508 13970 8520
rect 19705 8517 19717 8520
rect 19751 8517 19763 8551
rect 19705 8511 19763 8517
rect 19886 8508 19892 8560
rect 19944 8508 19950 8560
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 16025 8483 16083 8489
rect 16025 8480 16037 8483
rect 8260 8452 16037 8480
rect 8260 8440 8266 8452
rect 16025 8449 16037 8452
rect 16071 8449 16083 8483
rect 16025 8443 16083 8449
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 17865 8483 17923 8489
rect 17865 8480 17877 8483
rect 16172 8452 17877 8480
rect 16172 8440 16178 8452
rect 17865 8449 17877 8452
rect 17911 8449 17923 8483
rect 19996 8480 20024 8588
rect 23017 8585 23029 8588
rect 23063 8585 23075 8619
rect 23017 8579 23075 8585
rect 23290 8576 23296 8628
rect 23348 8616 23354 8628
rect 23348 8588 25636 8616
rect 23348 8576 23354 8588
rect 21910 8548 21916 8560
rect 17865 8443 17923 8449
rect 17972 8452 20024 8480
rect 20364 8520 21916 8548
rect 12894 8372 12900 8424
rect 12952 8412 12958 8424
rect 16761 8415 16819 8421
rect 12952 8384 16344 8412
rect 12952 8372 12958 8384
rect 3970 8304 3976 8356
rect 4028 8344 4034 8356
rect 15473 8347 15531 8353
rect 15473 8344 15485 8347
rect 4028 8316 15485 8344
rect 4028 8304 4034 8316
rect 15473 8313 15485 8316
rect 15519 8313 15531 8347
rect 15473 8307 15531 8313
rect 16316 8276 16344 8384
rect 16761 8381 16773 8415
rect 16807 8412 16819 8415
rect 17126 8412 17132 8424
rect 16807 8384 17132 8412
rect 16807 8381 16819 8384
rect 16761 8375 16819 8381
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 17972 8412 18000 8452
rect 17236 8384 18000 8412
rect 16390 8304 16396 8356
rect 16448 8344 16454 8356
rect 17236 8344 17264 8384
rect 18138 8372 18144 8424
rect 18196 8412 18202 8424
rect 18601 8415 18659 8421
rect 18601 8412 18613 8415
rect 18196 8384 18613 8412
rect 18196 8372 18202 8384
rect 18601 8381 18613 8384
rect 18647 8412 18659 8415
rect 18874 8412 18880 8424
rect 18647 8384 18880 8412
rect 18647 8381 18659 8384
rect 18601 8375 18659 8381
rect 18874 8372 18880 8384
rect 18932 8372 18938 8424
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 20257 8415 20315 8421
rect 20257 8412 20269 8415
rect 19392 8384 20269 8412
rect 19392 8372 19398 8384
rect 20257 8381 20269 8384
rect 20303 8381 20315 8415
rect 20257 8375 20315 8381
rect 16448 8316 17264 8344
rect 16448 8304 16454 8316
rect 17310 8304 17316 8356
rect 17368 8304 17374 8356
rect 18509 8347 18567 8353
rect 17420 8316 18460 8344
rect 17420 8276 17448 8316
rect 16316 8248 17448 8276
rect 18432 8276 18460 8316
rect 18509 8313 18521 8347
rect 18555 8344 18567 8347
rect 19242 8344 19248 8356
rect 18555 8316 19248 8344
rect 18555 8313 18567 8316
rect 18509 8307 18567 8313
rect 19242 8304 19248 8316
rect 19300 8304 19306 8356
rect 19426 8304 19432 8356
rect 19484 8304 19490 8356
rect 20364 8344 20392 8520
rect 21910 8508 21916 8520
rect 21968 8508 21974 8560
rect 22002 8508 22008 8560
rect 22060 8548 22066 8560
rect 23658 8548 23664 8560
rect 22060 8520 23664 8548
rect 22060 8508 22066 8520
rect 23658 8508 23664 8520
rect 23716 8548 23722 8560
rect 23716 8520 24794 8548
rect 23716 8508 23722 8520
rect 21634 8440 21640 8492
rect 21692 8480 21698 8492
rect 22094 8480 22100 8492
rect 21692 8452 22100 8480
rect 21692 8440 21698 8452
rect 22094 8440 22100 8452
rect 22152 8480 22158 8492
rect 22370 8480 22376 8492
rect 22152 8452 22376 8480
rect 22152 8440 22158 8452
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 25608 8480 25636 8588
rect 25774 8576 25780 8628
rect 25832 8616 25838 8628
rect 29638 8616 29644 8628
rect 25832 8588 29644 8616
rect 25832 8576 25838 8588
rect 29638 8576 29644 8588
rect 29696 8576 29702 8628
rect 30190 8576 30196 8628
rect 30248 8616 30254 8628
rect 30248 8588 32352 8616
rect 30248 8576 30254 8588
rect 25866 8508 25872 8560
rect 25924 8548 25930 8560
rect 26329 8551 26387 8557
rect 26329 8548 26341 8551
rect 25924 8520 26341 8548
rect 25924 8508 25930 8520
rect 26329 8517 26341 8520
rect 26375 8517 26387 8551
rect 26329 8511 26387 8517
rect 26878 8508 26884 8560
rect 26936 8548 26942 8560
rect 28905 8551 28963 8557
rect 28905 8548 28917 8551
rect 26936 8520 28917 8548
rect 26936 8508 26942 8520
rect 28905 8517 28917 8520
rect 28951 8517 28963 8551
rect 31665 8551 31723 8557
rect 31665 8548 31677 8551
rect 28905 8511 28963 8517
rect 29564 8520 30406 8548
rect 31220 8520 31677 8548
rect 27065 8483 27123 8489
rect 27065 8480 27077 8483
rect 25608 8452 27077 8480
rect 27065 8449 27077 8452
rect 27111 8449 27123 8483
rect 27065 8443 27123 8449
rect 27798 8440 27804 8492
rect 27856 8480 27862 8492
rect 27893 8483 27951 8489
rect 27893 8480 27905 8483
rect 27856 8452 27905 8480
rect 27856 8440 27862 8452
rect 27893 8449 27905 8452
rect 27939 8449 27951 8483
rect 27893 8443 27951 8449
rect 28077 8483 28135 8489
rect 28077 8449 28089 8483
rect 28123 8449 28135 8483
rect 28077 8443 28135 8449
rect 20438 8372 20444 8424
rect 20496 8372 20502 8424
rect 20806 8372 20812 8424
rect 20864 8412 20870 8424
rect 21729 8415 21787 8421
rect 21729 8412 21741 8415
rect 20864 8384 21741 8412
rect 20864 8372 20870 8384
rect 21729 8381 21741 8384
rect 21775 8381 21787 8415
rect 21729 8375 21787 8381
rect 21910 8372 21916 8424
rect 21968 8372 21974 8424
rect 23382 8372 23388 8424
rect 23440 8412 23446 8424
rect 23569 8415 23627 8421
rect 23569 8412 23581 8415
rect 23440 8384 23581 8412
rect 23440 8372 23446 8384
rect 23569 8381 23581 8384
rect 23615 8381 23627 8415
rect 23569 8375 23627 8381
rect 24026 8372 24032 8424
rect 24084 8372 24090 8424
rect 24302 8372 24308 8424
rect 24360 8372 24366 8424
rect 24670 8372 24676 8424
rect 24728 8412 24734 8424
rect 25682 8412 25688 8424
rect 24728 8384 25688 8412
rect 24728 8372 24734 8384
rect 25682 8372 25688 8384
rect 25740 8372 25746 8424
rect 26050 8372 26056 8424
rect 26108 8372 26114 8424
rect 26418 8372 26424 8424
rect 26476 8412 26482 8424
rect 26970 8412 26976 8424
rect 26476 8384 26976 8412
rect 26476 8372 26482 8384
rect 26970 8372 26976 8384
rect 27028 8372 27034 8424
rect 28092 8412 28120 8443
rect 27172 8384 28120 8412
rect 19536 8316 20392 8344
rect 19536 8276 19564 8316
rect 21082 8304 21088 8356
rect 21140 8304 21146 8356
rect 21174 8304 21180 8356
rect 21232 8304 21238 8356
rect 22296 8316 22692 8344
rect 18432 8248 19564 8276
rect 19794 8236 19800 8288
rect 19852 8276 19858 8288
rect 22296 8276 22324 8316
rect 19852 8248 22324 8276
rect 19852 8236 19858 8248
rect 22370 8236 22376 8288
rect 22428 8276 22434 8288
rect 22557 8279 22615 8285
rect 22557 8276 22569 8279
rect 22428 8248 22569 8276
rect 22428 8236 22434 8248
rect 22557 8245 22569 8248
rect 22603 8245 22615 8279
rect 22664 8276 22692 8316
rect 23750 8304 23756 8356
rect 23808 8344 23814 8356
rect 23808 8316 24164 8344
rect 23808 8304 23814 8316
rect 23934 8276 23940 8288
rect 22664 8248 23940 8276
rect 22557 8239 22615 8245
rect 23934 8236 23940 8248
rect 23992 8236 23998 8288
rect 24136 8276 24164 8316
rect 25590 8304 25596 8356
rect 25648 8344 25654 8356
rect 27172 8344 27200 8384
rect 28166 8372 28172 8424
rect 28224 8372 28230 8424
rect 28813 8415 28871 8421
rect 28813 8381 28825 8415
rect 28859 8412 28871 8415
rect 29457 8415 29515 8421
rect 29457 8412 29469 8415
rect 28859 8384 29469 8412
rect 28859 8381 28871 8384
rect 28813 8375 28871 8381
rect 29457 8381 29469 8384
rect 29503 8381 29515 8415
rect 29457 8375 29515 8381
rect 25648 8316 27200 8344
rect 25648 8304 25654 8316
rect 27246 8304 27252 8356
rect 27304 8344 27310 8356
rect 27709 8347 27767 8353
rect 27709 8344 27721 8347
rect 27304 8316 27721 8344
rect 27304 8304 27310 8316
rect 27709 8313 27721 8316
rect 27755 8313 27767 8347
rect 27709 8307 27767 8313
rect 27890 8304 27896 8356
rect 27948 8304 27954 8356
rect 28074 8304 28080 8356
rect 28132 8344 28138 8356
rect 29564 8344 29592 8520
rect 31220 8480 31248 8520
rect 31665 8517 31677 8520
rect 31711 8517 31723 8551
rect 31665 8511 31723 8517
rect 31128 8452 31248 8480
rect 31757 8483 31815 8489
rect 29638 8372 29644 8424
rect 29696 8372 29702 8424
rect 29914 8372 29920 8424
rect 29972 8372 29978 8424
rect 30650 8372 30656 8424
rect 30708 8412 30714 8424
rect 31128 8412 31156 8452
rect 31757 8449 31769 8483
rect 31803 8480 31815 8483
rect 31938 8480 31944 8492
rect 31803 8452 31944 8480
rect 31803 8449 31815 8452
rect 31757 8443 31815 8449
rect 31938 8440 31944 8452
rect 31996 8440 32002 8492
rect 30708 8384 31156 8412
rect 30708 8372 30714 8384
rect 32214 8372 32220 8424
rect 32272 8372 32278 8424
rect 32324 8412 32352 8588
rect 32398 8576 32404 8628
rect 32456 8616 32462 8628
rect 33229 8619 33287 8625
rect 33229 8616 33241 8619
rect 32456 8588 33241 8616
rect 32456 8576 32462 8588
rect 33229 8585 33241 8588
rect 33275 8585 33287 8619
rect 33965 8619 34023 8625
rect 33229 8579 33287 8585
rect 33612 8588 33916 8616
rect 32861 8551 32919 8557
rect 32861 8517 32873 8551
rect 32907 8548 32919 8551
rect 33134 8548 33140 8560
rect 32907 8520 33140 8548
rect 32907 8517 32919 8520
rect 32861 8511 32919 8517
rect 33134 8508 33140 8520
rect 33192 8508 33198 8560
rect 33042 8440 33048 8492
rect 33100 8440 33106 8492
rect 33229 8483 33287 8489
rect 33229 8480 33241 8483
rect 33152 8452 33241 8480
rect 32398 8412 32404 8424
rect 32324 8384 32404 8412
rect 32398 8372 32404 8384
rect 32456 8412 32462 8424
rect 33152 8412 33180 8452
rect 33229 8449 33241 8452
rect 33275 8449 33287 8483
rect 33229 8443 33287 8449
rect 33502 8440 33508 8492
rect 33560 8440 33566 8492
rect 33612 8489 33640 8588
rect 33888 8548 33916 8588
rect 33965 8585 33977 8619
rect 34011 8616 34023 8619
rect 34011 8588 36952 8616
rect 34011 8585 34023 8588
rect 33965 8579 34023 8585
rect 34146 8548 34152 8560
rect 33888 8520 34152 8548
rect 34146 8508 34152 8520
rect 34204 8548 34210 8560
rect 34790 8548 34796 8560
rect 34204 8520 34796 8548
rect 34204 8508 34210 8520
rect 34790 8508 34796 8520
rect 34848 8508 34854 8560
rect 35066 8508 35072 8560
rect 35124 8508 35130 8560
rect 33597 8483 33655 8489
rect 33597 8449 33609 8483
rect 33643 8449 33655 8483
rect 33597 8443 33655 8449
rect 33778 8440 33784 8492
rect 33836 8440 33842 8492
rect 33870 8440 33876 8492
rect 33928 8480 33934 8492
rect 34422 8480 34428 8492
rect 33928 8452 34428 8480
rect 33928 8440 33934 8452
rect 34422 8440 34428 8452
rect 34480 8440 34486 8492
rect 36078 8440 36084 8492
rect 36136 8480 36142 8492
rect 36722 8480 36728 8492
rect 36136 8452 36728 8480
rect 36136 8440 36142 8452
rect 36722 8440 36728 8452
rect 36780 8440 36786 8492
rect 36924 8489 36952 8588
rect 36909 8483 36967 8489
rect 36909 8449 36921 8483
rect 36955 8449 36967 8483
rect 36909 8443 36967 8449
rect 32456 8384 33180 8412
rect 33244 8384 34192 8412
rect 32456 8372 32462 8384
rect 28132 8316 29592 8344
rect 28132 8304 28138 8316
rect 26694 8276 26700 8288
rect 24136 8248 26700 8276
rect 26694 8236 26700 8248
rect 26752 8236 26758 8288
rect 29564 8276 29592 8316
rect 31110 8304 31116 8356
rect 31168 8344 31174 8356
rect 33244 8344 33272 8384
rect 34164 8356 34192 8384
rect 34606 8372 34612 8424
rect 34664 8372 34670 8424
rect 34793 8415 34851 8421
rect 34793 8381 34805 8415
rect 34839 8381 34851 8415
rect 34793 8375 34851 8381
rect 31168 8316 33272 8344
rect 33689 8347 33747 8353
rect 31168 8304 31174 8316
rect 33689 8313 33701 8347
rect 33735 8344 33747 8347
rect 33870 8344 33876 8356
rect 33735 8316 33876 8344
rect 33735 8313 33747 8316
rect 33689 8307 33747 8313
rect 33870 8304 33876 8316
rect 33928 8304 33934 8356
rect 34146 8304 34152 8356
rect 34204 8344 34210 8356
rect 34808 8344 34836 8375
rect 35066 8372 35072 8424
rect 35124 8412 35130 8424
rect 35710 8412 35716 8424
rect 35124 8384 35716 8412
rect 35124 8372 35130 8384
rect 35710 8372 35716 8384
rect 35768 8372 35774 8424
rect 35802 8372 35808 8424
rect 35860 8412 35866 8424
rect 36817 8415 36875 8421
rect 36817 8412 36829 8415
rect 35860 8384 36829 8412
rect 35860 8372 35866 8384
rect 36817 8381 36829 8384
rect 36863 8381 36875 8415
rect 36817 8375 36875 8381
rect 37182 8372 37188 8424
rect 37240 8412 37246 8424
rect 38749 8415 38807 8421
rect 38749 8412 38761 8415
rect 37240 8384 38761 8412
rect 37240 8372 37246 8384
rect 38749 8381 38761 8384
rect 38795 8381 38807 8415
rect 38749 8375 38807 8381
rect 39298 8372 39304 8424
rect 39356 8372 39362 8424
rect 39945 8415 40003 8421
rect 39945 8381 39957 8415
rect 39991 8412 40003 8415
rect 40221 8415 40279 8421
rect 40221 8412 40233 8415
rect 39991 8384 40233 8412
rect 39991 8381 40003 8384
rect 39945 8375 40003 8381
rect 40221 8381 40233 8384
rect 40267 8381 40279 8415
rect 40221 8375 40279 8381
rect 34204 8316 34836 8344
rect 34204 8304 34210 8316
rect 37642 8304 37648 8356
rect 37700 8344 37706 8356
rect 38197 8347 38255 8353
rect 38197 8344 38209 8347
rect 37700 8316 38209 8344
rect 37700 8304 37706 8316
rect 38197 8313 38209 8316
rect 38243 8313 38255 8347
rect 38197 8307 38255 8313
rect 40865 8347 40923 8353
rect 40865 8313 40877 8347
rect 40911 8344 40923 8347
rect 41414 8344 41420 8356
rect 40911 8316 41420 8344
rect 40911 8313 40923 8316
rect 40865 8307 40923 8313
rect 41414 8304 41420 8316
rect 41472 8304 41478 8356
rect 31202 8276 31208 8288
rect 29564 8248 31208 8276
rect 31202 8236 31208 8248
rect 31260 8236 31266 8288
rect 31662 8236 31668 8288
rect 31720 8276 31726 8288
rect 31941 8279 31999 8285
rect 31941 8276 31953 8279
rect 31720 8248 31953 8276
rect 31720 8236 31726 8248
rect 31941 8245 31953 8248
rect 31987 8245 31999 8279
rect 31941 8239 31999 8245
rect 33318 8236 33324 8288
rect 33376 8276 33382 8288
rect 34057 8279 34115 8285
rect 34057 8276 34069 8279
rect 33376 8248 34069 8276
rect 33376 8236 33382 8248
rect 34057 8245 34069 8248
rect 34103 8245 34115 8279
rect 34057 8239 34115 8245
rect 37550 8236 37556 8288
rect 37608 8236 37614 8288
rect 2024 8186 77924 8208
rect 2024 8134 5134 8186
rect 5186 8134 5198 8186
rect 5250 8134 5262 8186
rect 5314 8134 5326 8186
rect 5378 8134 5390 8186
rect 5442 8134 35854 8186
rect 35906 8134 35918 8186
rect 35970 8134 35982 8186
rect 36034 8134 36046 8186
rect 36098 8134 36110 8186
rect 36162 8134 66574 8186
rect 66626 8134 66638 8186
rect 66690 8134 66702 8186
rect 66754 8134 66766 8186
rect 66818 8134 66830 8186
rect 66882 8134 77924 8186
rect 2024 8112 77924 8134
rect 16669 8075 16727 8081
rect 16669 8041 16681 8075
rect 16715 8072 16727 8075
rect 17954 8072 17960 8084
rect 16715 8044 17960 8072
rect 16715 8041 16727 8044
rect 16669 8035 16727 8041
rect 17954 8032 17960 8044
rect 18012 8032 18018 8084
rect 18141 8075 18199 8081
rect 18141 8041 18153 8075
rect 18187 8072 18199 8075
rect 19150 8072 19156 8084
rect 18187 8044 19156 8072
rect 18187 8041 18199 8044
rect 18141 8035 18199 8041
rect 19150 8032 19156 8044
rect 19208 8032 19214 8084
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 19794 8072 19800 8084
rect 19659 8044 19800 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 19794 8032 19800 8044
rect 19852 8032 19858 8084
rect 21085 8075 21143 8081
rect 21085 8041 21097 8075
rect 21131 8072 21143 8075
rect 21910 8072 21916 8084
rect 21131 8044 21916 8072
rect 21131 8041 21143 8044
rect 21085 8035 21143 8041
rect 21910 8032 21916 8044
rect 21968 8032 21974 8084
rect 22186 8072 22192 8084
rect 22066 8044 22192 8072
rect 22066 8004 22094 8044
rect 22186 8032 22192 8044
rect 22244 8032 22250 8084
rect 22462 8032 22468 8084
rect 22520 8072 22526 8084
rect 26329 8075 26387 8081
rect 26329 8072 26341 8075
rect 22520 8044 26341 8072
rect 22520 8032 22526 8044
rect 26329 8041 26341 8044
rect 26375 8041 26387 8075
rect 26329 8035 26387 8041
rect 26510 8032 26516 8084
rect 26568 8072 26574 8084
rect 27065 8075 27123 8081
rect 27065 8072 27077 8075
rect 26568 8044 27077 8072
rect 26568 8032 26574 8044
rect 27065 8041 27077 8044
rect 27111 8041 27123 8075
rect 27065 8035 27123 8041
rect 27522 8032 27528 8084
rect 27580 8072 27586 8084
rect 27580 8044 29868 8072
rect 27580 8032 27586 8044
rect 20456 7976 22094 8004
rect 11146 7896 11152 7948
rect 11204 7936 11210 7948
rect 17497 7939 17555 7945
rect 17497 7936 17509 7939
rect 11204 7908 17509 7936
rect 11204 7896 11210 7908
rect 17497 7905 17509 7908
rect 17543 7905 17555 7939
rect 17497 7899 17555 7905
rect 18322 7896 18328 7948
rect 18380 7936 18386 7948
rect 18969 7939 19027 7945
rect 18969 7936 18981 7939
rect 18380 7908 18981 7936
rect 18380 7896 18386 7908
rect 18969 7905 18981 7908
rect 19015 7936 19027 7939
rect 19426 7936 19432 7948
rect 19015 7908 19432 7936
rect 19015 7905 19027 7908
rect 18969 7899 19027 7905
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 14829 7871 14887 7877
rect 14829 7868 14841 7871
rect 6972 7840 14841 7868
rect 6972 7828 6978 7840
rect 14829 7837 14841 7840
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 15378 7828 15384 7880
rect 15436 7828 15442 7880
rect 16298 7828 16304 7880
rect 16356 7828 16362 7880
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7868 17279 7871
rect 17402 7868 17408 7880
rect 17267 7840 17408 7868
rect 17267 7837 17279 7840
rect 17221 7831 17279 7837
rect 17402 7828 17408 7840
rect 17460 7828 17466 7880
rect 18782 7828 18788 7880
rect 18840 7828 18846 7880
rect 20456 7877 20484 7976
rect 23566 7964 23572 8016
rect 23624 8004 23630 8016
rect 23934 8004 23940 8016
rect 23624 7976 23940 8004
rect 23624 7964 23630 7976
rect 23934 7964 23940 7976
rect 23992 7964 23998 8016
rect 24210 7964 24216 8016
rect 24268 7964 24274 8016
rect 24397 8007 24455 8013
rect 24397 7973 24409 8007
rect 24443 8004 24455 8007
rect 24762 8004 24768 8016
rect 24443 7976 24768 8004
rect 24443 7973 24455 7976
rect 24397 7967 24455 7973
rect 24762 7964 24768 7976
rect 24820 7964 24826 8016
rect 25498 7964 25504 8016
rect 25556 8004 25562 8016
rect 28077 8007 28135 8013
rect 28077 8004 28089 8007
rect 25556 7976 28089 8004
rect 25556 7964 25562 7976
rect 28077 7973 28089 7976
rect 28123 8004 28135 8007
rect 28258 8004 28264 8016
rect 28123 7976 28264 8004
rect 28123 7973 28135 7976
rect 28077 7967 28135 7973
rect 28258 7964 28264 7976
rect 28316 7964 28322 8016
rect 29546 7964 29552 8016
rect 29604 7964 29610 8016
rect 21634 7936 21640 7948
rect 20732 7908 21640 7936
rect 20732 7877 20760 7908
rect 21634 7896 21640 7908
rect 21692 7896 21698 7948
rect 21726 7896 21732 7948
rect 21784 7896 21790 7948
rect 22097 7939 22155 7945
rect 22097 7905 22109 7939
rect 22143 7936 22155 7939
rect 24026 7936 24032 7948
rect 22143 7908 24032 7936
rect 22143 7905 22155 7908
rect 22097 7899 22155 7905
rect 24026 7896 24032 7908
rect 24084 7896 24090 7948
rect 24118 7896 24124 7948
rect 24176 7896 24182 7948
rect 24228 7936 24256 7964
rect 24228 7908 24440 7936
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 20625 7871 20683 7877
rect 20625 7837 20637 7871
rect 20671 7837 20683 7871
rect 20625 7831 20683 7837
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7837 20775 7871
rect 20717 7831 20775 7837
rect 20809 7871 20867 7877
rect 20809 7837 20821 7871
rect 20855 7868 20867 7871
rect 21177 7871 21235 7877
rect 21177 7868 21189 7871
rect 20855 7840 21189 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 21177 7837 21189 7840
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 18598 7760 18604 7812
rect 18656 7800 18662 7812
rect 20640 7800 20668 7831
rect 23934 7828 23940 7880
rect 23992 7868 23998 7880
rect 24412 7877 24440 7908
rect 25866 7896 25872 7948
rect 25924 7936 25930 7948
rect 26237 7939 26295 7945
rect 26237 7936 26249 7939
rect 25924 7908 26249 7936
rect 25924 7896 25930 7908
rect 26237 7905 26249 7908
rect 26283 7905 26295 7939
rect 26237 7899 26295 7905
rect 26694 7896 26700 7948
rect 26752 7936 26758 7948
rect 26752 7908 27936 7936
rect 26752 7896 26758 7908
rect 24213 7871 24271 7877
rect 24213 7868 24225 7871
rect 23992 7840 24225 7868
rect 23992 7828 23998 7840
rect 24213 7837 24225 7840
rect 24259 7837 24271 7871
rect 24213 7831 24271 7837
rect 24397 7871 24455 7877
rect 24397 7837 24409 7871
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 25038 7828 25044 7880
rect 25096 7868 25102 7880
rect 26050 7868 26056 7880
rect 25096 7840 26056 7868
rect 25096 7828 25102 7840
rect 26050 7828 26056 7840
rect 26108 7828 26114 7880
rect 26973 7871 27031 7877
rect 26973 7837 26985 7871
rect 27019 7868 27031 7871
rect 27522 7868 27528 7880
rect 27019 7840 27528 7868
rect 27019 7837 27031 7840
rect 26973 7831 27031 7837
rect 27522 7828 27528 7840
rect 27580 7828 27586 7880
rect 27614 7828 27620 7880
rect 27672 7828 27678 7880
rect 27798 7828 27804 7880
rect 27856 7828 27862 7880
rect 27908 7868 27936 7908
rect 28810 7896 28816 7948
rect 28868 7896 28874 7948
rect 28905 7939 28963 7945
rect 28905 7905 28917 7939
rect 28951 7936 28963 7939
rect 29086 7936 29092 7948
rect 28951 7908 29092 7936
rect 28951 7905 28963 7908
rect 28905 7899 28963 7905
rect 29086 7896 29092 7908
rect 29144 7896 29150 7948
rect 29840 7936 29868 8044
rect 29914 8032 29920 8084
rect 29972 8072 29978 8084
rect 30285 8075 30343 8081
rect 30285 8072 30297 8075
rect 29972 8044 30297 8072
rect 29972 8032 29978 8044
rect 30285 8041 30297 8044
rect 30331 8041 30343 8075
rect 30285 8035 30343 8041
rect 30374 8032 30380 8084
rect 30432 8072 30438 8084
rect 30469 8075 30527 8081
rect 30469 8072 30481 8075
rect 30432 8044 30481 8072
rect 30432 8032 30438 8044
rect 30469 8041 30481 8044
rect 30515 8041 30527 8075
rect 34701 8075 34759 8081
rect 34701 8072 34713 8075
rect 30469 8035 30527 8041
rect 30576 8044 34713 8072
rect 30190 7964 30196 8016
rect 30248 8004 30254 8016
rect 30576 8004 30604 8044
rect 34701 8041 34713 8044
rect 34747 8041 34759 8075
rect 34701 8035 34759 8041
rect 34882 8032 34888 8084
rect 34940 8072 34946 8084
rect 35621 8075 35679 8081
rect 35621 8072 35633 8075
rect 34940 8044 35633 8072
rect 34940 8032 34946 8044
rect 35621 8041 35633 8044
rect 35667 8041 35679 8075
rect 35621 8035 35679 8041
rect 37550 8032 37556 8084
rect 37608 8072 37614 8084
rect 37749 8075 37807 8081
rect 37749 8072 37761 8075
rect 37608 8044 37761 8072
rect 37608 8032 37614 8044
rect 37749 8041 37761 8044
rect 37795 8041 37807 8075
rect 37749 8035 37807 8041
rect 30248 7976 30604 8004
rect 30248 7964 30254 7976
rect 30834 7964 30840 8016
rect 30892 8004 30898 8016
rect 31757 8007 31815 8013
rect 31757 8004 31769 8007
rect 30892 7976 31769 8004
rect 30892 7964 30898 7976
rect 31757 7973 31769 7976
rect 31803 7973 31815 8007
rect 31757 7967 31815 7973
rect 33502 7936 33508 7948
rect 29840 7908 31892 7936
rect 28077 7871 28135 7877
rect 28077 7868 28089 7871
rect 27908 7840 28089 7868
rect 18656 7772 20668 7800
rect 18656 7760 18662 7772
rect 22370 7760 22376 7812
rect 22428 7760 22434 7812
rect 23658 7800 23664 7812
rect 23598 7772 23664 7800
rect 23658 7760 23664 7772
rect 23716 7760 23722 7812
rect 24489 7803 24547 7809
rect 24489 7800 24501 7803
rect 23768 7772 24501 7800
rect 10226 7692 10232 7744
rect 10284 7732 10290 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 10284 7704 14657 7732
rect 10284 7692 10290 7704
rect 14645 7701 14657 7704
rect 14691 7701 14703 7735
rect 14645 7695 14703 7701
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 15749 7735 15807 7741
rect 15749 7732 15761 7735
rect 14884 7704 15761 7732
rect 14884 7692 14890 7704
rect 15749 7701 15761 7704
rect 15795 7701 15807 7735
rect 15749 7695 15807 7701
rect 18230 7692 18236 7744
rect 18288 7692 18294 7744
rect 19794 7692 19800 7744
rect 19852 7692 19858 7744
rect 21818 7692 21824 7744
rect 21876 7732 21882 7744
rect 23768 7732 23796 7772
rect 24489 7769 24501 7772
rect 24535 7769 24547 7803
rect 24489 7763 24547 7769
rect 25682 7760 25688 7812
rect 25740 7800 25746 7812
rect 27816 7800 27844 7828
rect 25740 7772 27844 7800
rect 28000 7800 28028 7840
rect 28077 7837 28089 7840
rect 28123 7837 28135 7871
rect 28077 7831 28135 7837
rect 28534 7828 28540 7880
rect 28592 7868 28598 7880
rect 29641 7871 29699 7877
rect 29641 7868 29653 7871
rect 28592 7840 29653 7868
rect 28592 7828 28598 7840
rect 29641 7837 29653 7840
rect 29687 7837 29699 7871
rect 29641 7831 29699 7837
rect 30650 7828 30656 7880
rect 30708 7828 30714 7880
rect 30852 7877 30880 7908
rect 30837 7871 30895 7877
rect 30837 7837 30849 7871
rect 30883 7837 30895 7871
rect 30837 7831 30895 7837
rect 30929 7871 30987 7877
rect 30929 7837 30941 7871
rect 30975 7868 30987 7871
rect 31202 7868 31208 7880
rect 30975 7840 31208 7868
rect 30975 7837 30987 7840
rect 30929 7831 30987 7837
rect 31202 7828 31208 7840
rect 31260 7828 31266 7880
rect 31386 7828 31392 7880
rect 31444 7868 31450 7880
rect 31573 7871 31631 7877
rect 31573 7868 31585 7871
rect 31444 7840 31585 7868
rect 31444 7828 31450 7840
rect 31573 7837 31585 7840
rect 31619 7837 31631 7871
rect 31573 7831 31631 7837
rect 31754 7828 31760 7880
rect 31812 7828 31818 7880
rect 31864 7877 31892 7908
rect 32048 7908 33508 7936
rect 31849 7871 31907 7877
rect 31849 7837 31861 7871
rect 31895 7837 31907 7871
rect 31849 7831 31907 7837
rect 29546 7800 29552 7812
rect 28000 7772 29552 7800
rect 25740 7760 25746 7772
rect 29546 7760 29552 7772
rect 29604 7760 29610 7812
rect 29914 7760 29920 7812
rect 29972 7800 29978 7812
rect 31021 7803 31079 7809
rect 31021 7800 31033 7803
rect 29972 7772 31033 7800
rect 29972 7760 29978 7772
rect 31021 7769 31033 7772
rect 31067 7769 31079 7803
rect 31220 7800 31248 7828
rect 32048 7809 32076 7908
rect 33502 7896 33508 7908
rect 33560 7896 33566 7948
rect 33870 7896 33876 7948
rect 33928 7896 33934 7948
rect 34146 7896 34152 7948
rect 34204 7896 34210 7948
rect 38657 7939 38715 7945
rect 38657 7936 38669 7939
rect 36004 7908 38669 7936
rect 34241 7871 34299 7877
rect 34241 7837 34253 7871
rect 34287 7837 34299 7871
rect 34241 7831 34299 7837
rect 32033 7803 32091 7809
rect 32033 7800 32045 7803
rect 31220 7772 32045 7800
rect 31021 7763 31079 7769
rect 32033 7769 32045 7772
rect 32079 7769 32091 7803
rect 32033 7763 32091 7769
rect 32125 7803 32183 7809
rect 32125 7769 32137 7803
rect 32171 7769 32183 7803
rect 32125 7763 32183 7769
rect 21876 7704 23796 7732
rect 21876 7692 21882 7704
rect 24762 7692 24768 7744
rect 24820 7732 24826 7744
rect 25593 7735 25651 7741
rect 25593 7732 25605 7735
rect 24820 7704 25605 7732
rect 24820 7692 24826 7704
rect 25593 7701 25605 7704
rect 25639 7701 25651 7735
rect 25593 7695 25651 7701
rect 27154 7692 27160 7744
rect 27212 7732 27218 7744
rect 27893 7735 27951 7741
rect 27893 7732 27905 7735
rect 27212 7704 27905 7732
rect 27212 7692 27218 7704
rect 27893 7701 27905 7704
rect 27939 7701 27951 7735
rect 27893 7695 27951 7701
rect 27982 7692 27988 7744
rect 28040 7732 28046 7744
rect 28169 7735 28227 7741
rect 28169 7732 28181 7735
rect 28040 7704 28181 7732
rect 28040 7692 28046 7704
rect 28169 7701 28181 7704
rect 28215 7701 28227 7735
rect 28169 7695 28227 7701
rect 29086 7692 29092 7744
rect 29144 7732 29150 7744
rect 30190 7732 30196 7744
rect 29144 7704 30196 7732
rect 29144 7692 29150 7704
rect 30190 7692 30196 7704
rect 30248 7692 30254 7744
rect 30282 7692 30288 7744
rect 30340 7732 30346 7744
rect 30834 7732 30840 7744
rect 30340 7704 30840 7732
rect 30340 7692 30346 7704
rect 30834 7692 30840 7704
rect 30892 7692 30898 7744
rect 31386 7692 31392 7744
rect 31444 7732 31450 7744
rect 32140 7732 32168 7763
rect 32398 7760 32404 7812
rect 32456 7800 32462 7812
rect 32456 7772 32706 7800
rect 32456 7760 32462 7772
rect 31444 7704 32168 7732
rect 31444 7692 31450 7704
rect 32306 7692 32312 7744
rect 32364 7732 32370 7744
rect 34256 7732 34284 7831
rect 34330 7828 34336 7880
rect 34388 7868 34394 7880
rect 34517 7871 34575 7877
rect 34517 7868 34529 7871
rect 34388 7840 34529 7868
rect 34388 7828 34394 7840
rect 34517 7837 34529 7840
rect 34563 7837 34575 7871
rect 34517 7831 34575 7837
rect 34790 7828 34796 7880
rect 34848 7828 34854 7880
rect 34882 7828 34888 7880
rect 34940 7868 34946 7880
rect 35621 7871 35679 7877
rect 35621 7868 35633 7871
rect 34940 7840 35633 7868
rect 34940 7828 34946 7840
rect 35621 7837 35633 7840
rect 35667 7837 35679 7871
rect 35621 7831 35679 7837
rect 35805 7871 35863 7877
rect 35805 7837 35817 7871
rect 35851 7837 35863 7871
rect 35805 7831 35863 7837
rect 34422 7760 34428 7812
rect 34480 7800 34486 7812
rect 35820 7800 35848 7831
rect 36004 7812 36032 7908
rect 38657 7905 38669 7908
rect 38703 7905 38715 7939
rect 38657 7899 38715 7905
rect 40037 7939 40095 7945
rect 40037 7905 40049 7939
rect 40083 7936 40095 7939
rect 40402 7936 40408 7948
rect 40083 7908 40408 7936
rect 40083 7905 40095 7908
rect 40037 7899 40095 7905
rect 40402 7896 40408 7908
rect 40460 7896 40466 7948
rect 38013 7871 38071 7877
rect 38013 7837 38025 7871
rect 38059 7868 38071 7871
rect 38194 7868 38200 7880
rect 38059 7840 38200 7868
rect 38059 7837 38071 7840
rect 38013 7831 38071 7837
rect 38194 7828 38200 7840
rect 38252 7828 38258 7880
rect 40313 7871 40371 7877
rect 40313 7837 40325 7871
rect 40359 7837 40371 7871
rect 40313 7831 40371 7837
rect 40589 7871 40647 7877
rect 40589 7837 40601 7871
rect 40635 7868 40647 7871
rect 41598 7868 41604 7880
rect 40635 7840 41604 7868
rect 40635 7837 40647 7840
rect 40589 7831 40647 7837
rect 34480 7772 35848 7800
rect 34480 7760 34486 7772
rect 35986 7760 35992 7812
rect 36044 7760 36050 7812
rect 38378 7800 38384 7812
rect 37306 7772 38384 7800
rect 32364 7704 34284 7732
rect 32364 7692 32370 7704
rect 34330 7692 34336 7744
rect 34388 7692 34394 7744
rect 35437 7735 35495 7741
rect 35437 7701 35449 7735
rect 35483 7732 35495 7735
rect 35618 7732 35624 7744
rect 35483 7704 35624 7732
rect 35483 7701 35495 7704
rect 35437 7695 35495 7701
rect 35618 7692 35624 7704
rect 35676 7692 35682 7744
rect 36722 7692 36728 7744
rect 36780 7732 36786 7744
rect 37384 7732 37412 7772
rect 38378 7760 38384 7772
rect 38436 7760 38442 7812
rect 40328 7800 40356 7831
rect 41598 7828 41604 7840
rect 41656 7828 41662 7880
rect 40862 7800 40868 7812
rect 40328 7772 40868 7800
rect 40862 7760 40868 7772
rect 40920 7760 40926 7812
rect 36780 7704 37412 7732
rect 36780 7692 36786 7704
rect 37458 7692 37464 7744
rect 37516 7732 37522 7744
rect 38105 7735 38163 7741
rect 38105 7732 38117 7735
rect 37516 7704 38117 7732
rect 37516 7692 37522 7704
rect 38105 7701 38117 7704
rect 38151 7701 38163 7735
rect 38105 7695 38163 7701
rect 39206 7692 39212 7744
rect 39264 7732 39270 7744
rect 39393 7735 39451 7741
rect 39393 7732 39405 7735
rect 39264 7704 39405 7732
rect 39264 7692 39270 7704
rect 39393 7701 39405 7704
rect 39439 7701 39451 7735
rect 39393 7695 39451 7701
rect 40126 7692 40132 7744
rect 40184 7692 40190 7744
rect 40494 7692 40500 7744
rect 40552 7692 40558 7744
rect 2024 7642 77924 7664
rect 2024 7590 5794 7642
rect 5846 7590 5858 7642
rect 5910 7590 5922 7642
rect 5974 7590 5986 7642
rect 6038 7590 6050 7642
rect 6102 7590 36514 7642
rect 36566 7590 36578 7642
rect 36630 7590 36642 7642
rect 36694 7590 36706 7642
rect 36758 7590 36770 7642
rect 36822 7590 67234 7642
rect 67286 7590 67298 7642
rect 67350 7590 67362 7642
rect 67414 7590 67426 7642
rect 67478 7590 67490 7642
rect 67542 7590 77924 7642
rect 2024 7568 77924 7590
rect 10778 7488 10784 7540
rect 10836 7528 10842 7540
rect 10836 7500 15424 7528
rect 10836 7488 10842 7500
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 11112 7364 12725 7392
rect 11112 7352 11118 7364
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 14274 7352 14280 7404
rect 14332 7352 14338 7404
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 15396 7401 15424 7500
rect 16298 7488 16304 7540
rect 16356 7528 16362 7540
rect 17589 7531 17647 7537
rect 17589 7528 17601 7531
rect 16356 7500 17601 7528
rect 16356 7488 16362 7500
rect 17589 7497 17601 7500
rect 17635 7497 17647 7531
rect 17589 7491 17647 7497
rect 20349 7531 20407 7537
rect 20349 7497 20361 7531
rect 20395 7528 20407 7531
rect 22278 7528 22284 7540
rect 20395 7500 22284 7528
rect 20395 7497 20407 7500
rect 20349 7491 20407 7497
rect 22278 7488 22284 7500
rect 22336 7488 22342 7540
rect 23382 7488 23388 7540
rect 23440 7488 23446 7540
rect 27614 7528 27620 7540
rect 23492 7500 27620 7528
rect 16482 7420 16488 7472
rect 16540 7460 16546 7472
rect 19702 7460 19708 7472
rect 16540 7432 17908 7460
rect 16540 7420 16546 7432
rect 15381 7395 15439 7401
rect 14516 7364 15240 7392
rect 14516 7352 14522 7364
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7293 15163 7327
rect 15212 7324 15240 7364
rect 15381 7361 15393 7395
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 17880 7401 17908 7432
rect 18064 7432 19708 7460
rect 17773 7395 17831 7401
rect 17773 7392 17785 7395
rect 15528 7364 17785 7392
rect 15528 7352 15534 7364
rect 17773 7361 17785 7364
rect 17819 7361 17831 7395
rect 17773 7355 17831 7361
rect 17865 7395 17923 7401
rect 17865 7361 17877 7395
rect 17911 7361 17923 7395
rect 17865 7355 17923 7361
rect 16577 7327 16635 7333
rect 16577 7324 16589 7327
rect 15212 7296 16589 7324
rect 15105 7287 15163 7293
rect 16577 7293 16589 7296
rect 16623 7293 16635 7327
rect 16577 7287 16635 7293
rect 17405 7327 17463 7333
rect 17405 7293 17417 7327
rect 17451 7324 17463 7327
rect 18064 7324 18092 7432
rect 19702 7420 19708 7432
rect 19760 7420 19766 7472
rect 21818 7460 21824 7472
rect 21100 7432 21824 7460
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7392 18199 7395
rect 18969 7395 19027 7401
rect 18969 7392 18981 7395
rect 18187 7364 18981 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 18969 7361 18981 7364
rect 19015 7361 19027 7395
rect 18969 7355 19027 7361
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 20714 7392 20720 7404
rect 19659 7364 20720 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 20714 7352 20720 7364
rect 20772 7352 20778 7404
rect 21100 7401 21128 7432
rect 21818 7420 21824 7432
rect 21876 7420 21882 7472
rect 22020 7432 22876 7460
rect 21085 7395 21143 7401
rect 21085 7361 21097 7395
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 21174 7352 21180 7404
rect 21232 7352 21238 7404
rect 21270 7395 21328 7401
rect 21270 7361 21282 7395
rect 21316 7361 21328 7395
rect 21270 7355 21328 7361
rect 17451 7296 18092 7324
rect 18233 7327 18291 7333
rect 17451 7293 17463 7296
rect 17405 7287 17463 7293
rect 18233 7293 18245 7327
rect 18279 7293 18291 7327
rect 19426 7324 19432 7336
rect 18233 7287 18291 7293
rect 18708 7296 19432 7324
rect 14461 7259 14519 7265
rect 14461 7225 14473 7259
rect 14507 7256 14519 7259
rect 15120 7256 15148 7287
rect 14507 7228 15148 7256
rect 14507 7225 14519 7228
rect 14461 7219 14519 7225
rect 15194 7216 15200 7268
rect 15252 7256 15258 7268
rect 16761 7259 16819 7265
rect 16761 7256 16773 7259
rect 15252 7228 16773 7256
rect 15252 7216 15258 7228
rect 16761 7225 16773 7228
rect 16807 7225 16819 7259
rect 18248 7256 18276 7287
rect 16761 7219 16819 7225
rect 16868 7228 18276 7256
rect 12342 7148 12348 7200
rect 12400 7188 12406 7200
rect 12529 7191 12587 7197
rect 12529 7188 12541 7191
rect 12400 7160 12541 7188
rect 12400 7148 12406 7160
rect 12529 7157 12541 7160
rect 12575 7157 12587 7191
rect 12529 7151 12587 7157
rect 14550 7148 14556 7200
rect 14608 7148 14614 7200
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 15470 7188 15476 7200
rect 15068 7160 15476 7188
rect 15068 7148 15074 7160
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 15838 7148 15844 7200
rect 15896 7188 15902 7200
rect 15933 7191 15991 7197
rect 15933 7188 15945 7191
rect 15896 7160 15945 7188
rect 15896 7148 15902 7160
rect 15933 7157 15945 7160
rect 15979 7157 15991 7191
rect 15933 7151 15991 7157
rect 16022 7148 16028 7200
rect 16080 7148 16086 7200
rect 16206 7148 16212 7200
rect 16264 7188 16270 7200
rect 16868 7188 16896 7228
rect 16264 7160 16896 7188
rect 18049 7191 18107 7197
rect 16264 7148 16270 7160
rect 18049 7157 18061 7191
rect 18095 7188 18107 7191
rect 18708 7188 18736 7296
rect 19426 7284 19432 7296
rect 19484 7284 19490 7336
rect 19797 7327 19855 7333
rect 19797 7293 19809 7327
rect 19843 7324 19855 7327
rect 20441 7327 20499 7333
rect 20441 7324 20453 7327
rect 19843 7296 20453 7324
rect 19843 7293 19855 7296
rect 19797 7287 19855 7293
rect 20441 7293 20453 7296
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 20622 7284 20628 7336
rect 20680 7324 20686 7336
rect 21285 7324 21313 7355
rect 21450 7352 21456 7404
rect 21508 7352 21514 7404
rect 21542 7352 21548 7404
rect 21600 7352 21606 7404
rect 21634 7352 21640 7404
rect 21692 7401 21698 7404
rect 21692 7392 21700 7401
rect 22020 7392 22048 7432
rect 21692 7364 22048 7392
rect 21692 7355 21700 7364
rect 21692 7352 21698 7355
rect 21726 7324 21732 7336
rect 20680 7296 21732 7324
rect 20680 7284 20686 7296
rect 21726 7284 21732 7296
rect 21784 7284 21790 7336
rect 22002 7284 22008 7336
rect 22060 7284 22066 7336
rect 22554 7284 22560 7336
rect 22612 7324 22618 7336
rect 22741 7327 22799 7333
rect 22741 7324 22753 7327
rect 22612 7296 22753 7324
rect 22612 7284 22618 7296
rect 22741 7293 22753 7296
rect 22787 7293 22799 7327
rect 22848 7324 22876 7432
rect 23014 7420 23020 7472
rect 23072 7460 23078 7472
rect 23492 7460 23520 7500
rect 27614 7488 27620 7500
rect 27672 7488 27678 7540
rect 29549 7531 29607 7537
rect 29549 7497 29561 7531
rect 29595 7528 29607 7531
rect 29822 7528 29828 7540
rect 29595 7500 29828 7528
rect 29595 7497 29607 7500
rect 29549 7491 29607 7497
rect 29822 7488 29828 7500
rect 29880 7488 29886 7540
rect 30190 7488 30196 7540
rect 30248 7528 30254 7540
rect 31662 7528 31668 7540
rect 30248 7500 31668 7528
rect 30248 7488 30254 7500
rect 31662 7488 31668 7500
rect 31720 7488 31726 7540
rect 32214 7488 32220 7540
rect 32272 7488 32278 7540
rect 32858 7488 32864 7540
rect 32916 7528 32922 7540
rect 33042 7528 33048 7540
rect 32916 7500 33048 7528
rect 32916 7488 32922 7500
rect 33042 7488 33048 7500
rect 33100 7488 33106 7540
rect 33965 7531 34023 7537
rect 33965 7497 33977 7531
rect 34011 7528 34023 7531
rect 34606 7528 34612 7540
rect 34011 7500 34612 7528
rect 34011 7497 34023 7500
rect 33965 7491 34023 7497
rect 34606 7488 34612 7500
rect 34664 7488 34670 7540
rect 34701 7531 34759 7537
rect 34701 7497 34713 7531
rect 34747 7528 34759 7531
rect 36262 7528 36268 7540
rect 34747 7500 36268 7528
rect 34747 7497 34759 7500
rect 34701 7491 34759 7497
rect 36262 7488 36268 7500
rect 36320 7488 36326 7540
rect 23072 7432 23520 7460
rect 23072 7420 23078 7432
rect 24486 7420 24492 7472
rect 24544 7460 24550 7472
rect 25317 7463 25375 7469
rect 25317 7460 25329 7463
rect 24544 7432 25329 7460
rect 24544 7420 24550 7432
rect 25317 7429 25329 7432
rect 25363 7429 25375 7463
rect 25317 7423 25375 7429
rect 26786 7420 26792 7472
rect 26844 7460 26850 7472
rect 27341 7463 27399 7469
rect 27341 7460 27353 7463
rect 26844 7432 27353 7460
rect 26844 7420 26850 7432
rect 27341 7429 27353 7432
rect 27387 7429 27399 7463
rect 27341 7423 27399 7429
rect 26418 7352 26424 7404
rect 26476 7352 26482 7404
rect 26970 7352 26976 7404
rect 27028 7392 27034 7404
rect 27065 7395 27123 7401
rect 27065 7392 27077 7395
rect 27028 7364 27077 7392
rect 27028 7352 27034 7364
rect 27065 7361 27077 7364
rect 27111 7361 27123 7395
rect 27356 7392 27384 7423
rect 27430 7420 27436 7472
rect 27488 7420 27494 7472
rect 27522 7420 27528 7472
rect 27580 7420 27586 7472
rect 29638 7420 29644 7472
rect 29696 7460 29702 7472
rect 30282 7460 30288 7472
rect 29696 7432 30288 7460
rect 29696 7420 29702 7432
rect 28166 7392 28172 7404
rect 27356 7364 28172 7392
rect 27065 7355 27123 7361
rect 28166 7352 28172 7364
rect 28224 7352 28230 7404
rect 28261 7395 28319 7401
rect 28261 7361 28273 7395
rect 28307 7392 28319 7395
rect 28718 7392 28724 7404
rect 28307 7364 28724 7392
rect 28307 7361 28319 7364
rect 28261 7355 28319 7361
rect 28718 7352 28724 7364
rect 28776 7352 28782 7404
rect 29748 7401 29776 7432
rect 30282 7420 30288 7432
rect 30340 7420 30346 7472
rect 31386 7420 31392 7472
rect 31444 7460 31450 7472
rect 32125 7463 32183 7469
rect 32125 7460 32137 7463
rect 31444 7432 32137 7460
rect 31444 7420 31450 7432
rect 32125 7429 32137 7432
rect 32171 7460 32183 7463
rect 32171 7432 32812 7460
rect 32171 7429 32183 7432
rect 32125 7423 32183 7429
rect 29733 7395 29791 7401
rect 29733 7361 29745 7395
rect 29779 7361 29791 7395
rect 29733 7355 29791 7361
rect 31110 7352 31116 7404
rect 31168 7352 31174 7404
rect 31662 7352 31668 7404
rect 31720 7392 31726 7404
rect 31849 7395 31907 7401
rect 31849 7392 31861 7395
rect 31720 7364 31861 7392
rect 31720 7352 31726 7364
rect 31849 7361 31861 7364
rect 31895 7361 31907 7395
rect 31849 7355 31907 7361
rect 31941 7395 31999 7401
rect 31941 7361 31953 7395
rect 31987 7392 31999 7395
rect 32306 7392 32312 7404
rect 31987 7364 32312 7392
rect 31987 7361 31999 7364
rect 31941 7355 31999 7361
rect 32306 7352 32312 7364
rect 32364 7352 32370 7404
rect 32490 7352 32496 7404
rect 32548 7352 32554 7404
rect 32784 7392 32812 7432
rect 33134 7420 33140 7472
rect 33192 7460 33198 7472
rect 33192 7432 34560 7460
rect 33192 7420 33198 7432
rect 33226 7392 33232 7404
rect 32784 7364 33232 7392
rect 33226 7352 33232 7364
rect 33284 7392 33290 7404
rect 33321 7395 33379 7401
rect 33321 7392 33333 7395
rect 33284 7364 33333 7392
rect 33284 7352 33290 7364
rect 33321 7361 33333 7364
rect 33367 7361 33379 7395
rect 33321 7355 33379 7361
rect 33502 7352 33508 7404
rect 33560 7392 33566 7404
rect 34054 7392 34060 7404
rect 33560 7364 34060 7392
rect 33560 7352 33566 7364
rect 34054 7352 34060 7364
rect 34112 7352 34118 7404
rect 34532 7401 34560 7432
rect 34517 7395 34575 7401
rect 34517 7361 34529 7395
rect 34563 7361 34575 7395
rect 34517 7355 34575 7361
rect 35710 7352 35716 7404
rect 35768 7392 35774 7404
rect 37093 7395 37151 7401
rect 37093 7392 37105 7395
rect 35768 7364 37105 7392
rect 35768 7352 35774 7364
rect 37093 7361 37105 7364
rect 37139 7361 37151 7395
rect 37093 7355 37151 7361
rect 37458 7352 37464 7404
rect 37516 7352 37522 7404
rect 38562 7352 38568 7404
rect 38620 7392 38626 7404
rect 40589 7395 40647 7401
rect 40589 7392 40601 7395
rect 38620 7364 40601 7392
rect 38620 7352 38626 7364
rect 40589 7361 40601 7364
rect 40635 7361 40647 7395
rect 40589 7355 40647 7361
rect 41414 7352 41420 7404
rect 41472 7352 41478 7404
rect 23658 7324 23664 7336
rect 22848 7296 23664 7324
rect 22741 7287 22799 7293
rect 23658 7284 23664 7296
rect 23716 7284 23722 7336
rect 23753 7327 23811 7333
rect 23753 7293 23765 7327
rect 23799 7324 23811 7327
rect 23934 7324 23940 7336
rect 23799 7296 23940 7324
rect 23799 7293 23811 7296
rect 23753 7287 23811 7293
rect 23934 7284 23940 7296
rect 23992 7284 23998 7336
rect 24121 7327 24179 7333
rect 24121 7293 24133 7327
rect 24167 7324 24179 7327
rect 24394 7324 24400 7336
rect 24167 7296 24400 7324
rect 24167 7293 24179 7296
rect 24121 7287 24179 7293
rect 24394 7284 24400 7296
rect 24452 7284 24458 7336
rect 24946 7284 24952 7336
rect 25004 7284 25010 7336
rect 25038 7284 25044 7336
rect 25096 7284 25102 7336
rect 28905 7327 28963 7333
rect 28905 7324 28917 7327
rect 28736 7296 28917 7324
rect 18877 7259 18935 7265
rect 18877 7225 18889 7259
rect 18923 7256 18935 7259
rect 23198 7256 23204 7268
rect 18923 7228 23204 7256
rect 18923 7225 18935 7228
rect 18877 7219 18935 7225
rect 23198 7216 23204 7228
rect 23256 7216 23262 7268
rect 24762 7256 24768 7268
rect 23308 7228 24768 7256
rect 18095 7160 18736 7188
rect 18095 7157 18107 7160
rect 18049 7151 18107 7157
rect 18782 7148 18788 7200
rect 18840 7188 18846 7200
rect 20714 7188 20720 7200
rect 18840 7160 20720 7188
rect 18840 7148 18846 7160
rect 20714 7148 20720 7160
rect 20772 7148 20778 7200
rect 21818 7148 21824 7200
rect 21876 7148 21882 7200
rect 22002 7148 22008 7200
rect 22060 7188 22066 7200
rect 22186 7188 22192 7200
rect 22060 7160 22192 7188
rect 22060 7148 22066 7160
rect 22186 7148 22192 7160
rect 22244 7148 22250 7200
rect 22554 7148 22560 7200
rect 22612 7148 22618 7200
rect 22830 7148 22836 7200
rect 22888 7188 22894 7200
rect 23308 7188 23336 7228
rect 24762 7216 24768 7228
rect 24820 7216 24826 7268
rect 27154 7216 27160 7268
rect 27212 7216 27218 7268
rect 28534 7256 28540 7268
rect 27264 7228 28540 7256
rect 22888 7160 23336 7188
rect 22888 7148 22894 7160
rect 23474 7148 23480 7200
rect 23532 7148 23538 7200
rect 23658 7148 23664 7200
rect 23716 7188 23722 7200
rect 24305 7191 24363 7197
rect 24305 7188 24317 7191
rect 23716 7160 24317 7188
rect 23716 7148 23722 7160
rect 24305 7157 24317 7160
rect 24351 7157 24363 7191
rect 24305 7151 24363 7157
rect 25866 7148 25872 7200
rect 25924 7188 25930 7200
rect 27264 7188 27292 7228
rect 28534 7216 28540 7228
rect 28592 7216 28598 7268
rect 25924 7160 27292 7188
rect 27709 7191 27767 7197
rect 25924 7148 25930 7160
rect 27709 7157 27721 7191
rect 27755 7188 27767 7191
rect 27798 7188 27804 7200
rect 27755 7160 27804 7188
rect 27755 7157 27767 7160
rect 27709 7151 27767 7157
rect 27798 7148 27804 7160
rect 27856 7148 27862 7200
rect 28736 7188 28764 7296
rect 28905 7293 28917 7296
rect 28951 7293 28963 7327
rect 30009 7327 30067 7333
rect 30009 7324 30021 7327
rect 28905 7287 28963 7293
rect 29472 7296 30021 7324
rect 28813 7259 28871 7265
rect 28813 7225 28825 7259
rect 28859 7256 28871 7259
rect 29472 7256 29500 7296
rect 30009 7293 30021 7296
rect 30055 7293 30067 7327
rect 31128 7324 31156 7352
rect 30009 7287 30067 7293
rect 31036 7296 31156 7324
rect 31757 7327 31815 7333
rect 28859 7228 29500 7256
rect 28859 7225 28871 7228
rect 28813 7219 28871 7225
rect 30190 7188 30196 7200
rect 28736 7160 30196 7188
rect 30190 7148 30196 7160
rect 30248 7148 30254 7200
rect 31036 7188 31064 7296
rect 31757 7293 31769 7327
rect 31803 7293 31815 7327
rect 31757 7287 31815 7293
rect 32052 7327 32110 7333
rect 32052 7293 32064 7327
rect 32098 7324 32110 7327
rect 32401 7327 32459 7333
rect 32401 7324 32413 7327
rect 32098 7296 32413 7324
rect 32098 7293 32110 7296
rect 32052 7287 32110 7293
rect 32401 7293 32413 7296
rect 32447 7293 32459 7327
rect 32401 7287 32459 7293
rect 32769 7327 32827 7333
rect 32769 7293 32781 7327
rect 32815 7293 32827 7327
rect 32769 7287 32827 7293
rect 31772 7256 31800 7287
rect 32214 7256 32220 7268
rect 31772 7228 32220 7256
rect 32214 7216 32220 7228
rect 32272 7216 32278 7268
rect 32398 7188 32404 7200
rect 31036 7160 32404 7188
rect 32398 7148 32404 7160
rect 32456 7148 32462 7200
rect 32784 7188 32812 7287
rect 32858 7284 32864 7336
rect 32916 7284 32922 7336
rect 34330 7284 34336 7336
rect 34388 7284 34394 7336
rect 34422 7284 34428 7336
rect 34480 7324 34486 7336
rect 34793 7327 34851 7333
rect 34793 7324 34805 7327
rect 34480 7296 34805 7324
rect 34480 7284 34486 7296
rect 34793 7293 34805 7296
rect 34839 7293 34851 7327
rect 34793 7287 34851 7293
rect 36449 7327 36507 7333
rect 36449 7293 36461 7327
rect 36495 7324 36507 7327
rect 36541 7327 36599 7333
rect 36541 7324 36553 7327
rect 36495 7296 36553 7324
rect 36495 7293 36507 7296
rect 36449 7287 36507 7293
rect 36541 7293 36553 7296
rect 36587 7293 36599 7327
rect 36541 7287 36599 7293
rect 38013 7327 38071 7333
rect 38013 7293 38025 7327
rect 38059 7324 38071 7327
rect 38749 7327 38807 7333
rect 38749 7324 38761 7327
rect 38059 7296 38761 7324
rect 38059 7293 38071 7296
rect 38013 7287 38071 7293
rect 38749 7293 38761 7296
rect 38795 7293 38807 7327
rect 38749 7287 38807 7293
rect 39761 7327 39819 7333
rect 39761 7293 39773 7327
rect 39807 7324 39819 7327
rect 40037 7327 40095 7333
rect 40037 7324 40049 7327
rect 39807 7296 40049 7324
rect 39807 7293 39819 7296
rect 39761 7287 39819 7293
rect 40037 7293 40049 7296
rect 40083 7293 40095 7327
rect 40037 7287 40095 7293
rect 35526 7216 35532 7268
rect 35584 7256 35590 7268
rect 35805 7259 35863 7265
rect 35805 7256 35817 7259
rect 35584 7228 35817 7256
rect 35584 7216 35590 7228
rect 35805 7225 35817 7228
rect 35851 7225 35863 7259
rect 35805 7219 35863 7225
rect 37458 7216 37464 7268
rect 37516 7256 37522 7268
rect 39117 7259 39175 7265
rect 39117 7256 39129 7259
rect 37516 7228 39129 7256
rect 37516 7216 37522 7228
rect 39117 7225 39129 7228
rect 39163 7225 39175 7259
rect 39117 7219 39175 7225
rect 34238 7188 34244 7200
rect 32784 7160 34244 7188
rect 34238 7148 34244 7160
rect 34296 7148 34302 7200
rect 35437 7191 35495 7197
rect 35437 7157 35449 7191
rect 35483 7188 35495 7191
rect 35710 7188 35716 7200
rect 35483 7160 35716 7188
rect 35483 7157 35495 7160
rect 35437 7151 35495 7157
rect 35710 7148 35716 7160
rect 35768 7148 35774 7200
rect 37274 7148 37280 7200
rect 37332 7188 37338 7200
rect 38197 7191 38255 7197
rect 38197 7188 38209 7191
rect 37332 7160 38209 7188
rect 37332 7148 37338 7160
rect 38197 7157 38209 7160
rect 38243 7157 38255 7191
rect 38197 7151 38255 7157
rect 40678 7148 40684 7200
rect 40736 7188 40742 7200
rect 40773 7191 40831 7197
rect 40773 7188 40785 7191
rect 40736 7160 40785 7188
rect 40736 7148 40742 7160
rect 40773 7157 40785 7160
rect 40819 7157 40831 7191
rect 40773 7151 40831 7157
rect 2024 7098 77924 7120
rect 2024 7046 5134 7098
rect 5186 7046 5198 7098
rect 5250 7046 5262 7098
rect 5314 7046 5326 7098
rect 5378 7046 5390 7098
rect 5442 7046 35854 7098
rect 35906 7046 35918 7098
rect 35970 7046 35982 7098
rect 36034 7046 36046 7098
rect 36098 7046 36110 7098
rect 36162 7046 66574 7098
rect 66626 7046 66638 7098
rect 66690 7046 66702 7098
rect 66754 7046 66766 7098
rect 66818 7046 66830 7098
rect 66882 7046 77924 7098
rect 2024 7024 77924 7046
rect 14274 6984 14280 6996
rect 6886 6956 14280 6984
rect 4522 6876 4528 6928
rect 4580 6916 4586 6928
rect 6886 6916 6914 6956
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 15838 6944 15844 6996
rect 15896 6984 15902 6996
rect 18782 6984 18788 6996
rect 15896 6956 18788 6984
rect 15896 6944 15902 6956
rect 18782 6944 18788 6956
rect 18840 6944 18846 6996
rect 19886 6984 19892 6996
rect 19168 6956 19892 6984
rect 4580 6888 6914 6916
rect 4580 6876 4586 6888
rect 10962 6876 10968 6928
rect 11020 6916 11026 6928
rect 11020 6888 12664 6916
rect 11020 6876 11026 6888
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 4396 6820 12541 6848
rect 4396 6808 4402 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12636 6848 12664 6888
rect 14642 6876 14648 6928
rect 14700 6916 14706 6928
rect 16482 6916 16488 6928
rect 14700 6888 16488 6916
rect 14700 6876 14706 6888
rect 16482 6876 16488 6888
rect 16540 6876 16546 6928
rect 19168 6916 19196 6956
rect 19886 6944 19892 6956
rect 19944 6984 19950 6996
rect 20428 6987 20486 6993
rect 19944 6956 20300 6984
rect 19944 6944 19950 6956
rect 17696 6888 19196 6916
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 12636 6820 13277 6848
rect 12529 6811 12587 6817
rect 13265 6817 13277 6820
rect 13311 6817 13323 6851
rect 15565 6851 15623 6857
rect 13265 6811 13323 6817
rect 13832 6820 15516 6848
rect 10594 6740 10600 6792
rect 10652 6740 10658 6792
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 11149 6783 11207 6789
rect 10744 6752 11100 6780
rect 10744 6740 10750 6752
rect 11072 6712 11100 6752
rect 11149 6749 11161 6783
rect 11195 6780 11207 6783
rect 11606 6780 11612 6792
rect 11195 6752 11612 6780
rect 11195 6749 11207 6752
rect 11149 6743 11207 6749
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 11790 6740 11796 6792
rect 11848 6740 11854 6792
rect 12434 6740 12440 6792
rect 12492 6740 12498 6792
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 11241 6715 11299 6721
rect 11241 6712 11253 6715
rect 11072 6684 11253 6712
rect 11241 6681 11253 6684
rect 11287 6681 11299 6715
rect 11241 6675 11299 6681
rect 11330 6672 11336 6724
rect 11388 6712 11394 6724
rect 13096 6712 13124 6743
rect 11388 6684 13124 6712
rect 11388 6672 11394 6684
rect 8386 6604 8392 6656
rect 8444 6644 8450 6656
rect 12253 6647 12311 6653
rect 12253 6644 12265 6647
rect 8444 6616 12265 6644
rect 8444 6604 8450 6616
rect 12253 6613 12265 6616
rect 12299 6613 12311 6647
rect 12253 6607 12311 6613
rect 12526 6604 12532 6656
rect 12584 6644 12590 6656
rect 13832 6644 13860 6820
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6780 14887 6783
rect 14918 6780 14924 6792
rect 14875 6752 14924 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 15488 6780 15516 6820
rect 15565 6817 15577 6851
rect 15611 6848 15623 6851
rect 16298 6848 16304 6860
rect 15611 6820 16304 6848
rect 15611 6817 15623 6820
rect 15565 6811 15623 6817
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 17696 6848 17724 6888
rect 16408 6820 17724 6848
rect 15488 6752 15608 6780
rect 13909 6715 13967 6721
rect 13909 6681 13921 6715
rect 13955 6712 13967 6715
rect 15470 6712 15476 6724
rect 13955 6684 15476 6712
rect 13955 6681 13967 6684
rect 13909 6675 13967 6681
rect 15470 6672 15476 6684
rect 15528 6672 15534 6724
rect 15580 6712 15608 6752
rect 15654 6740 15660 6792
rect 15712 6740 15718 6792
rect 16408 6780 16436 6820
rect 17770 6808 17776 6860
rect 17828 6808 17834 6860
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 20272 6848 20300 6956
rect 20428 6953 20440 6987
rect 20474 6984 20486 6987
rect 20530 6984 20536 6996
rect 20474 6956 20536 6984
rect 20474 6953 20486 6956
rect 20428 6947 20486 6953
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 22465 6987 22523 6993
rect 22465 6984 22477 6987
rect 21468 6956 22477 6984
rect 21468 6848 21496 6956
rect 22465 6953 22477 6956
rect 22511 6953 22523 6987
rect 22465 6947 22523 6953
rect 22738 6944 22744 6996
rect 22796 6984 22802 6996
rect 23382 6984 23388 6996
rect 22796 6956 23388 6984
rect 22796 6944 22802 6956
rect 23382 6944 23388 6956
rect 23440 6944 23446 6996
rect 24121 6987 24179 6993
rect 23584 6956 23888 6984
rect 21818 6876 21824 6928
rect 21876 6916 21882 6928
rect 21876 6888 22508 6916
rect 21876 6876 21882 6888
rect 22370 6848 22376 6860
rect 18104 6820 20208 6848
rect 20272 6820 21496 6848
rect 22296 6820 22376 6848
rect 18104 6808 18110 6820
rect 20180 6792 20208 6820
rect 16224 6752 16436 6780
rect 16224 6712 16252 6752
rect 16482 6740 16488 6792
rect 16540 6740 16546 6792
rect 17037 6783 17095 6789
rect 17037 6749 17049 6783
rect 17083 6780 17095 6783
rect 17862 6780 17868 6792
rect 17083 6752 17868 6780
rect 17083 6749 17095 6752
rect 17037 6743 17095 6749
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 17957 6783 18015 6789
rect 17957 6749 17969 6783
rect 18003 6749 18015 6783
rect 17957 6743 18015 6749
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6780 18751 6783
rect 19058 6780 19064 6792
rect 18739 6752 19064 6780
rect 18739 6749 18751 6752
rect 18693 6743 18751 6749
rect 15580 6684 16252 6712
rect 16301 6715 16359 6721
rect 16301 6681 16313 6715
rect 16347 6712 16359 6715
rect 17972 6712 18000 6743
rect 19058 6740 19064 6752
rect 19116 6740 19122 6792
rect 19245 6783 19303 6789
rect 19245 6749 19257 6783
rect 19291 6780 19303 6783
rect 19334 6780 19340 6792
rect 19291 6752 19340 6780
rect 19291 6749 19303 6752
rect 19245 6743 19303 6749
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 19610 6740 19616 6792
rect 19668 6780 19674 6792
rect 19889 6783 19947 6789
rect 19889 6780 19901 6783
rect 19668 6752 19901 6780
rect 19668 6740 19674 6752
rect 19889 6749 19901 6752
rect 19935 6749 19947 6783
rect 19889 6743 19947 6749
rect 20162 6740 20168 6792
rect 20220 6740 20226 6792
rect 22186 6740 22192 6792
rect 22244 6740 22250 6792
rect 20530 6712 20536 6724
rect 16347 6684 17908 6712
rect 17972 6684 20536 6712
rect 16347 6681 16359 6684
rect 16301 6675 16359 6681
rect 12584 6616 13860 6644
rect 12584 6604 12590 6616
rect 14274 6604 14280 6656
rect 14332 6604 14338 6656
rect 14366 6604 14372 6656
rect 14424 6644 14430 6656
rect 15105 6647 15163 6653
rect 15105 6644 15117 6647
rect 14424 6616 15117 6644
rect 14424 6604 14430 6616
rect 15105 6613 15117 6616
rect 15151 6613 15163 6647
rect 15105 6607 15163 6613
rect 17129 6647 17187 6653
rect 17129 6613 17141 6647
rect 17175 6644 17187 6647
rect 17218 6644 17224 6656
rect 17175 6616 17224 6644
rect 17175 6613 17187 6616
rect 17129 6607 17187 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 17880 6644 17908 6684
rect 20530 6672 20536 6684
rect 20588 6672 20594 6724
rect 22094 6712 22100 6724
rect 21666 6684 22100 6712
rect 22094 6672 22100 6684
rect 22152 6672 22158 6724
rect 22296 6721 22324 6820
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 22281 6715 22339 6721
rect 22281 6681 22293 6715
rect 22327 6681 22339 6715
rect 22480 6712 22508 6888
rect 22646 6876 22652 6928
rect 22704 6916 22710 6928
rect 23584 6916 23612 6956
rect 22704 6888 23612 6916
rect 22704 6876 22710 6888
rect 22833 6851 22891 6857
rect 22833 6817 22845 6851
rect 22879 6848 22891 6851
rect 22922 6848 22928 6860
rect 22879 6820 22928 6848
rect 22879 6817 22891 6820
rect 22833 6811 22891 6817
rect 22922 6808 22928 6820
rect 22980 6808 22986 6860
rect 23290 6808 23296 6860
rect 23348 6848 23354 6860
rect 23385 6851 23443 6857
rect 23385 6848 23397 6851
rect 23348 6820 23397 6848
rect 23348 6808 23354 6820
rect 23385 6817 23397 6820
rect 23431 6817 23443 6851
rect 23385 6811 23443 6817
rect 23474 6808 23480 6860
rect 23532 6808 23538 6860
rect 23860 6848 23888 6956
rect 24121 6953 24133 6987
rect 24167 6984 24179 6987
rect 24486 6984 24492 6996
rect 24167 6956 24492 6984
rect 24167 6953 24179 6956
rect 24121 6947 24179 6953
rect 24486 6944 24492 6956
rect 24544 6944 24550 6996
rect 25866 6944 25872 6996
rect 25924 6944 25930 6996
rect 27430 6944 27436 6996
rect 27488 6984 27494 6996
rect 30558 6984 30564 6996
rect 27488 6956 30564 6984
rect 27488 6944 27494 6956
rect 30558 6944 30564 6956
rect 30616 6944 30622 6996
rect 31018 6944 31024 6996
rect 31076 6944 31082 6996
rect 32493 6987 32551 6993
rect 32493 6953 32505 6987
rect 32539 6984 32551 6987
rect 32858 6984 32864 6996
rect 32539 6956 32864 6984
rect 32539 6953 32551 6956
rect 32493 6947 32551 6953
rect 32858 6944 32864 6956
rect 32916 6944 32922 6996
rect 34701 6987 34759 6993
rect 34701 6953 34713 6987
rect 34747 6984 34759 6987
rect 35158 6984 35164 6996
rect 34747 6956 35164 6984
rect 34747 6953 34759 6956
rect 34701 6947 34759 6953
rect 35158 6944 35164 6956
rect 35216 6944 35222 6996
rect 35897 6987 35955 6993
rect 35897 6953 35909 6987
rect 35943 6984 35955 6987
rect 36354 6984 36360 6996
rect 35943 6956 36360 6984
rect 35943 6953 35955 6956
rect 35897 6947 35955 6953
rect 36354 6944 36360 6956
rect 36412 6944 36418 6996
rect 24026 6876 24032 6928
rect 24084 6916 24090 6928
rect 25038 6916 25044 6928
rect 24084 6888 25044 6916
rect 24084 6876 24090 6888
rect 25038 6876 25044 6888
rect 25096 6916 25102 6928
rect 25096 6888 26740 6916
rect 25096 6876 25102 6888
rect 24118 6848 24124 6860
rect 23860 6820 24124 6848
rect 24118 6808 24124 6820
rect 24176 6808 24182 6860
rect 24486 6808 24492 6860
rect 24544 6848 24550 6860
rect 26712 6857 26740 6888
rect 28166 6876 28172 6928
rect 28224 6916 28230 6928
rect 28224 6888 30420 6916
rect 28224 6876 28230 6888
rect 24857 6851 24915 6857
rect 24857 6848 24869 6851
rect 24544 6820 24869 6848
rect 24544 6808 24550 6820
rect 24857 6817 24869 6820
rect 24903 6817 24915 6851
rect 24857 6811 24915 6817
rect 26697 6851 26755 6857
rect 26697 6817 26709 6851
rect 26743 6817 26755 6851
rect 26697 6811 26755 6817
rect 26970 6808 26976 6860
rect 27028 6848 27034 6860
rect 28442 6848 28448 6860
rect 27028 6820 28448 6848
rect 27028 6808 27034 6820
rect 28442 6808 28448 6820
rect 28500 6808 28506 6860
rect 28626 6808 28632 6860
rect 28684 6848 28690 6860
rect 28721 6851 28779 6857
rect 28721 6848 28733 6851
rect 28684 6820 28733 6848
rect 28684 6808 28690 6820
rect 28721 6817 28733 6820
rect 28767 6817 28779 6851
rect 28721 6811 28779 6817
rect 29549 6851 29607 6857
rect 29549 6817 29561 6851
rect 29595 6848 29607 6851
rect 29914 6848 29920 6860
rect 29595 6820 29920 6848
rect 29595 6817 29607 6820
rect 29549 6811 29607 6817
rect 29914 6808 29920 6820
rect 29972 6808 29978 6860
rect 30098 6808 30104 6860
rect 30156 6848 30162 6860
rect 30193 6851 30251 6857
rect 30193 6848 30205 6851
rect 30156 6820 30205 6848
rect 30156 6808 30162 6820
rect 30193 6817 30205 6820
rect 30239 6817 30251 6851
rect 30193 6811 30251 6817
rect 22554 6740 22560 6792
rect 22612 6780 22618 6792
rect 23566 6780 23572 6792
rect 22612 6752 23572 6780
rect 22612 6740 22618 6752
rect 23566 6740 23572 6752
rect 23624 6740 23630 6792
rect 23750 6740 23756 6792
rect 23808 6780 23814 6792
rect 23934 6780 23940 6792
rect 23808 6752 23940 6780
rect 23808 6740 23814 6752
rect 23934 6740 23940 6752
rect 23992 6740 23998 6792
rect 24213 6783 24271 6789
rect 24213 6749 24225 6783
rect 24259 6749 24271 6783
rect 24213 6743 24271 6749
rect 25317 6783 25375 6789
rect 25317 6749 25329 6783
rect 25363 6749 25375 6783
rect 25317 6743 25375 6749
rect 24228 6712 24256 6743
rect 22480 6684 24256 6712
rect 22281 6675 22339 6681
rect 18138 6644 18144 6656
rect 17880 6616 18144 6644
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 18506 6604 18512 6656
rect 18564 6604 18570 6656
rect 19334 6604 19340 6656
rect 19392 6604 19398 6656
rect 22491 6647 22549 6653
rect 22491 6613 22503 6647
rect 22537 6644 22549 6647
rect 23106 6644 23112 6656
rect 22537 6616 23112 6644
rect 22537 6613 22549 6616
rect 22491 6607 22549 6613
rect 23106 6604 23112 6616
rect 23164 6604 23170 6656
rect 23934 6604 23940 6656
rect 23992 6644 23998 6656
rect 25332 6644 25360 6743
rect 25498 6740 25504 6792
rect 25556 6740 25562 6792
rect 25685 6783 25743 6789
rect 25685 6749 25697 6783
rect 25731 6780 25743 6783
rect 25866 6780 25872 6792
rect 25731 6752 25872 6780
rect 25731 6749 25743 6752
rect 25685 6743 25743 6749
rect 25866 6740 25872 6752
rect 25924 6740 25930 6792
rect 26050 6740 26056 6792
rect 26108 6740 26114 6792
rect 28258 6780 28264 6792
rect 28106 6752 28264 6780
rect 28258 6740 28264 6752
rect 28316 6780 28322 6792
rect 28534 6780 28540 6792
rect 28316 6752 28540 6780
rect 28316 6740 28322 6752
rect 28534 6740 28540 6752
rect 28592 6740 28598 6792
rect 30392 6780 30420 6888
rect 30576 6857 30604 6944
rect 31386 6916 31392 6928
rect 30760 6888 31392 6916
rect 30561 6851 30619 6857
rect 30561 6817 30573 6851
rect 30607 6817 30619 6851
rect 30561 6811 30619 6817
rect 30650 6808 30656 6860
rect 30708 6808 30714 6860
rect 30760 6789 30788 6888
rect 31386 6876 31392 6888
rect 31444 6876 31450 6928
rect 31754 6876 31760 6928
rect 31812 6916 31818 6928
rect 34606 6916 34612 6928
rect 31812 6888 34612 6916
rect 31812 6876 31818 6888
rect 30837 6851 30895 6857
rect 30837 6817 30849 6851
rect 30883 6848 30895 6851
rect 31662 6848 31668 6860
rect 30883 6820 31668 6848
rect 30883 6817 30895 6820
rect 30837 6811 30895 6817
rect 31662 6808 31668 6820
rect 31720 6808 31726 6860
rect 33226 6848 33232 6860
rect 31772 6820 33232 6848
rect 30745 6783 30803 6789
rect 30745 6780 30757 6783
rect 30392 6752 30757 6780
rect 30745 6749 30757 6752
rect 30791 6749 30803 6783
rect 30745 6743 30803 6749
rect 31110 6740 31116 6792
rect 31168 6740 31174 6792
rect 31772 6789 31800 6820
rect 33226 6808 33232 6820
rect 33284 6808 33290 6860
rect 33336 6857 33364 6888
rect 34606 6876 34612 6888
rect 34664 6876 34670 6928
rect 35250 6876 35256 6928
rect 35308 6876 35314 6928
rect 35434 6876 35440 6928
rect 35492 6876 35498 6928
rect 35728 6888 35940 6916
rect 33321 6851 33379 6857
rect 33321 6817 33333 6851
rect 33367 6817 33379 6851
rect 33321 6811 33379 6817
rect 33965 6851 34023 6857
rect 33965 6817 33977 6851
rect 34011 6848 34023 6851
rect 34422 6848 34428 6860
rect 34011 6820 34428 6848
rect 34011 6817 34023 6820
rect 33965 6811 34023 6817
rect 34422 6808 34428 6820
rect 34480 6808 34486 6860
rect 34698 6808 34704 6860
rect 34756 6848 34762 6860
rect 35268 6848 35296 6876
rect 35728 6848 35756 6888
rect 34756 6820 35020 6848
rect 35268 6820 35756 6848
rect 35912 6848 35940 6888
rect 36449 6851 36507 6857
rect 36449 6848 36461 6851
rect 35912 6820 36461 6848
rect 34756 6808 34762 6820
rect 31757 6783 31815 6789
rect 31757 6749 31769 6783
rect 31803 6749 31815 6783
rect 31757 6743 31815 6749
rect 31846 6740 31852 6792
rect 31904 6740 31910 6792
rect 31938 6740 31944 6792
rect 31996 6780 32002 6792
rect 31996 6752 32720 6780
rect 31996 6740 32002 6752
rect 25593 6715 25651 6721
rect 25593 6681 25605 6715
rect 25639 6712 25651 6715
rect 26326 6712 26332 6724
rect 25639 6684 26332 6712
rect 25639 6681 25651 6684
rect 25593 6675 25651 6681
rect 26326 6672 26332 6684
rect 26384 6672 26390 6724
rect 26605 6715 26663 6721
rect 26605 6681 26617 6715
rect 26651 6712 26663 6715
rect 26973 6715 27031 6721
rect 26973 6712 26985 6715
rect 26651 6684 26985 6712
rect 26651 6681 26663 6684
rect 26605 6675 26663 6681
rect 26973 6681 26985 6684
rect 27019 6681 27031 6715
rect 26973 6675 27031 6681
rect 30466 6672 30472 6724
rect 30524 6712 30530 6724
rect 32585 6715 32643 6721
rect 32585 6712 32597 6715
rect 30524 6684 32597 6712
rect 30524 6672 30530 6684
rect 32585 6681 32597 6684
rect 32631 6681 32643 6715
rect 32692 6712 32720 6752
rect 33134 6740 33140 6792
rect 33192 6740 33198 6792
rect 33502 6740 33508 6792
rect 33560 6780 33566 6792
rect 34057 6783 34115 6789
rect 34057 6780 34069 6783
rect 33560 6752 34069 6780
rect 33560 6740 33566 6752
rect 34057 6749 34069 6752
rect 34103 6749 34115 6783
rect 34793 6783 34851 6789
rect 34793 6780 34805 6783
rect 34057 6743 34115 6749
rect 34164 6752 34805 6780
rect 34164 6712 34192 6752
rect 34793 6749 34805 6752
rect 34839 6749 34851 6783
rect 34793 6743 34851 6749
rect 34882 6740 34888 6792
rect 34940 6740 34946 6792
rect 34992 6780 35020 6820
rect 36449 6817 36461 6820
rect 36495 6817 36507 6851
rect 36449 6811 36507 6817
rect 37369 6851 37427 6857
rect 37369 6817 37381 6851
rect 37415 6848 37427 6851
rect 38194 6848 38200 6860
rect 37415 6820 38200 6848
rect 37415 6817 37427 6820
rect 37369 6811 37427 6817
rect 38194 6808 38200 6820
rect 38252 6808 38258 6860
rect 39390 6808 39396 6860
rect 39448 6848 39454 6860
rect 40037 6851 40095 6857
rect 40037 6848 40049 6851
rect 39448 6820 40049 6848
rect 39448 6808 39454 6820
rect 40037 6817 40049 6820
rect 40083 6817 40095 6851
rect 40037 6811 40095 6817
rect 40218 6808 40224 6860
rect 40276 6848 40282 6860
rect 40773 6851 40831 6857
rect 40773 6848 40785 6851
rect 40276 6820 40785 6848
rect 40276 6808 40282 6820
rect 40773 6817 40785 6820
rect 40819 6817 40831 6851
rect 42797 6851 42855 6857
rect 42797 6848 42809 6851
rect 40773 6811 40831 6817
rect 41386 6820 42809 6848
rect 35158 6780 35164 6792
rect 34992 6752 35164 6780
rect 35158 6740 35164 6752
rect 35216 6740 35222 6792
rect 35253 6761 35311 6767
rect 35253 6727 35265 6761
rect 35299 6758 35311 6761
rect 35299 6730 35388 6758
rect 35802 6740 35808 6792
rect 35860 6740 35866 6792
rect 36633 6783 36691 6789
rect 36633 6749 36645 6783
rect 36679 6749 36691 6783
rect 41386 6780 41414 6820
rect 42797 6817 42809 6820
rect 42843 6817 42855 6851
rect 42797 6811 42855 6817
rect 36633 6743 36691 6749
rect 38948 6752 41414 6780
rect 42153 6783 42211 6789
rect 35299 6727 35311 6730
rect 32692 6684 34192 6712
rect 32585 6675 32643 6681
rect 34238 6672 34244 6724
rect 34296 6712 34302 6724
rect 34422 6712 34428 6724
rect 34296 6684 34428 6712
rect 34296 6672 34302 6684
rect 34422 6672 34428 6684
rect 34480 6672 34486 6724
rect 34606 6672 34612 6724
rect 34664 6712 34670 6724
rect 35253 6721 35311 6727
rect 35069 6715 35127 6721
rect 35069 6712 35081 6715
rect 34664 6684 35081 6712
rect 34664 6672 34670 6684
rect 35069 6681 35081 6684
rect 35115 6681 35127 6715
rect 35069 6675 35127 6681
rect 23992 6616 25360 6644
rect 23992 6604 23998 6616
rect 28258 6604 28264 6656
rect 28316 6644 28322 6656
rect 28905 6647 28963 6653
rect 28905 6644 28917 6647
rect 28316 6616 28917 6644
rect 28316 6604 28322 6616
rect 28905 6613 28917 6616
rect 28951 6613 28963 6647
rect 28905 6607 28963 6613
rect 28994 6604 29000 6656
rect 29052 6644 29058 6656
rect 29641 6647 29699 6653
rect 29641 6644 29653 6647
rect 29052 6616 29653 6644
rect 29052 6604 29058 6616
rect 29641 6613 29653 6616
rect 29687 6613 29699 6647
rect 29641 6607 29699 6613
rect 29914 6604 29920 6656
rect 29972 6644 29978 6656
rect 31202 6644 31208 6656
rect 29972 6616 31208 6644
rect 29972 6604 29978 6616
rect 31202 6604 31208 6616
rect 31260 6604 31266 6656
rect 31938 6604 31944 6656
rect 31996 6644 32002 6656
rect 33502 6644 33508 6656
rect 31996 6616 33508 6644
rect 31996 6604 32002 6616
rect 33502 6604 33508 6616
rect 33560 6604 33566 6656
rect 34054 6604 34060 6656
rect 34112 6644 34118 6656
rect 35158 6644 35164 6656
rect 34112 6616 35164 6644
rect 34112 6604 34118 6616
rect 35158 6604 35164 6616
rect 35216 6644 35222 6656
rect 35360 6644 35388 6730
rect 35986 6672 35992 6724
rect 36044 6712 36050 6724
rect 36044 6684 36308 6712
rect 36044 6672 36050 6684
rect 35216 6616 35388 6644
rect 35713 6647 35771 6653
rect 35216 6604 35222 6616
rect 35713 6613 35725 6647
rect 35759 6644 35771 6647
rect 35894 6644 35900 6656
rect 35759 6616 35900 6644
rect 35759 6613 35771 6616
rect 35713 6607 35771 6613
rect 35894 6604 35900 6616
rect 35952 6604 35958 6656
rect 36280 6644 36308 6684
rect 36354 6672 36360 6724
rect 36412 6712 36418 6724
rect 36648 6712 36676 6743
rect 36412 6684 36676 6712
rect 37277 6715 37335 6721
rect 36412 6672 36418 6684
rect 37277 6681 37289 6715
rect 37323 6712 37335 6715
rect 37645 6715 37703 6721
rect 37645 6712 37657 6715
rect 37323 6684 37657 6712
rect 37323 6681 37335 6684
rect 37277 6675 37335 6681
rect 37645 6681 37657 6684
rect 37691 6681 37703 6715
rect 37645 6675 37703 6681
rect 38378 6672 38384 6724
rect 38436 6672 38442 6724
rect 38948 6644 38976 6752
rect 42153 6749 42165 6783
rect 42199 6780 42211 6783
rect 44082 6780 44088 6792
rect 42199 6752 44088 6780
rect 42199 6749 42211 6752
rect 42153 6743 42211 6749
rect 44082 6740 44088 6752
rect 44140 6740 44146 6792
rect 39574 6672 39580 6724
rect 39632 6712 39638 6724
rect 40221 6715 40279 6721
rect 40221 6712 40233 6715
rect 39632 6684 40233 6712
rect 39632 6672 39638 6684
rect 40221 6681 40233 6684
rect 40267 6681 40279 6715
rect 40221 6675 40279 6681
rect 40405 6715 40463 6721
rect 40405 6681 40417 6715
rect 40451 6712 40463 6715
rect 43346 6712 43352 6724
rect 40451 6684 43352 6712
rect 40451 6681 40463 6684
rect 40405 6675 40463 6681
rect 43346 6672 43352 6684
rect 43404 6672 43410 6724
rect 36280 6616 38976 6644
rect 39114 6604 39120 6656
rect 39172 6644 39178 6656
rect 39485 6647 39543 6653
rect 39485 6644 39497 6647
rect 39172 6616 39497 6644
rect 39172 6604 39178 6616
rect 39485 6613 39497 6616
rect 39531 6613 39543 6647
rect 39485 6607 39543 6613
rect 40586 6604 40592 6656
rect 40644 6604 40650 6656
rect 41414 6604 41420 6656
rect 41472 6604 41478 6656
rect 41506 6604 41512 6656
rect 41564 6604 41570 6656
rect 41782 6604 41788 6656
rect 41840 6644 41846 6656
rect 42245 6647 42303 6653
rect 42245 6644 42257 6647
rect 41840 6616 42257 6644
rect 41840 6604 41846 6616
rect 42245 6613 42257 6616
rect 42291 6613 42303 6647
rect 42245 6607 42303 6613
rect 2024 6554 77924 6576
rect 2024 6502 5794 6554
rect 5846 6502 5858 6554
rect 5910 6502 5922 6554
rect 5974 6502 5986 6554
rect 6038 6502 6050 6554
rect 6102 6502 36514 6554
rect 36566 6502 36578 6554
rect 36630 6502 36642 6554
rect 36694 6502 36706 6554
rect 36758 6502 36770 6554
rect 36822 6502 67234 6554
rect 67286 6502 67298 6554
rect 67350 6502 67362 6554
rect 67414 6502 67426 6554
rect 67478 6502 67490 6554
rect 67542 6502 77924 6554
rect 2024 6480 77924 6502
rect 7006 6400 7012 6452
rect 7064 6440 7070 6452
rect 10686 6440 10692 6452
rect 7064 6412 10692 6440
rect 7064 6400 7070 6412
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 13354 6440 13360 6452
rect 11664 6412 13360 6440
rect 11664 6400 11670 6412
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 13725 6443 13783 6449
rect 13725 6409 13737 6443
rect 13771 6440 13783 6443
rect 15654 6440 15660 6452
rect 13771 6412 15660 6440
rect 13771 6409 13783 6412
rect 13725 6403 13783 6409
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 15933 6443 15991 6449
rect 15933 6409 15945 6443
rect 15979 6440 15991 6443
rect 16114 6440 16120 6452
rect 15979 6412 16120 6440
rect 15979 6409 15991 6412
rect 15933 6403 15991 6409
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 16666 6400 16672 6452
rect 16724 6400 16730 6452
rect 18414 6400 18420 6452
rect 18472 6400 18478 6452
rect 20806 6440 20812 6452
rect 19996 6412 20812 6440
rect 10594 6332 10600 6384
rect 10652 6372 10658 6384
rect 13630 6372 13636 6384
rect 10652 6344 13636 6372
rect 10652 6332 10658 6344
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 16761 6375 16819 6381
rect 16761 6372 16773 6375
rect 14476 6344 16773 6372
rect 8110 6264 8116 6316
rect 8168 6304 8174 6316
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 8168 6276 9689 6304
rect 8168 6264 8174 6276
rect 9677 6273 9689 6276
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 12161 6307 12219 6313
rect 12161 6304 12173 6307
rect 10827 6276 12173 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 12161 6273 12173 6276
rect 12207 6273 12219 6307
rect 12161 6267 12219 6273
rect 12710 6264 12716 6316
rect 12768 6264 12774 6316
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6304 13967 6307
rect 14476 6304 14504 6344
rect 16761 6341 16773 6344
rect 16807 6341 16819 6375
rect 16761 6335 16819 6341
rect 18325 6375 18383 6381
rect 18325 6341 18337 6375
rect 18371 6372 18383 6375
rect 19996 6372 20024 6412
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 21082 6400 21088 6452
rect 21140 6440 21146 6452
rect 21729 6443 21787 6449
rect 21729 6440 21741 6443
rect 21140 6412 21741 6440
rect 21140 6400 21146 6412
rect 21729 6409 21741 6412
rect 21775 6409 21787 6443
rect 23753 6443 23811 6449
rect 23753 6440 23765 6443
rect 21729 6403 21787 6409
rect 22020 6412 23765 6440
rect 21634 6372 21640 6384
rect 18371 6344 20024 6372
rect 20656 6344 21640 6372
rect 18371 6341 18383 6344
rect 18325 6335 18383 6341
rect 13955 6276 14504 6304
rect 13955 6273 13967 6276
rect 13909 6267 13967 6273
rect 14550 6264 14556 6316
rect 14608 6264 14614 6316
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 16390 6304 16396 6316
rect 16163 6276 16396 6304
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 17773 6307 17831 6313
rect 17773 6273 17785 6307
rect 17819 6304 17831 6307
rect 19334 6304 19340 6316
rect 17819 6276 19340 6304
rect 17819 6273 17831 6276
rect 17773 6267 17831 6273
rect 19334 6264 19340 6276
rect 19392 6264 19398 6316
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 19889 6307 19947 6313
rect 19889 6304 19901 6307
rect 19484 6276 19901 6304
rect 19484 6264 19490 6276
rect 19889 6273 19901 6276
rect 19935 6273 19947 6307
rect 20656 6304 20684 6344
rect 21634 6332 21640 6344
rect 21692 6332 21698 6384
rect 19889 6267 19947 6273
rect 20180 6276 20684 6304
rect 20717 6307 20775 6313
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 10321 6239 10379 6245
rect 10321 6236 10333 6239
rect 8996 6208 10333 6236
rect 8996 6196 9002 6208
rect 10321 6205 10333 6208
rect 10367 6205 10379 6239
rect 10321 6199 10379 6205
rect 11333 6239 11391 6245
rect 11333 6205 11345 6239
rect 11379 6236 11391 6239
rect 12250 6236 12256 6248
rect 11379 6208 12256 6236
rect 11379 6205 11391 6208
rect 11333 6199 11391 6205
rect 12250 6196 12256 6208
rect 12308 6196 12314 6248
rect 13173 6239 13231 6245
rect 13173 6205 13185 6239
rect 13219 6236 13231 6239
rect 15194 6236 15200 6248
rect 13219 6208 15200 6236
rect 13219 6205 13231 6208
rect 13173 6199 13231 6205
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6236 15439 6239
rect 16574 6236 16580 6248
rect 15427 6208 16580 6236
rect 15427 6205 15439 6208
rect 15381 6199 15439 6205
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 17313 6239 17371 6245
rect 17313 6205 17325 6239
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 3786 6128 3792 6180
rect 3844 6168 3850 6180
rect 11790 6168 11796 6180
rect 3844 6140 11796 6168
rect 3844 6128 3850 6140
rect 11790 6128 11796 6140
rect 11848 6128 11854 6180
rect 11882 6128 11888 6180
rect 11940 6168 11946 6180
rect 17328 6168 17356 6199
rect 18138 6196 18144 6248
rect 18196 6236 18202 6248
rect 18598 6236 18604 6248
rect 18196 6208 18604 6236
rect 18196 6196 18202 6208
rect 18598 6196 18604 6208
rect 18656 6196 18662 6248
rect 18969 6239 19027 6245
rect 18969 6205 18981 6239
rect 19015 6205 19027 6239
rect 18969 6199 19027 6205
rect 11940 6140 17356 6168
rect 11940 6128 11946 6140
rect 17586 6128 17592 6180
rect 17644 6168 17650 6180
rect 18984 6168 19012 6199
rect 19150 6196 19156 6248
rect 19208 6196 19214 6248
rect 19794 6196 19800 6248
rect 19852 6236 19858 6248
rect 20180 6236 20208 6276
rect 20717 6273 20729 6307
rect 20763 6304 20775 6307
rect 22020 6304 22048 6412
rect 23753 6409 23765 6412
rect 23799 6409 23811 6443
rect 23753 6403 23811 6409
rect 24394 6400 24400 6452
rect 24452 6440 24458 6452
rect 24670 6440 24676 6452
rect 24452 6412 24676 6440
rect 24452 6400 24458 6412
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 25133 6443 25191 6449
rect 25133 6409 25145 6443
rect 25179 6440 25191 6443
rect 25774 6440 25780 6452
rect 25179 6412 25780 6440
rect 25179 6409 25191 6412
rect 25133 6403 25191 6409
rect 25774 6400 25780 6412
rect 25832 6400 25838 6452
rect 26050 6400 26056 6452
rect 26108 6440 26114 6452
rect 26881 6443 26939 6449
rect 26881 6440 26893 6443
rect 26108 6412 26893 6440
rect 26108 6400 26114 6412
rect 26881 6409 26893 6412
rect 26927 6409 26939 6443
rect 26881 6403 26939 6409
rect 27246 6400 27252 6452
rect 27304 6400 27310 6452
rect 27341 6443 27399 6449
rect 27341 6409 27353 6443
rect 27387 6440 27399 6443
rect 27890 6440 27896 6452
rect 27387 6412 27896 6440
rect 27387 6409 27399 6412
rect 27341 6403 27399 6409
rect 27890 6400 27896 6412
rect 27948 6400 27954 6452
rect 28813 6443 28871 6449
rect 28813 6409 28825 6443
rect 28859 6440 28871 6443
rect 28902 6440 28908 6452
rect 28859 6412 28908 6440
rect 28859 6409 28871 6412
rect 28813 6403 28871 6409
rect 28902 6400 28908 6412
rect 28960 6400 28966 6452
rect 30282 6400 30288 6452
rect 30340 6400 30346 6452
rect 30374 6400 30380 6452
rect 30432 6440 30438 6452
rect 34146 6440 34152 6452
rect 30432 6412 34152 6440
rect 30432 6400 30438 6412
rect 22189 6375 22247 6381
rect 22189 6372 22201 6375
rect 20763 6276 22048 6304
rect 22112 6344 22201 6372
rect 20763 6273 20775 6276
rect 20717 6267 20775 6273
rect 19852 6208 20208 6236
rect 19852 6196 19858 6208
rect 20254 6196 20260 6248
rect 20312 6236 20318 6248
rect 21821 6239 21879 6245
rect 21821 6236 21833 6239
rect 20312 6208 21833 6236
rect 20312 6196 20318 6208
rect 21821 6205 21833 6208
rect 21867 6205 21879 6239
rect 21821 6199 21879 6205
rect 22002 6196 22008 6248
rect 22060 6196 22066 6248
rect 22112 6236 22140 6344
rect 22189 6341 22201 6344
rect 22235 6341 22247 6375
rect 22189 6335 22247 6341
rect 22405 6375 22463 6381
rect 22405 6341 22417 6375
rect 22451 6372 22463 6375
rect 22646 6372 22652 6384
rect 22451 6344 22652 6372
rect 22451 6341 22463 6344
rect 22405 6335 22463 6341
rect 22646 6332 22652 6344
rect 22704 6332 22710 6384
rect 28166 6372 28172 6384
rect 24044 6344 28172 6372
rect 22741 6307 22799 6313
rect 22741 6304 22753 6307
rect 22664 6276 22753 6304
rect 22664 6248 22692 6276
rect 22741 6273 22753 6276
rect 22787 6273 22799 6307
rect 23750 6304 23756 6316
rect 22741 6267 22799 6273
rect 22848 6276 23756 6304
rect 22186 6236 22192 6248
rect 22112 6208 22192 6236
rect 22186 6196 22192 6208
rect 22244 6236 22250 6248
rect 22554 6236 22560 6248
rect 22244 6208 22560 6236
rect 22244 6196 22250 6208
rect 22554 6196 22560 6208
rect 22612 6196 22618 6248
rect 22646 6196 22652 6248
rect 22704 6196 22710 6248
rect 20533 6171 20591 6177
rect 17644 6140 18920 6168
rect 18984 6140 20484 6168
rect 17644 6128 17650 6140
rect 7926 6060 7932 6112
rect 7984 6100 7990 6112
rect 9493 6103 9551 6109
rect 9493 6100 9505 6103
rect 7984 6072 9505 6100
rect 7984 6060 7990 6072
rect 9493 6069 9505 6072
rect 9539 6069 9551 6103
rect 9493 6063 9551 6069
rect 9766 6060 9772 6112
rect 9824 6060 9830 6112
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 11609 6103 11667 6109
rect 11609 6100 11621 6103
rect 9916 6072 11621 6100
rect 9916 6060 9922 6072
rect 11609 6069 11621 6072
rect 11655 6069 11667 6103
rect 11609 6063 11667 6069
rect 12710 6060 12716 6112
rect 12768 6060 12774 6112
rect 14461 6103 14519 6109
rect 14461 6069 14473 6103
rect 14507 6100 14519 6103
rect 14642 6100 14648 6112
rect 14507 6072 14648 6100
rect 14507 6069 14519 6072
rect 14461 6063 14519 6069
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 15197 6103 15255 6109
rect 15197 6069 15209 6103
rect 15243 6100 15255 6103
rect 18690 6100 18696 6112
rect 15243 6072 18696 6100
rect 15243 6069 15255 6072
rect 15197 6063 15255 6069
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 18892 6100 18920 6140
rect 20254 6100 20260 6112
rect 18892 6072 20260 6100
rect 20254 6060 20260 6072
rect 20312 6060 20318 6112
rect 20456 6100 20484 6140
rect 20533 6137 20545 6171
rect 20579 6168 20591 6171
rect 22848 6168 22876 6276
rect 23750 6264 23756 6276
rect 23808 6264 23814 6316
rect 23109 6239 23167 6245
rect 23109 6205 23121 6239
rect 23155 6236 23167 6239
rect 23290 6236 23296 6248
rect 23155 6208 23296 6236
rect 23155 6205 23167 6208
rect 23109 6199 23167 6205
rect 23290 6196 23296 6208
rect 23348 6196 23354 6248
rect 23474 6196 23480 6248
rect 23532 6236 23538 6248
rect 24044 6236 24072 6344
rect 28166 6332 28172 6344
rect 28224 6332 28230 6384
rect 31478 6372 31484 6384
rect 28736 6344 31484 6372
rect 24118 6264 24124 6316
rect 24176 6304 24182 6316
rect 25225 6307 25283 6313
rect 25225 6304 25237 6307
rect 24176 6276 25237 6304
rect 24176 6264 24182 6276
rect 25225 6273 25237 6276
rect 25271 6273 25283 6307
rect 25225 6267 25283 6273
rect 25406 6264 25412 6316
rect 25464 6304 25470 6316
rect 25682 6304 25688 6316
rect 25464 6276 25688 6304
rect 25464 6264 25470 6276
rect 25682 6264 25688 6276
rect 25740 6264 25746 6316
rect 26510 6264 26516 6316
rect 26568 6264 26574 6316
rect 27448 6276 28212 6304
rect 23532 6208 24072 6236
rect 23532 6196 23538 6208
rect 24394 6196 24400 6248
rect 24452 6196 24458 6248
rect 24489 6239 24547 6245
rect 24489 6205 24501 6239
rect 24535 6205 24547 6239
rect 24489 6199 24547 6205
rect 20579 6140 22876 6168
rect 22925 6171 22983 6177
rect 20579 6137 20591 6140
rect 20533 6131 20591 6137
rect 22925 6137 22937 6171
rect 22971 6168 22983 6171
rect 24504 6168 24532 6199
rect 25774 6196 25780 6248
rect 25832 6196 25838 6248
rect 25866 6196 25872 6248
rect 25924 6236 25930 6248
rect 27448 6236 27476 6276
rect 25924 6208 27476 6236
rect 25924 6196 25930 6208
rect 27522 6196 27528 6248
rect 27580 6196 27586 6248
rect 28184 6236 28212 6276
rect 28258 6264 28264 6316
rect 28316 6264 28322 6316
rect 28736 6236 28764 6344
rect 31478 6332 31484 6344
rect 31536 6332 31542 6384
rect 31846 6332 31852 6384
rect 31904 6332 31910 6384
rect 32122 6332 32128 6384
rect 32180 6372 32186 6384
rect 32677 6375 32735 6381
rect 32677 6372 32689 6375
rect 32180 6344 32689 6372
rect 32180 6332 32186 6344
rect 32677 6341 32689 6344
rect 32723 6341 32735 6375
rect 32677 6335 32735 6341
rect 29733 6307 29791 6313
rect 29733 6273 29745 6307
rect 29779 6304 29791 6307
rect 30098 6304 30104 6316
rect 29779 6276 30104 6304
rect 29779 6273 29791 6276
rect 29733 6267 29791 6273
rect 30098 6264 30104 6276
rect 30156 6264 30162 6316
rect 30466 6264 30472 6316
rect 30524 6264 30530 6316
rect 31757 6307 31815 6313
rect 31757 6273 31769 6307
rect 31803 6304 31815 6307
rect 31938 6304 31944 6316
rect 31803 6276 31944 6304
rect 31803 6273 31815 6276
rect 31757 6267 31815 6273
rect 31938 6264 31944 6276
rect 31996 6264 32002 6316
rect 32214 6264 32220 6316
rect 32272 6304 32278 6316
rect 33060 6313 33088 6412
rect 34146 6400 34152 6412
rect 34204 6400 34210 6452
rect 34238 6400 34244 6452
rect 34296 6440 34302 6452
rect 35986 6440 35992 6452
rect 34296 6412 35992 6440
rect 34296 6400 34302 6412
rect 35986 6400 35992 6412
rect 36044 6400 36050 6452
rect 36354 6400 36360 6452
rect 36412 6440 36418 6452
rect 36541 6443 36599 6449
rect 36541 6440 36553 6443
rect 36412 6412 36553 6440
rect 36412 6400 36418 6412
rect 36541 6409 36553 6412
rect 36587 6409 36599 6443
rect 36541 6403 36599 6409
rect 38608 6400 38614 6452
rect 38666 6440 38672 6452
rect 40586 6440 40592 6452
rect 38666 6412 40592 6440
rect 38666 6400 38672 6412
rect 40586 6400 40592 6412
rect 40644 6400 40650 6452
rect 40862 6400 40868 6452
rect 40920 6440 40926 6452
rect 40920 6412 43024 6440
rect 40920 6400 40926 6412
rect 33226 6332 33232 6384
rect 33284 6372 33290 6384
rect 33321 6375 33379 6381
rect 33321 6372 33333 6375
rect 33284 6344 33333 6372
rect 33284 6332 33290 6344
rect 33321 6341 33333 6344
rect 33367 6341 33379 6375
rect 33321 6335 33379 6341
rect 33778 6332 33784 6384
rect 33836 6332 33842 6384
rect 34606 6332 34612 6384
rect 34664 6372 34670 6384
rect 35069 6375 35127 6381
rect 35069 6372 35081 6375
rect 34664 6344 35081 6372
rect 34664 6332 34670 6344
rect 35069 6341 35081 6344
rect 35115 6341 35127 6375
rect 37369 6375 37427 6381
rect 37369 6372 37381 6375
rect 35069 6335 35127 6341
rect 36096 6344 37381 6372
rect 32585 6307 32643 6313
rect 32585 6304 32597 6307
rect 32272 6276 32597 6304
rect 32272 6264 32278 6276
rect 32585 6273 32597 6276
rect 32631 6273 32643 6307
rect 32585 6267 32643 6273
rect 33045 6307 33103 6313
rect 33045 6273 33057 6307
rect 33091 6273 33103 6307
rect 33045 6267 33103 6273
rect 35434 6264 35440 6316
rect 35492 6304 35498 6316
rect 36096 6313 36124 6344
rect 37369 6341 37381 6344
rect 37415 6341 37427 6375
rect 37369 6335 37427 6341
rect 38378 6332 38384 6384
rect 38436 6372 38442 6384
rect 38930 6372 38936 6384
rect 38436 6344 38936 6372
rect 38436 6332 38442 6344
rect 38930 6332 38936 6344
rect 38988 6332 38994 6384
rect 40494 6372 40500 6384
rect 39776 6344 40500 6372
rect 35897 6307 35955 6313
rect 35897 6304 35909 6307
rect 35492 6276 35909 6304
rect 35492 6264 35498 6276
rect 35897 6273 35909 6276
rect 35943 6273 35955 6307
rect 35897 6267 35955 6273
rect 36081 6307 36139 6313
rect 36081 6273 36093 6307
rect 36127 6273 36139 6307
rect 36081 6267 36139 6273
rect 36170 6264 36176 6316
rect 36228 6264 36234 6316
rect 36262 6264 36268 6316
rect 36320 6264 36326 6316
rect 37826 6264 37832 6316
rect 37884 6304 37890 6316
rect 37921 6307 37979 6313
rect 37921 6304 37933 6307
rect 37884 6276 37933 6304
rect 37884 6264 37890 6276
rect 37921 6273 37933 6276
rect 37967 6273 37979 6307
rect 37921 6267 37979 6273
rect 38194 6264 38200 6316
rect 38252 6264 38258 6316
rect 28184 6208 28764 6236
rect 28810 6196 28816 6248
rect 28868 6236 28874 6248
rect 29457 6239 29515 6245
rect 29457 6236 29469 6239
rect 28868 6208 29469 6236
rect 28868 6196 28874 6208
rect 29457 6205 29469 6208
rect 29503 6205 29515 6239
rect 29457 6199 29515 6205
rect 29822 6196 29828 6248
rect 29880 6236 29886 6248
rect 31113 6239 31171 6245
rect 31113 6236 31125 6239
rect 29880 6208 31125 6236
rect 29880 6196 29886 6208
rect 31113 6205 31125 6208
rect 31159 6205 31171 6239
rect 32401 6239 32459 6245
rect 32401 6236 32413 6239
rect 31113 6199 31171 6205
rect 31220 6208 32413 6236
rect 22971 6140 24532 6168
rect 22971 6137 22983 6140
rect 22925 6131 22983 6137
rect 25498 6128 25504 6180
rect 25556 6168 25562 6180
rect 28905 6171 28963 6177
rect 28905 6168 28917 6171
rect 25556 6140 28917 6168
rect 25556 6128 25562 6140
rect 28905 6137 28917 6140
rect 28951 6137 28963 6171
rect 28905 6131 28963 6137
rect 30466 6128 30472 6180
rect 30524 6168 30530 6180
rect 31220 6168 31248 6208
rect 32401 6205 32413 6208
rect 32447 6205 32459 6239
rect 32401 6199 32459 6205
rect 32508 6208 35664 6236
rect 30524 6140 31248 6168
rect 30524 6128 30530 6140
rect 32214 6128 32220 6180
rect 32272 6168 32278 6180
rect 32508 6168 32536 6208
rect 35636 6168 35664 6208
rect 35710 6196 35716 6248
rect 35768 6196 35774 6248
rect 37274 6196 37280 6248
rect 37332 6196 37338 6248
rect 38473 6239 38531 6245
rect 38473 6236 38485 6239
rect 38304 6208 38485 6236
rect 32272 6140 32536 6168
rect 32600 6140 32904 6168
rect 35636 6140 37044 6168
rect 32272 6128 32278 6140
rect 21082 6100 21088 6112
rect 20456 6072 21088 6100
rect 21082 6060 21088 6072
rect 21140 6060 21146 6112
rect 21266 6060 21272 6112
rect 21324 6060 21330 6112
rect 21358 6060 21364 6112
rect 21416 6060 21422 6112
rect 21450 6060 21456 6112
rect 21508 6100 21514 6112
rect 21634 6100 21640 6112
rect 21508 6072 21640 6100
rect 21508 6060 21514 6072
rect 21634 6060 21640 6072
rect 21692 6060 21698 6112
rect 22002 6060 22008 6112
rect 22060 6100 22066 6112
rect 22186 6100 22192 6112
rect 22060 6072 22192 6100
rect 22060 6060 22066 6072
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 22278 6060 22284 6112
rect 22336 6100 22342 6112
rect 22373 6103 22431 6109
rect 22373 6100 22385 6103
rect 22336 6072 22385 6100
rect 22336 6060 22342 6072
rect 22373 6069 22385 6072
rect 22419 6069 22431 6103
rect 22373 6063 22431 6069
rect 22554 6060 22560 6112
rect 22612 6060 22618 6112
rect 23661 6103 23719 6109
rect 23661 6069 23673 6103
rect 23707 6100 23719 6103
rect 25038 6100 25044 6112
rect 23707 6072 25044 6100
rect 23707 6069 23719 6072
rect 23661 6063 23719 6069
rect 25038 6060 25044 6072
rect 25096 6060 25102 6112
rect 25314 6060 25320 6112
rect 25372 6100 25378 6112
rect 25961 6103 26019 6109
rect 25961 6100 25973 6103
rect 25372 6072 25973 6100
rect 25372 6060 25378 6072
rect 25961 6069 25973 6072
rect 26007 6069 26019 6103
rect 25961 6063 26019 6069
rect 27430 6060 27436 6112
rect 27488 6100 27494 6112
rect 30834 6100 30840 6112
rect 27488 6072 30840 6100
rect 27488 6060 27494 6072
rect 30834 6060 30840 6072
rect 30892 6060 30898 6112
rect 31021 6103 31079 6109
rect 31021 6069 31033 6103
rect 31067 6100 31079 6103
rect 32600 6100 32628 6140
rect 31067 6072 32628 6100
rect 32876 6100 32904 6140
rect 33870 6100 33876 6112
rect 32876 6072 33876 6100
rect 31067 6069 31079 6072
rect 31021 6063 31079 6069
rect 33870 6060 33876 6072
rect 33928 6060 33934 6112
rect 35161 6103 35219 6109
rect 35161 6069 35173 6103
rect 35207 6100 35219 6103
rect 35434 6100 35440 6112
rect 35207 6072 35440 6100
rect 35207 6069 35219 6072
rect 35161 6063 35219 6069
rect 35434 6060 35440 6072
rect 35492 6060 35498 6112
rect 36633 6103 36691 6109
rect 36633 6069 36645 6103
rect 36679 6100 36691 6103
rect 36906 6100 36912 6112
rect 36679 6072 36912 6100
rect 36679 6069 36691 6072
rect 36633 6063 36691 6069
rect 36906 6060 36912 6072
rect 36964 6060 36970 6112
rect 37016 6100 37044 6140
rect 37550 6128 37556 6180
rect 37608 6168 37614 6180
rect 38304 6168 38332 6208
rect 38473 6205 38485 6208
rect 38519 6205 38531 6239
rect 38473 6199 38531 6205
rect 38562 6196 38568 6248
rect 38620 6236 38626 6248
rect 39776 6236 39804 6344
rect 40494 6332 40500 6344
rect 40552 6372 40558 6384
rect 42518 6372 42524 6384
rect 40552 6344 42524 6372
rect 40552 6332 40558 6344
rect 42518 6332 42524 6344
rect 42576 6372 42582 6384
rect 42797 6375 42855 6381
rect 42797 6372 42809 6375
rect 42576 6344 42809 6372
rect 42576 6332 42582 6344
rect 42797 6341 42809 6344
rect 42843 6341 42855 6375
rect 42797 6335 42855 6341
rect 41414 6264 41420 6316
rect 41472 6304 41478 6316
rect 42996 6313 43024 6412
rect 41785 6307 41843 6313
rect 41785 6304 41797 6307
rect 41472 6276 41797 6304
rect 41472 6264 41478 6276
rect 41785 6273 41797 6276
rect 41831 6273 41843 6307
rect 42705 6307 42763 6313
rect 42705 6304 42717 6307
rect 41785 6267 41843 6273
rect 41892 6276 42717 6304
rect 38620 6208 39804 6236
rect 38620 6196 38626 6208
rect 40218 6196 40224 6248
rect 40276 6196 40282 6248
rect 40589 6239 40647 6245
rect 40589 6205 40601 6239
rect 40635 6236 40647 6239
rect 41233 6239 41291 6245
rect 41233 6236 41245 6239
rect 40635 6208 41245 6236
rect 40635 6205 40647 6208
rect 40589 6199 40647 6205
rect 41233 6205 41245 6208
rect 41279 6205 41291 6239
rect 41233 6199 41291 6205
rect 41322 6196 41328 6248
rect 41380 6236 41386 6248
rect 41892 6236 41920 6276
rect 42705 6273 42717 6276
rect 42751 6273 42763 6307
rect 42705 6267 42763 6273
rect 42981 6307 43039 6313
rect 42981 6273 42993 6307
rect 43027 6304 43039 6307
rect 43070 6304 43076 6316
rect 43027 6276 43076 6304
rect 43027 6273 43039 6276
rect 42981 6267 43039 6273
rect 43070 6264 43076 6276
rect 43128 6264 43134 6316
rect 41380 6208 41920 6236
rect 41380 6196 41386 6208
rect 41966 6196 41972 6248
rect 42024 6196 42030 6248
rect 37608 6140 38332 6168
rect 37608 6128 37614 6140
rect 39850 6100 39856 6112
rect 37016 6072 39856 6100
rect 39850 6060 39856 6072
rect 39908 6060 39914 6112
rect 41138 6060 41144 6112
rect 41196 6060 41202 6112
rect 42610 6060 42616 6112
rect 42668 6060 42674 6112
rect 42794 6060 42800 6112
rect 42852 6100 42858 6112
rect 43165 6103 43223 6109
rect 43165 6100 43177 6103
rect 42852 6072 43177 6100
rect 42852 6060 42858 6072
rect 43165 6069 43177 6072
rect 43211 6069 43223 6103
rect 43165 6063 43223 6069
rect 2024 6010 77924 6032
rect 2024 5958 5134 6010
rect 5186 5958 5198 6010
rect 5250 5958 5262 6010
rect 5314 5958 5326 6010
rect 5378 5958 5390 6010
rect 5442 5958 35854 6010
rect 35906 5958 35918 6010
rect 35970 5958 35982 6010
rect 36034 5958 36046 6010
rect 36098 5958 36110 6010
rect 36162 5958 66574 6010
rect 66626 5958 66638 6010
rect 66690 5958 66702 6010
rect 66754 5958 66766 6010
rect 66818 5958 66830 6010
rect 66882 5958 77924 6010
rect 2024 5936 77924 5958
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 9766 5896 9772 5908
rect 3660 5868 9772 5896
rect 3660 5856 3666 5868
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 10134 5856 10140 5908
rect 10192 5856 10198 5908
rect 11146 5856 11152 5908
rect 11204 5856 11210 5908
rect 12434 5896 12440 5908
rect 11256 5868 12440 5896
rect 7558 5788 7564 5840
rect 7616 5828 7622 5840
rect 9858 5828 9864 5840
rect 7616 5800 9864 5828
rect 7616 5788 7622 5800
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 7834 5720 7840 5772
rect 7892 5760 7898 5772
rect 11256 5760 11284 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 14093 5899 14151 5905
rect 12728 5868 14044 5896
rect 12728 5760 12756 5868
rect 14016 5828 14044 5868
rect 14093 5865 14105 5899
rect 14139 5896 14151 5899
rect 14458 5896 14464 5908
rect 14139 5868 14464 5896
rect 14139 5865 14151 5868
rect 14093 5859 14151 5865
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 14829 5899 14887 5905
rect 14829 5865 14841 5899
rect 14875 5896 14887 5899
rect 15102 5896 15108 5908
rect 14875 5868 15108 5896
rect 14875 5865 14887 5868
rect 14829 5859 14887 5865
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 18414 5896 18420 5908
rect 16408 5868 18420 5896
rect 15562 5828 15568 5840
rect 14016 5800 15568 5828
rect 15562 5788 15568 5800
rect 15620 5788 15626 5840
rect 7892 5732 11284 5760
rect 12406 5732 12756 5760
rect 12805 5763 12863 5769
rect 7892 5720 7898 5732
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 9585 5695 9643 5701
rect 9585 5692 9597 5695
rect 8352 5664 9597 5692
rect 8352 5652 8358 5664
rect 9585 5661 9597 5664
rect 9631 5661 9643 5695
rect 9585 5655 9643 5661
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 8018 5584 8024 5636
rect 8076 5624 8082 5636
rect 9968 5624 9996 5655
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 10505 5695 10563 5701
rect 10505 5692 10517 5695
rect 10376 5664 10517 5692
rect 10376 5652 10382 5664
rect 10505 5661 10517 5664
rect 10551 5661 10563 5695
rect 10505 5655 10563 5661
rect 10686 5652 10692 5704
rect 10744 5692 10750 5704
rect 11330 5692 11336 5704
rect 10744 5664 11336 5692
rect 10744 5652 10750 5664
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 11422 5652 11428 5704
rect 11480 5652 11486 5704
rect 11514 5652 11520 5704
rect 11572 5652 11578 5704
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5692 11943 5695
rect 12406 5692 12434 5732
rect 12805 5729 12817 5763
rect 12851 5760 12863 5763
rect 16022 5760 16028 5772
rect 12851 5732 16028 5760
rect 12851 5729 12863 5732
rect 12805 5723 12863 5729
rect 16022 5720 16028 5732
rect 16080 5720 16086 5772
rect 16298 5720 16304 5772
rect 16356 5720 16362 5772
rect 11931 5664 12434 5692
rect 12529 5695 12587 5701
rect 11931 5661 11943 5664
rect 11885 5655 11943 5661
rect 12529 5661 12541 5695
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 13814 5692 13820 5704
rect 13587 5664 13820 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 8076 5596 9996 5624
rect 11793 5627 11851 5633
rect 8076 5584 8082 5596
rect 11793 5593 11805 5627
rect 11839 5624 11851 5627
rect 12434 5624 12440 5636
rect 11839 5596 12440 5624
rect 11839 5593 11851 5596
rect 11793 5587 11851 5593
rect 12434 5584 12440 5596
rect 12492 5584 12498 5636
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 9033 5559 9091 5565
rect 9033 5556 9045 5559
rect 4764 5528 9045 5556
rect 4764 5516 4770 5528
rect 9033 5525 9045 5528
rect 9079 5525 9091 5559
rect 9033 5519 9091 5525
rect 9766 5516 9772 5568
rect 9824 5556 9830 5568
rect 11977 5559 12035 5565
rect 11977 5556 11989 5559
rect 9824 5528 11989 5556
rect 9824 5516 9830 5528
rect 11977 5525 11989 5528
rect 12023 5525 12035 5559
rect 11977 5519 12035 5525
rect 12066 5516 12072 5568
rect 12124 5556 12130 5568
rect 12544 5556 12572 5655
rect 13814 5652 13820 5664
rect 13872 5652 13878 5704
rect 14090 5652 14096 5704
rect 14148 5692 14154 5704
rect 14185 5695 14243 5701
rect 14185 5692 14197 5695
rect 14148 5664 14197 5692
rect 14148 5652 14154 5664
rect 14185 5661 14197 5664
rect 14231 5661 14243 5695
rect 15841 5695 15899 5701
rect 14185 5655 14243 5661
rect 14844 5664 15424 5692
rect 13357 5627 13415 5633
rect 13357 5593 13369 5627
rect 13403 5624 13415 5627
rect 14734 5624 14740 5636
rect 13403 5596 14740 5624
rect 13403 5593 13415 5596
rect 13357 5587 13415 5593
rect 14734 5584 14740 5596
rect 14792 5584 14798 5636
rect 12124 5528 12572 5556
rect 12124 5516 12130 5528
rect 13262 5516 13268 5568
rect 13320 5556 13326 5568
rect 14844 5556 14872 5664
rect 15286 5584 15292 5636
rect 15344 5584 15350 5636
rect 15396 5624 15424 5664
rect 15841 5661 15853 5695
rect 15887 5692 15899 5695
rect 16408 5692 16436 5868
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 18509 5899 18567 5905
rect 18509 5865 18521 5899
rect 18555 5896 18567 5899
rect 18598 5896 18604 5908
rect 18555 5868 18604 5896
rect 18555 5865 18567 5868
rect 18509 5859 18567 5865
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 19245 5899 19303 5905
rect 19245 5865 19257 5899
rect 19291 5896 19303 5899
rect 19426 5896 19432 5908
rect 19291 5868 19432 5896
rect 19291 5865 19303 5868
rect 19245 5859 19303 5865
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 20533 5899 20591 5905
rect 20533 5896 20545 5899
rect 19576 5868 20545 5896
rect 19576 5856 19582 5868
rect 20533 5865 20545 5868
rect 20579 5865 20591 5899
rect 20533 5859 20591 5865
rect 20717 5899 20775 5905
rect 20717 5865 20729 5899
rect 20763 5896 20775 5899
rect 21174 5896 21180 5908
rect 20763 5868 21180 5896
rect 20763 5865 20775 5868
rect 20717 5859 20775 5865
rect 21174 5856 21180 5868
rect 21232 5856 21238 5908
rect 22922 5896 22928 5908
rect 21284 5868 22928 5896
rect 16482 5788 16488 5840
rect 16540 5828 16546 5840
rect 21284 5828 21312 5868
rect 22922 5856 22928 5868
rect 22980 5856 22986 5908
rect 24762 5896 24768 5908
rect 23032 5868 24768 5896
rect 16540 5800 21312 5828
rect 16540 5788 16546 5800
rect 21726 5788 21732 5840
rect 21784 5828 21790 5840
rect 23032 5828 23060 5868
rect 24762 5856 24768 5868
rect 24820 5856 24826 5908
rect 25133 5899 25191 5905
rect 25133 5865 25145 5899
rect 25179 5896 25191 5899
rect 27522 5896 27528 5908
rect 25179 5868 27528 5896
rect 25179 5865 25191 5868
rect 25133 5859 25191 5865
rect 27522 5856 27528 5868
rect 27580 5856 27586 5908
rect 33778 5896 33784 5908
rect 30300 5868 33784 5896
rect 23474 5828 23480 5840
rect 21784 5800 23060 5828
rect 23124 5800 23480 5828
rect 21784 5788 21790 5800
rect 17037 5763 17095 5769
rect 17037 5729 17049 5763
rect 17083 5760 17095 5763
rect 19150 5760 19156 5772
rect 17083 5732 19156 5760
rect 17083 5729 17095 5732
rect 17037 5723 17095 5729
rect 19150 5720 19156 5732
rect 19208 5720 19214 5772
rect 19334 5720 19340 5772
rect 19392 5720 19398 5772
rect 20438 5760 20444 5772
rect 20088 5732 20444 5760
rect 17129 5695 17187 5701
rect 17129 5692 17141 5695
rect 15887 5664 16436 5692
rect 16500 5664 17141 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 16500 5624 16528 5664
rect 17129 5661 17141 5664
rect 17175 5661 17187 5695
rect 17129 5655 17187 5661
rect 17678 5652 17684 5704
rect 17736 5692 17742 5704
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 17736 5664 17877 5692
rect 17736 5652 17742 5664
rect 17865 5661 17877 5664
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 18601 5695 18659 5701
rect 18601 5661 18613 5695
rect 18647 5661 18659 5695
rect 18601 5655 18659 5661
rect 15396 5596 16528 5624
rect 16574 5584 16580 5636
rect 16632 5624 16638 5636
rect 18616 5624 18644 5655
rect 18690 5652 18696 5704
rect 18748 5692 18754 5704
rect 20088 5692 20116 5732
rect 20438 5720 20444 5732
rect 20496 5720 20502 5772
rect 21637 5763 21695 5769
rect 21637 5729 21649 5763
rect 21683 5760 21695 5763
rect 21818 5760 21824 5772
rect 21683 5732 21824 5760
rect 21683 5729 21695 5732
rect 21637 5723 21695 5729
rect 21818 5720 21824 5732
rect 21876 5720 21882 5772
rect 22373 5763 22431 5769
rect 22373 5729 22385 5763
rect 22419 5760 22431 5763
rect 22462 5760 22468 5772
rect 22419 5732 22468 5760
rect 22419 5729 22431 5732
rect 22373 5723 22431 5729
rect 22462 5720 22468 5732
rect 22520 5720 22526 5772
rect 22925 5763 22983 5769
rect 22925 5729 22937 5763
rect 22971 5760 22983 5763
rect 23014 5760 23020 5772
rect 22971 5732 23020 5760
rect 22971 5729 22983 5732
rect 22925 5723 22983 5729
rect 23014 5720 23020 5732
rect 23072 5720 23078 5772
rect 23124 5769 23152 5800
rect 23474 5788 23480 5800
rect 23532 5788 23538 5840
rect 23661 5831 23719 5837
rect 23661 5797 23673 5831
rect 23707 5828 23719 5831
rect 23750 5828 23756 5840
rect 23707 5800 23756 5828
rect 23707 5797 23719 5800
rect 23661 5791 23719 5797
rect 23750 5788 23756 5800
rect 23808 5788 23814 5840
rect 23842 5788 23848 5840
rect 23900 5828 23906 5840
rect 24302 5828 24308 5840
rect 23900 5800 24308 5828
rect 23900 5788 23906 5800
rect 24302 5788 24308 5800
rect 24360 5788 24366 5840
rect 24397 5831 24455 5837
rect 24397 5797 24409 5831
rect 24443 5828 24455 5831
rect 26970 5828 26976 5840
rect 24443 5800 26976 5828
rect 24443 5797 24455 5800
rect 24397 5791 24455 5797
rect 26970 5788 26976 5800
rect 27028 5788 27034 5840
rect 28169 5831 28227 5837
rect 28169 5797 28181 5831
rect 28215 5797 28227 5831
rect 28169 5791 28227 5797
rect 23109 5763 23167 5769
rect 23109 5729 23121 5763
rect 23155 5729 23167 5763
rect 23109 5723 23167 5729
rect 23566 5720 23572 5772
rect 23624 5760 23630 5772
rect 28184 5760 28212 5791
rect 30300 5769 30328 5868
rect 33778 5856 33784 5868
rect 33836 5856 33842 5908
rect 34701 5899 34759 5905
rect 34701 5865 34713 5899
rect 34747 5896 34759 5899
rect 35250 5896 35256 5908
rect 34747 5868 35256 5896
rect 34747 5865 34759 5868
rect 34701 5859 34759 5865
rect 35250 5856 35256 5868
rect 35308 5856 35314 5908
rect 35710 5856 35716 5908
rect 35768 5896 35774 5908
rect 35986 5896 35992 5908
rect 35768 5868 35992 5896
rect 35768 5856 35774 5868
rect 35986 5856 35992 5868
rect 36044 5896 36050 5908
rect 36446 5896 36452 5908
rect 36044 5868 36452 5896
rect 36044 5856 36050 5868
rect 36446 5856 36452 5868
rect 36504 5856 36510 5908
rect 36817 5899 36875 5905
rect 36817 5865 36829 5899
rect 36863 5896 36875 5899
rect 37550 5896 37556 5908
rect 36863 5868 37556 5896
rect 36863 5865 36875 5868
rect 36817 5859 36875 5865
rect 37550 5856 37556 5868
rect 37608 5856 37614 5908
rect 38654 5856 38660 5908
rect 38712 5896 38718 5908
rect 39574 5896 39580 5908
rect 38712 5868 39580 5896
rect 38712 5856 38718 5868
rect 39574 5856 39580 5868
rect 39632 5856 39638 5908
rect 41509 5899 41567 5905
rect 41509 5865 41521 5899
rect 41555 5896 41567 5899
rect 41598 5896 41604 5908
rect 41555 5868 41604 5896
rect 41555 5865 41567 5868
rect 41509 5859 41567 5865
rect 41598 5856 41604 5868
rect 41656 5856 41662 5908
rect 32125 5831 32183 5837
rect 30760 5800 31984 5828
rect 30285 5763 30343 5769
rect 23624 5732 30236 5760
rect 23624 5720 23630 5732
rect 18748 5664 20116 5692
rect 20165 5695 20223 5701
rect 18748 5652 18754 5664
rect 20165 5661 20177 5695
rect 20211 5692 20223 5695
rect 20714 5692 20720 5704
rect 20211 5664 20720 5692
rect 20211 5661 20223 5664
rect 20165 5655 20223 5661
rect 20714 5652 20720 5664
rect 20772 5652 20778 5704
rect 20898 5652 20904 5704
rect 20956 5652 20962 5704
rect 22646 5692 22652 5704
rect 21008 5664 22652 5692
rect 21008 5624 21036 5664
rect 22646 5652 22652 5664
rect 22704 5652 22710 5704
rect 23750 5692 23756 5704
rect 23400 5664 23756 5692
rect 16632 5596 18644 5624
rect 18708 5596 21036 5624
rect 16632 5584 16638 5596
rect 13320 5528 14872 5556
rect 13320 5516 13326 5528
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 16025 5559 16083 5565
rect 16025 5556 16037 5559
rect 15252 5528 16037 5556
rect 15252 5516 15258 5528
rect 16025 5525 16037 5528
rect 16071 5556 16083 5559
rect 16298 5556 16304 5568
rect 16071 5528 16304 5556
rect 16071 5525 16083 5528
rect 16025 5519 16083 5525
rect 16298 5516 16304 5528
rect 16356 5516 16362 5568
rect 16390 5516 16396 5568
rect 16448 5516 16454 5568
rect 17773 5559 17831 5565
rect 17773 5525 17785 5559
rect 17819 5556 17831 5559
rect 17862 5556 17868 5568
rect 17819 5528 17868 5556
rect 17819 5525 17831 5528
rect 17773 5519 17831 5525
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18708 5556 18736 5596
rect 21266 5584 21272 5636
rect 21324 5624 21330 5636
rect 23400 5624 23428 5664
rect 23750 5652 23756 5664
rect 23808 5652 23814 5704
rect 23842 5652 23848 5704
rect 23900 5652 23906 5704
rect 24486 5652 24492 5704
rect 24544 5652 24550 5704
rect 25498 5652 25504 5704
rect 25556 5652 25562 5704
rect 25958 5652 25964 5704
rect 26016 5692 26022 5704
rect 26145 5695 26203 5701
rect 26145 5692 26157 5695
rect 26016 5664 26157 5692
rect 26016 5652 26022 5664
rect 26145 5661 26157 5664
rect 26191 5661 26203 5695
rect 26145 5655 26203 5661
rect 29549 5695 29607 5701
rect 29549 5661 29561 5695
rect 29595 5692 29607 5695
rect 30098 5692 30104 5704
rect 29595 5664 30104 5692
rect 29595 5661 29607 5664
rect 29549 5655 29607 5661
rect 30098 5652 30104 5664
rect 30156 5652 30162 5704
rect 30208 5692 30236 5732
rect 30285 5729 30297 5763
rect 30331 5729 30343 5763
rect 30285 5723 30343 5729
rect 30760 5692 30788 5800
rect 30834 5720 30840 5772
rect 30892 5760 30898 5772
rect 31021 5763 31079 5769
rect 31021 5760 31033 5763
rect 30892 5732 31033 5760
rect 30892 5720 30898 5732
rect 31021 5729 31033 5732
rect 31067 5729 31079 5763
rect 31021 5723 31079 5729
rect 30208 5664 30788 5692
rect 21324 5596 21680 5624
rect 21324 5584 21330 5596
rect 18012 5528 18736 5556
rect 18012 5516 18018 5528
rect 19426 5516 19432 5568
rect 19484 5556 19490 5568
rect 19981 5559 20039 5565
rect 19981 5556 19993 5559
rect 19484 5528 19993 5556
rect 19484 5516 19490 5528
rect 19981 5525 19993 5528
rect 20027 5525 20039 5559
rect 19981 5519 20039 5525
rect 20346 5516 20352 5568
rect 20404 5556 20410 5568
rect 20533 5559 20591 5565
rect 20533 5556 20545 5559
rect 20404 5528 20545 5556
rect 20404 5516 20410 5528
rect 20533 5525 20545 5528
rect 20579 5525 20591 5559
rect 20533 5519 20591 5525
rect 21358 5516 21364 5568
rect 21416 5556 21422 5568
rect 21453 5559 21511 5565
rect 21453 5556 21465 5559
rect 21416 5528 21465 5556
rect 21416 5516 21422 5528
rect 21453 5525 21465 5528
rect 21499 5525 21511 5559
rect 21652 5556 21680 5596
rect 22066 5596 23428 5624
rect 22066 5556 22094 5596
rect 23474 5584 23480 5636
rect 23532 5624 23538 5636
rect 26881 5627 26939 5633
rect 26881 5624 26893 5627
rect 23532 5596 26893 5624
rect 23532 5584 23538 5596
rect 26881 5593 26893 5596
rect 26927 5593 26939 5627
rect 26881 5587 26939 5593
rect 26970 5584 26976 5636
rect 27028 5624 27034 5636
rect 30837 5627 30895 5633
rect 30837 5624 30849 5627
rect 27028 5596 30849 5624
rect 27028 5584 27034 5596
rect 30837 5593 30849 5596
rect 30883 5593 30895 5627
rect 30837 5587 30895 5593
rect 21652 5528 22094 5556
rect 21453 5519 21511 5525
rect 22186 5516 22192 5568
rect 22244 5516 22250 5568
rect 22278 5516 22284 5568
rect 22336 5556 22342 5568
rect 22462 5556 22468 5568
rect 22336 5528 22468 5556
rect 22336 5516 22342 5528
rect 22462 5516 22468 5528
rect 22520 5516 22526 5568
rect 22554 5516 22560 5568
rect 22612 5556 22618 5568
rect 25406 5556 25412 5568
rect 22612 5528 25412 5556
rect 22612 5516 22618 5528
rect 25406 5516 25412 5528
rect 25464 5516 25470 5568
rect 26050 5516 26056 5568
rect 26108 5516 26114 5568
rect 26789 5559 26847 5565
rect 26789 5525 26801 5559
rect 26835 5556 26847 5559
rect 27246 5556 27252 5568
rect 26835 5528 27252 5556
rect 26835 5525 26847 5528
rect 26789 5519 26847 5525
rect 27246 5516 27252 5528
rect 27304 5516 27310 5568
rect 27890 5516 27896 5568
rect 27948 5556 27954 5568
rect 28905 5559 28963 5565
rect 28905 5556 28917 5559
rect 27948 5528 28917 5556
rect 27948 5516 27954 5528
rect 28905 5525 28917 5528
rect 28951 5525 28963 5559
rect 28905 5519 28963 5525
rect 29178 5516 29184 5568
rect 29236 5556 29242 5568
rect 29641 5559 29699 5565
rect 29641 5556 29653 5559
rect 29236 5528 29653 5556
rect 29236 5516 29242 5528
rect 29641 5525 29653 5528
rect 29687 5525 29699 5559
rect 29641 5519 29699 5525
rect 30190 5516 30196 5568
rect 30248 5556 30254 5568
rect 30469 5559 30527 5565
rect 30469 5556 30481 5559
rect 30248 5528 30481 5556
rect 30248 5516 30254 5528
rect 30469 5525 30481 5528
rect 30515 5525 30527 5559
rect 30469 5519 30527 5525
rect 30650 5516 30656 5568
rect 30708 5556 30714 5568
rect 30929 5559 30987 5565
rect 30929 5556 30941 5559
rect 30708 5528 30941 5556
rect 30708 5516 30714 5528
rect 30929 5525 30941 5528
rect 30975 5525 30987 5559
rect 31036 5556 31064 5723
rect 31202 5720 31208 5772
rect 31260 5760 31266 5772
rect 31956 5760 31984 5800
rect 32125 5797 32137 5831
rect 32171 5828 32183 5831
rect 33502 5828 33508 5840
rect 32171 5800 33508 5828
rect 32171 5797 32183 5800
rect 32125 5791 32183 5797
rect 33502 5788 33508 5800
rect 33560 5788 33566 5840
rect 34146 5828 34152 5840
rect 34072 5800 34152 5828
rect 34072 5769 34100 5800
rect 34146 5788 34152 5800
rect 34204 5788 34210 5840
rect 34256 5800 34468 5828
rect 34057 5763 34115 5769
rect 31260 5732 31892 5760
rect 31956 5732 32352 5760
rect 31260 5720 31266 5732
rect 31478 5652 31484 5704
rect 31536 5652 31542 5704
rect 31573 5695 31631 5701
rect 31573 5661 31585 5695
rect 31619 5692 31631 5695
rect 31662 5692 31668 5704
rect 31619 5664 31668 5692
rect 31619 5661 31631 5664
rect 31573 5655 31631 5661
rect 31662 5652 31668 5664
rect 31720 5652 31726 5704
rect 31864 5701 31892 5732
rect 31849 5695 31907 5701
rect 31849 5661 31861 5695
rect 31895 5661 31907 5695
rect 31849 5655 31907 5661
rect 31938 5652 31944 5704
rect 31996 5652 32002 5704
rect 31757 5627 31815 5633
rect 31757 5593 31769 5627
rect 31803 5624 31815 5627
rect 32214 5624 32220 5636
rect 31803 5596 32220 5624
rect 31803 5593 31815 5596
rect 31757 5587 31815 5593
rect 32214 5584 32220 5596
rect 32272 5584 32278 5636
rect 32324 5633 32352 5732
rect 34057 5729 34069 5763
rect 34103 5729 34115 5763
rect 34057 5723 34115 5729
rect 33686 5652 33692 5704
rect 33744 5692 33750 5704
rect 34149 5695 34207 5701
rect 34149 5692 34161 5695
rect 33744 5664 34161 5692
rect 33744 5652 33750 5664
rect 34149 5661 34161 5664
rect 34195 5661 34207 5695
rect 34149 5655 34207 5661
rect 32309 5627 32367 5633
rect 32309 5593 32321 5627
rect 32355 5624 32367 5627
rect 34256 5624 34284 5800
rect 34330 5720 34336 5772
rect 34388 5720 34394 5772
rect 34440 5760 34468 5800
rect 36262 5788 36268 5840
rect 36320 5828 36326 5840
rect 38841 5831 38899 5837
rect 38841 5828 38853 5831
rect 36320 5800 38853 5828
rect 36320 5788 36326 5800
rect 38841 5797 38853 5800
rect 38887 5797 38899 5831
rect 38841 5791 38899 5797
rect 38948 5800 40448 5828
rect 34440 5732 36952 5760
rect 34348 5692 34376 5720
rect 34517 5695 34575 5701
rect 34517 5692 34529 5695
rect 34348 5664 34529 5692
rect 34517 5661 34529 5664
rect 34563 5661 34575 5695
rect 34517 5655 34575 5661
rect 35437 5695 35495 5701
rect 35437 5661 35449 5695
rect 35483 5692 35495 5695
rect 35526 5692 35532 5704
rect 35483 5664 35532 5692
rect 35483 5661 35495 5664
rect 35437 5655 35495 5661
rect 35526 5652 35532 5664
rect 35584 5652 35590 5704
rect 35805 5695 35863 5701
rect 35805 5661 35817 5695
rect 35851 5661 35863 5695
rect 35805 5655 35863 5661
rect 32355 5596 34284 5624
rect 32355 5593 32367 5596
rect 32309 5587 32367 5593
rect 34330 5584 34336 5636
rect 34388 5584 34394 5636
rect 34425 5627 34483 5633
rect 34425 5593 34437 5627
rect 34471 5593 34483 5627
rect 34425 5587 34483 5593
rect 33686 5556 33692 5568
rect 31036 5528 33692 5556
rect 30929 5519 30987 5525
rect 33686 5516 33692 5528
rect 33744 5516 33750 5568
rect 33962 5516 33968 5568
rect 34020 5556 34026 5568
rect 34440 5556 34468 5587
rect 34020 5528 34468 5556
rect 34020 5516 34026 5528
rect 34698 5516 34704 5568
rect 34756 5556 34762 5568
rect 34793 5559 34851 5565
rect 34793 5556 34805 5559
rect 34756 5528 34805 5556
rect 34756 5516 34762 5528
rect 34793 5525 34805 5528
rect 34839 5525 34851 5559
rect 34793 5519 34851 5525
rect 34974 5516 34980 5568
rect 35032 5556 35038 5568
rect 35621 5559 35679 5565
rect 35621 5556 35633 5559
rect 35032 5528 35633 5556
rect 35032 5516 35038 5528
rect 35621 5525 35633 5528
rect 35667 5525 35679 5559
rect 35820 5556 35848 5655
rect 35986 5652 35992 5704
rect 36044 5652 36050 5704
rect 36081 5695 36139 5701
rect 36081 5661 36093 5695
rect 36127 5661 36139 5695
rect 36081 5655 36139 5661
rect 36096 5624 36124 5655
rect 36170 5652 36176 5704
rect 36228 5652 36234 5704
rect 36924 5701 36952 5732
rect 37274 5720 37280 5772
rect 37332 5760 37338 5772
rect 38948 5760 38976 5800
rect 37332 5732 38976 5760
rect 37332 5720 37338 5732
rect 39114 5720 39120 5772
rect 39172 5720 39178 5772
rect 36909 5695 36967 5701
rect 36909 5661 36921 5695
rect 36955 5661 36967 5695
rect 36909 5655 36967 5661
rect 37826 5652 37832 5704
rect 37884 5692 37890 5704
rect 38562 5692 38568 5704
rect 37884 5664 38568 5692
rect 37884 5652 37890 5664
rect 38562 5652 38568 5664
rect 38620 5652 38626 5704
rect 38933 5695 38991 5701
rect 38933 5661 38945 5695
rect 38979 5692 38991 5695
rect 39390 5692 39396 5704
rect 38979 5664 39396 5692
rect 38979 5661 38991 5664
rect 38933 5655 38991 5661
rect 39390 5652 39396 5664
rect 39448 5652 39454 5704
rect 39669 5695 39727 5701
rect 39669 5661 39681 5695
rect 39715 5692 39727 5695
rect 40313 5695 40371 5701
rect 40313 5692 40325 5695
rect 39715 5664 40325 5692
rect 39715 5661 39727 5664
rect 39669 5655 39727 5661
rect 40313 5661 40325 5664
rect 40359 5661 40371 5695
rect 40420 5692 40448 5800
rect 41414 5788 41420 5840
rect 41472 5828 41478 5840
rect 42981 5831 43039 5837
rect 42981 5828 42993 5831
rect 41472 5800 42993 5828
rect 41472 5788 41478 5800
rect 42981 5797 42993 5800
rect 43027 5797 43039 5831
rect 42981 5791 43039 5797
rect 41138 5720 41144 5772
rect 41196 5760 41202 5772
rect 41325 5763 41383 5769
rect 41325 5760 41337 5763
rect 41196 5732 41337 5760
rect 41196 5720 41202 5732
rect 41325 5729 41337 5732
rect 41371 5729 41383 5763
rect 41325 5723 41383 5729
rect 42610 5720 42616 5772
rect 42668 5760 42674 5772
rect 43533 5763 43591 5769
rect 43533 5760 43545 5763
rect 42668 5732 43545 5760
rect 42668 5720 42674 5732
rect 43533 5729 43545 5732
rect 43579 5729 43591 5763
rect 43533 5723 43591 5729
rect 41782 5692 41788 5704
rect 40420 5664 41788 5692
rect 40313 5655 40371 5661
rect 41782 5652 41788 5664
rect 41840 5652 41846 5704
rect 42058 5652 42064 5704
rect 42116 5652 42122 5704
rect 42889 5695 42947 5701
rect 42889 5661 42901 5695
rect 42935 5692 42947 5695
rect 42978 5692 42984 5704
rect 42935 5664 42984 5692
rect 42935 5661 42947 5664
rect 42889 5655 42947 5661
rect 42978 5652 42984 5664
rect 43036 5652 43042 5704
rect 43162 5652 43168 5704
rect 43220 5692 43226 5704
rect 43717 5695 43775 5701
rect 43717 5692 43729 5695
rect 43220 5664 43729 5692
rect 43220 5652 43226 5664
rect 43717 5661 43729 5664
rect 43763 5661 43775 5695
rect 43717 5655 43775 5661
rect 44729 5695 44787 5701
rect 44729 5661 44741 5695
rect 44775 5692 44787 5695
rect 45922 5692 45928 5704
rect 44775 5664 45928 5692
rect 44775 5661 44787 5664
rect 44729 5655 44787 5661
rect 45922 5652 45928 5664
rect 45980 5652 45986 5704
rect 46569 5695 46627 5701
rect 46569 5661 46581 5695
rect 46615 5692 46627 5695
rect 48774 5692 48780 5704
rect 46615 5664 48780 5692
rect 46615 5661 46627 5664
rect 46569 5655 46627 5661
rect 48774 5652 48780 5664
rect 48832 5652 48838 5704
rect 36262 5624 36268 5636
rect 36096 5596 36268 5624
rect 36262 5584 36268 5596
rect 36320 5584 36326 5636
rect 40862 5624 40868 5636
rect 36372 5596 40868 5624
rect 36372 5556 36400 5596
rect 40862 5584 40868 5596
rect 40920 5584 40926 5636
rect 45281 5627 45339 5633
rect 45281 5593 45293 5627
rect 45327 5624 45339 5627
rect 49786 5624 49792 5636
rect 45327 5596 49792 5624
rect 45327 5593 45339 5596
rect 45281 5587 45339 5593
rect 49786 5584 49792 5596
rect 49844 5584 49850 5636
rect 35820 5528 36400 5556
rect 35621 5519 35679 5525
rect 37826 5516 37832 5568
rect 37884 5556 37890 5568
rect 38194 5556 38200 5568
rect 37884 5528 38200 5556
rect 37884 5516 37890 5528
rect 38194 5516 38200 5528
rect 38252 5516 38258 5568
rect 39022 5516 39028 5568
rect 39080 5556 39086 5568
rect 39761 5559 39819 5565
rect 39761 5556 39773 5559
rect 39080 5528 39773 5556
rect 39080 5516 39086 5528
rect 39761 5525 39773 5528
rect 39807 5525 39819 5559
rect 39761 5519 39819 5525
rect 40494 5516 40500 5568
rect 40552 5556 40558 5568
rect 40773 5559 40831 5565
rect 40773 5556 40785 5559
rect 40552 5528 40785 5556
rect 40552 5516 40558 5528
rect 40773 5525 40785 5528
rect 40819 5525 40831 5559
rect 40773 5519 40831 5525
rect 41690 5516 41696 5568
rect 41748 5556 41754 5568
rect 42245 5559 42303 5565
rect 42245 5556 42257 5559
rect 41748 5528 42257 5556
rect 41748 5516 41754 5528
rect 42245 5525 42257 5528
rect 42291 5525 42303 5559
rect 42245 5519 42303 5525
rect 44266 5516 44272 5568
rect 44324 5516 44330 5568
rect 45925 5559 45983 5565
rect 45925 5525 45937 5559
rect 45971 5556 45983 5559
rect 46934 5556 46940 5568
rect 45971 5528 46940 5556
rect 45971 5525 45983 5528
rect 45925 5519 45983 5525
rect 46934 5516 46940 5528
rect 46992 5516 46998 5568
rect 2024 5466 77924 5488
rect 2024 5414 5794 5466
rect 5846 5414 5858 5466
rect 5910 5414 5922 5466
rect 5974 5414 5986 5466
rect 6038 5414 6050 5466
rect 6102 5414 36514 5466
rect 36566 5414 36578 5466
rect 36630 5414 36642 5466
rect 36694 5414 36706 5466
rect 36758 5414 36770 5466
rect 36822 5414 67234 5466
rect 67286 5414 67298 5466
rect 67350 5414 67362 5466
rect 67414 5414 67426 5466
rect 67478 5414 67490 5466
rect 67542 5414 77924 5466
rect 2024 5392 77924 5414
rect 8941 5355 8999 5361
rect 8941 5321 8953 5355
rect 8987 5352 8999 5355
rect 10686 5352 10692 5364
rect 8987 5324 10692 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 10778 5312 10784 5364
rect 10836 5312 10842 5364
rect 11517 5355 11575 5361
rect 11517 5321 11529 5355
rect 11563 5352 11575 5355
rect 11882 5352 11888 5364
rect 11563 5324 11888 5352
rect 11563 5321 11575 5324
rect 11517 5315 11575 5321
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 14461 5355 14519 5361
rect 14461 5321 14473 5355
rect 14507 5352 14519 5355
rect 15010 5352 15016 5364
rect 14507 5324 15016 5352
rect 14507 5321 14519 5324
rect 14461 5315 14519 5321
rect 15010 5312 15016 5324
rect 15068 5312 15074 5364
rect 15194 5312 15200 5364
rect 15252 5312 15258 5364
rect 15930 5312 15936 5364
rect 15988 5312 15994 5364
rect 18138 5312 18144 5364
rect 18196 5312 18202 5364
rect 18877 5355 18935 5361
rect 18877 5321 18889 5355
rect 18923 5352 18935 5355
rect 18966 5352 18972 5364
rect 18923 5324 18972 5352
rect 18923 5321 18935 5324
rect 18877 5315 18935 5321
rect 18966 5312 18972 5324
rect 19024 5312 19030 5364
rect 19150 5312 19156 5364
rect 19208 5352 19214 5364
rect 19208 5324 20392 5352
rect 19208 5312 19214 5324
rect 8573 5287 8631 5293
rect 8573 5253 8585 5287
rect 8619 5284 8631 5287
rect 12526 5284 12532 5296
rect 8619 5256 12532 5284
rect 8619 5253 8631 5256
rect 8573 5247 8631 5253
rect 12526 5244 12532 5256
rect 12584 5244 12590 5296
rect 12986 5244 12992 5296
rect 13044 5244 13050 5296
rect 13725 5287 13783 5293
rect 13725 5253 13737 5287
rect 13771 5284 13783 5287
rect 16206 5284 16212 5296
rect 13771 5256 16212 5284
rect 13771 5253 13783 5256
rect 13725 5247 13783 5253
rect 16206 5244 16212 5256
rect 16264 5244 16270 5296
rect 18506 5244 18512 5296
rect 18564 5284 18570 5296
rect 19245 5287 19303 5293
rect 19245 5284 19257 5287
rect 18564 5256 19257 5284
rect 18564 5244 18570 5256
rect 19245 5253 19257 5256
rect 19291 5253 19303 5287
rect 19245 5247 19303 5253
rect 20364 5228 20392 5324
rect 20530 5312 20536 5364
rect 20588 5352 20594 5364
rect 20809 5355 20867 5361
rect 20809 5352 20821 5355
rect 20588 5324 20821 5352
rect 20588 5312 20594 5324
rect 20809 5321 20821 5324
rect 20855 5321 20867 5355
rect 21542 5352 21548 5364
rect 20809 5315 20867 5321
rect 20916 5324 21548 5352
rect 20916 5284 20944 5324
rect 21542 5312 21548 5324
rect 21600 5352 21606 5364
rect 21600 5324 21685 5352
rect 21600 5312 21606 5324
rect 20656 5256 20944 5284
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5216 8079 5219
rect 9858 5216 9864 5228
rect 8067 5188 9864 5216
rect 8067 5185 8079 5188
rect 8021 5179 8079 5185
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5117 9551 5151
rect 9968 5148 9996 5179
rect 10226 5176 10232 5228
rect 10284 5176 10290 5228
rect 10410 5176 10416 5228
rect 10468 5216 10474 5228
rect 10873 5219 10931 5225
rect 10873 5216 10885 5219
rect 10468 5188 10885 5216
rect 10468 5176 10474 5188
rect 10873 5185 10885 5188
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 11606 5176 11612 5228
rect 11664 5176 11670 5228
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 12342 5216 12348 5228
rect 12299 5188 12348 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12342 5176 12348 5188
rect 12400 5176 12406 5228
rect 12621 5219 12679 5225
rect 12621 5185 12633 5219
rect 12667 5216 12679 5219
rect 15010 5216 15016 5228
rect 12667 5188 15016 5216
rect 12667 5185 12679 5188
rect 12621 5179 12679 5185
rect 12636 5148 12664 5179
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 16850 5216 16856 5228
rect 16715 5188 16856 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 17586 5176 17592 5228
rect 17644 5176 17650 5228
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 17865 5219 17923 5225
rect 17865 5216 17877 5219
rect 17736 5188 17877 5216
rect 17736 5176 17742 5188
rect 17865 5185 17877 5188
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 18969 5219 19027 5225
rect 18969 5216 18981 5219
rect 18196 5188 18981 5216
rect 18196 5176 18202 5188
rect 18969 5185 18981 5188
rect 19015 5185 19027 5219
rect 18969 5179 19027 5185
rect 20346 5176 20352 5228
rect 20404 5176 20410 5228
rect 9968 5120 12664 5148
rect 9493 5111 9551 5117
rect 9508 5080 9536 5111
rect 13170 5108 13176 5160
rect 13228 5108 13234 5160
rect 13814 5108 13820 5160
rect 13872 5108 13878 5160
rect 13906 5108 13912 5160
rect 13964 5148 13970 5160
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 13964 5120 14565 5148
rect 13964 5108 13970 5120
rect 14553 5117 14565 5120
rect 14599 5117 14611 5151
rect 14553 5111 14611 5117
rect 15286 5108 15292 5160
rect 15344 5108 15350 5160
rect 15746 5108 15752 5160
rect 15804 5148 15810 5160
rect 16298 5148 16304 5160
rect 15804 5120 16304 5148
rect 15804 5108 15810 5120
rect 16298 5108 16304 5120
rect 16356 5108 16362 5160
rect 16758 5108 16764 5160
rect 16816 5108 16822 5160
rect 18230 5108 18236 5160
rect 18288 5108 18294 5160
rect 18506 5108 18512 5160
rect 18564 5148 18570 5160
rect 20656 5148 20684 5256
rect 20990 5244 20996 5296
rect 21048 5284 21054 5296
rect 21657 5284 21685 5324
rect 21726 5312 21732 5364
rect 21784 5312 21790 5364
rect 21818 5312 21824 5364
rect 21876 5352 21882 5364
rect 23658 5352 23664 5364
rect 21876 5324 23664 5352
rect 21876 5312 21882 5324
rect 23658 5312 23664 5324
rect 23716 5312 23722 5364
rect 24026 5312 24032 5364
rect 24084 5312 24090 5364
rect 24854 5312 24860 5364
rect 24912 5352 24918 5364
rect 25041 5355 25099 5361
rect 25041 5352 25053 5355
rect 24912 5324 25053 5352
rect 24912 5312 24918 5324
rect 25041 5321 25053 5324
rect 25087 5321 25099 5355
rect 25041 5315 25099 5321
rect 26237 5355 26295 5361
rect 26237 5321 26249 5355
rect 26283 5352 26295 5355
rect 28810 5352 28816 5364
rect 26283 5324 28816 5352
rect 26283 5321 26295 5324
rect 26237 5315 26295 5321
rect 28810 5312 28816 5324
rect 28868 5312 28874 5364
rect 31846 5352 31852 5364
rect 28920 5324 31852 5352
rect 21048 5256 21404 5284
rect 21657 5256 21864 5284
rect 21048 5244 21054 5256
rect 20806 5216 20812 5228
rect 20732 5188 20812 5216
rect 20732 5157 20760 5188
rect 20806 5176 20812 5188
rect 20864 5216 20870 5228
rect 21177 5219 21235 5225
rect 21177 5216 21189 5219
rect 20864 5188 21189 5216
rect 20864 5176 20870 5188
rect 21177 5185 21189 5188
rect 21223 5185 21235 5219
rect 21177 5179 21235 5185
rect 21376 5157 21404 5256
rect 21450 5176 21456 5228
rect 21508 5216 21514 5228
rect 21836 5225 21864 5256
rect 22278 5244 22284 5296
rect 22336 5284 22342 5296
rect 22557 5287 22615 5293
rect 22557 5284 22569 5287
rect 22336 5256 22569 5284
rect 22336 5244 22342 5256
rect 22557 5253 22569 5256
rect 22603 5253 22615 5287
rect 22741 5287 22799 5293
rect 22741 5284 22753 5287
rect 22557 5247 22615 5253
rect 22664 5256 22753 5284
rect 21637 5219 21695 5225
rect 21637 5216 21649 5219
rect 21508 5188 21649 5216
rect 21508 5176 21514 5188
rect 21637 5185 21649 5188
rect 21683 5185 21695 5219
rect 21637 5179 21695 5185
rect 21821 5219 21879 5225
rect 21821 5185 21833 5219
rect 21867 5185 21879 5219
rect 22664 5216 22692 5256
rect 22741 5253 22753 5256
rect 22787 5284 22799 5287
rect 23566 5284 23572 5296
rect 22787 5256 23572 5284
rect 22787 5253 22799 5256
rect 22741 5247 22799 5253
rect 23566 5244 23572 5256
rect 23624 5244 23630 5296
rect 23842 5244 23848 5296
rect 23900 5284 23906 5296
rect 27893 5287 27951 5293
rect 27893 5284 27905 5287
rect 23900 5256 27905 5284
rect 23900 5244 23906 5256
rect 27893 5253 27905 5256
rect 27939 5253 27951 5287
rect 27893 5247 27951 5253
rect 28166 5244 28172 5296
rect 28224 5244 28230 5296
rect 24949 5219 25007 5225
rect 24949 5216 24961 5219
rect 21821 5179 21879 5185
rect 22572 5188 22692 5216
rect 22848 5188 24961 5216
rect 18564 5120 20684 5148
rect 20717 5151 20775 5157
rect 18564 5108 18570 5120
rect 20717 5117 20729 5151
rect 20763 5117 20775 5151
rect 20717 5111 20775 5117
rect 21269 5151 21327 5157
rect 21269 5117 21281 5151
rect 21315 5117 21327 5151
rect 21269 5111 21327 5117
rect 21361 5151 21419 5157
rect 21361 5117 21373 5151
rect 21407 5117 21419 5151
rect 21361 5111 21419 5117
rect 9508 5052 10364 5080
rect 9861 5015 9919 5021
rect 9861 4981 9873 5015
rect 9907 5012 9919 5015
rect 9950 5012 9956 5024
rect 9907 4984 9956 5012
rect 9907 4981 9919 4984
rect 9861 4975 9919 4981
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 10336 5012 10364 5052
rect 10410 5040 10416 5092
rect 10468 5080 10474 5092
rect 16025 5083 16083 5089
rect 16025 5080 16037 5083
rect 10468 5052 16037 5080
rect 10468 5040 10474 5052
rect 16025 5049 16037 5052
rect 16071 5049 16083 5083
rect 16025 5043 16083 5049
rect 17405 5083 17463 5089
rect 17405 5049 17417 5083
rect 17451 5080 17463 5083
rect 17451 5052 18644 5080
rect 17451 5049 17463 5052
rect 17405 5043 17463 5049
rect 12434 5012 12440 5024
rect 10336 4984 12440 5012
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 14550 4972 14556 5024
rect 14608 5012 14614 5024
rect 17586 5012 17592 5024
rect 14608 4984 17592 5012
rect 14608 4972 14614 4984
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 17957 5015 18015 5021
rect 17957 4981 17969 5015
rect 18003 5012 18015 5015
rect 18506 5012 18512 5024
rect 18003 4984 18512 5012
rect 18003 4981 18015 4984
rect 17957 4975 18015 4981
rect 18506 4972 18512 4984
rect 18564 4972 18570 5024
rect 18616 5012 18644 5052
rect 18892 5052 19104 5080
rect 18892 5012 18920 5052
rect 18616 4984 18920 5012
rect 19076 5012 19104 5052
rect 20438 5040 20444 5092
rect 20496 5080 20502 5092
rect 21284 5080 21312 5111
rect 21726 5108 21732 5160
rect 21784 5148 21790 5160
rect 21913 5151 21971 5157
rect 21913 5148 21925 5151
rect 21784 5120 21925 5148
rect 21784 5108 21790 5120
rect 21913 5117 21925 5120
rect 21959 5117 21971 5151
rect 21913 5111 21971 5117
rect 20496 5052 21312 5080
rect 20496 5040 20502 5052
rect 21818 5040 21824 5092
rect 21876 5080 21882 5092
rect 22572 5080 22600 5188
rect 21876 5052 22600 5080
rect 21876 5040 21882 5052
rect 22848 5012 22876 5188
rect 24949 5185 24961 5188
rect 24995 5185 25007 5219
rect 24949 5179 25007 5185
rect 25148 5188 25636 5216
rect 23106 5108 23112 5160
rect 23164 5148 23170 5160
rect 25148 5148 25176 5188
rect 23164 5120 25176 5148
rect 25225 5151 25283 5157
rect 23164 5108 23170 5120
rect 25225 5117 25237 5151
rect 25271 5148 25283 5151
rect 25406 5148 25412 5160
rect 25271 5120 25412 5148
rect 25271 5117 25283 5120
rect 25225 5111 25283 5117
rect 25406 5108 25412 5120
rect 25464 5108 25470 5160
rect 25608 5148 25636 5188
rect 25682 5176 25688 5228
rect 25740 5176 25746 5228
rect 26421 5219 26479 5225
rect 26421 5185 26433 5219
rect 26467 5216 26479 5219
rect 28718 5216 28724 5228
rect 26467 5188 28724 5216
rect 26467 5185 26479 5188
rect 26421 5179 26479 5185
rect 28718 5176 28724 5188
rect 28776 5176 28782 5228
rect 28920 5225 28948 5324
rect 31846 5312 31852 5324
rect 31904 5312 31910 5364
rect 32398 5352 32404 5364
rect 31956 5324 32404 5352
rect 30837 5287 30895 5293
rect 30837 5284 30849 5287
rect 29104 5256 30849 5284
rect 28905 5219 28963 5225
rect 28905 5185 28917 5219
rect 28951 5185 28963 5219
rect 28905 5179 28963 5185
rect 26878 5148 26884 5160
rect 25608 5120 26884 5148
rect 26878 5108 26884 5120
rect 26936 5108 26942 5160
rect 26970 5108 26976 5160
rect 27028 5148 27034 5160
rect 27065 5151 27123 5157
rect 27065 5148 27077 5151
rect 27028 5120 27077 5148
rect 27028 5108 27034 5120
rect 27065 5117 27077 5120
rect 27111 5117 27123 5151
rect 27617 5151 27675 5157
rect 27617 5148 27629 5151
rect 27065 5111 27123 5117
rect 27172 5120 27629 5148
rect 24118 5080 24124 5092
rect 23492 5052 24124 5080
rect 19076 4984 22876 5012
rect 23014 4972 23020 5024
rect 23072 5012 23078 5024
rect 23492 5012 23520 5052
rect 24118 5040 24124 5052
rect 24176 5040 24182 5092
rect 24302 5040 24308 5092
rect 24360 5080 24366 5092
rect 27172 5080 27200 5120
rect 27617 5117 27629 5120
rect 27663 5117 27675 5151
rect 27617 5111 27675 5117
rect 28813 5151 28871 5157
rect 28813 5117 28825 5151
rect 28859 5148 28871 5151
rect 28994 5148 29000 5160
rect 28859 5120 29000 5148
rect 28859 5117 28871 5120
rect 28813 5111 28871 5117
rect 28994 5108 29000 5120
rect 29052 5108 29058 5160
rect 24360 5052 27200 5080
rect 24360 5040 24366 5052
rect 27522 5040 27528 5092
rect 27580 5080 27586 5092
rect 29104 5080 29132 5256
rect 30837 5253 30849 5256
rect 30883 5253 30895 5287
rect 30837 5247 30895 5253
rect 29270 5176 29276 5228
rect 29328 5216 29334 5228
rect 29641 5219 29699 5225
rect 29641 5216 29653 5219
rect 29328 5188 29653 5216
rect 29328 5176 29334 5188
rect 29641 5185 29653 5188
rect 29687 5185 29699 5219
rect 29641 5179 29699 5185
rect 30374 5176 30380 5228
rect 30432 5216 30438 5228
rect 30561 5219 30619 5225
rect 30561 5216 30573 5219
rect 30432 5188 30573 5216
rect 30432 5176 30438 5188
rect 30561 5185 30573 5188
rect 30607 5185 30619 5219
rect 31956 5202 31984 5324
rect 32398 5312 32404 5324
rect 32456 5312 32462 5364
rect 32769 5355 32827 5361
rect 32769 5321 32781 5355
rect 32815 5352 32827 5355
rect 33134 5352 33140 5364
rect 32815 5324 33140 5352
rect 32815 5321 32827 5324
rect 32769 5315 32827 5321
rect 33134 5312 33140 5324
rect 33192 5312 33198 5364
rect 33686 5312 33692 5364
rect 33744 5352 33750 5364
rect 36814 5352 36820 5364
rect 33744 5324 36820 5352
rect 33744 5312 33750 5324
rect 33502 5244 33508 5296
rect 33560 5284 33566 5296
rect 33560 5256 34284 5284
rect 33560 5244 33566 5256
rect 30561 5179 30619 5185
rect 32306 5176 32312 5228
rect 32364 5216 32370 5228
rect 32861 5219 32919 5225
rect 32364 5188 32628 5216
rect 32364 5176 32370 5188
rect 29546 5108 29552 5160
rect 29604 5108 29610 5160
rect 32600 5157 32628 5188
rect 32861 5185 32873 5219
rect 32907 5216 32919 5219
rect 32907 5188 34008 5216
rect 32907 5185 32919 5188
rect 32861 5179 32919 5185
rect 30285 5151 30343 5157
rect 30285 5117 30297 5151
rect 30331 5148 30343 5151
rect 32585 5151 32643 5157
rect 30331 5120 32536 5148
rect 30331 5117 30343 5120
rect 30285 5111 30343 5117
rect 27580 5052 29132 5080
rect 27580 5040 27586 5052
rect 29362 5040 29368 5092
rect 29420 5080 29426 5092
rect 32508 5080 32536 5120
rect 32585 5117 32597 5151
rect 32631 5148 32643 5151
rect 32950 5148 32956 5160
rect 32631 5120 32956 5148
rect 32631 5117 32643 5120
rect 32585 5111 32643 5117
rect 32950 5108 32956 5120
rect 33008 5108 33014 5160
rect 33870 5108 33876 5160
rect 33928 5108 33934 5160
rect 33980 5148 34008 5188
rect 34054 5176 34060 5228
rect 34112 5176 34118 5228
rect 34256 5225 34284 5256
rect 34348 5225 34376 5324
rect 36814 5312 36820 5324
rect 36872 5312 36878 5364
rect 37461 5355 37519 5361
rect 37461 5321 37473 5355
rect 37507 5352 37519 5355
rect 39758 5352 39764 5364
rect 37507 5324 39764 5352
rect 37507 5321 37519 5324
rect 37461 5315 37519 5321
rect 39758 5312 39764 5324
rect 39816 5312 39822 5364
rect 39850 5312 39856 5364
rect 39908 5352 39914 5364
rect 41598 5352 41604 5364
rect 39908 5324 41604 5352
rect 39908 5312 39914 5324
rect 41598 5312 41604 5324
rect 41656 5312 41662 5364
rect 41785 5355 41843 5361
rect 41785 5321 41797 5355
rect 41831 5352 41843 5355
rect 42058 5352 42064 5364
rect 41831 5324 42064 5352
rect 41831 5321 41843 5324
rect 41785 5315 41843 5321
rect 42058 5312 42064 5324
rect 42116 5312 42122 5364
rect 42518 5312 42524 5364
rect 42576 5352 42582 5364
rect 42705 5355 42763 5361
rect 42705 5352 42717 5355
rect 42576 5324 42717 5352
rect 42576 5312 42582 5324
rect 42705 5321 42717 5324
rect 42751 5321 42763 5355
rect 42705 5315 42763 5321
rect 36538 5284 36544 5296
rect 34900 5256 36544 5284
rect 34241 5219 34299 5225
rect 34241 5185 34253 5219
rect 34287 5185 34299 5219
rect 34241 5179 34299 5185
rect 34333 5219 34391 5225
rect 34333 5185 34345 5219
rect 34379 5185 34391 5219
rect 34333 5179 34391 5185
rect 34425 5219 34483 5225
rect 34425 5185 34437 5219
rect 34471 5216 34483 5219
rect 34606 5216 34612 5228
rect 34471 5188 34612 5216
rect 34471 5185 34483 5188
rect 34425 5179 34483 5185
rect 34606 5176 34612 5188
rect 34664 5176 34670 5228
rect 34900 5225 34928 5256
rect 36538 5244 36544 5256
rect 36596 5244 36602 5296
rect 37734 5244 37740 5296
rect 37792 5284 37798 5296
rect 40126 5284 40132 5296
rect 37792 5256 40132 5284
rect 37792 5244 37798 5256
rect 40126 5244 40132 5256
rect 40184 5244 40190 5296
rect 42150 5244 42156 5296
rect 42208 5284 42214 5296
rect 44085 5287 44143 5293
rect 44085 5284 44097 5287
rect 42208 5256 44097 5284
rect 42208 5244 42214 5256
rect 44085 5253 44097 5256
rect 44131 5253 44143 5287
rect 44085 5247 44143 5253
rect 34885 5219 34943 5225
rect 34885 5185 34897 5219
rect 34931 5185 34943 5219
rect 34885 5179 34943 5185
rect 35158 5176 35164 5228
rect 35216 5216 35222 5228
rect 36078 5216 36084 5228
rect 35216 5188 36084 5216
rect 35216 5176 35222 5188
rect 36078 5176 36084 5188
rect 36136 5176 36142 5228
rect 36173 5219 36231 5225
rect 36173 5185 36185 5219
rect 36219 5216 36231 5219
rect 37369 5219 37427 5225
rect 37369 5216 37381 5219
rect 36219 5188 37381 5216
rect 36219 5185 36231 5188
rect 36173 5179 36231 5185
rect 37369 5185 37381 5188
rect 37415 5185 37427 5219
rect 37369 5179 37427 5185
rect 37550 5176 37556 5228
rect 37608 5216 37614 5228
rect 38841 5219 38899 5225
rect 37608 5188 38654 5216
rect 37608 5176 37614 5188
rect 35434 5148 35440 5160
rect 33980 5120 35440 5148
rect 35434 5108 35440 5120
rect 35492 5108 35498 5160
rect 35621 5151 35679 5157
rect 35621 5117 35633 5151
rect 35667 5148 35679 5151
rect 36446 5148 36452 5160
rect 35667 5120 36452 5148
rect 35667 5117 35679 5120
rect 35621 5111 35679 5117
rect 36446 5108 36452 5120
rect 36504 5108 36510 5160
rect 37660 5157 37688 5188
rect 38626 5160 38654 5188
rect 38841 5185 38853 5219
rect 38887 5216 38899 5219
rect 39669 5219 39727 5225
rect 39669 5216 39681 5219
rect 38887 5188 39681 5216
rect 38887 5185 38899 5188
rect 38841 5179 38899 5185
rect 39669 5185 39681 5188
rect 39715 5185 39727 5219
rect 39669 5179 39727 5185
rect 40494 5176 40500 5228
rect 40552 5176 40558 5228
rect 41049 5219 41107 5225
rect 41049 5185 41061 5219
rect 41095 5216 41107 5219
rect 42613 5219 42671 5225
rect 42613 5216 42625 5219
rect 41095 5188 42625 5216
rect 41095 5185 41107 5188
rect 41049 5179 41107 5185
rect 42613 5185 42625 5188
rect 42659 5185 42671 5219
rect 42613 5179 42671 5185
rect 42889 5219 42947 5225
rect 42889 5185 42901 5219
rect 42935 5216 42947 5219
rect 43070 5216 43076 5228
rect 42935 5188 43076 5216
rect 42935 5185 42947 5188
rect 42889 5179 42947 5185
rect 43070 5176 43076 5188
rect 43128 5216 43134 5228
rect 43530 5216 43536 5228
rect 43128 5188 43536 5216
rect 43128 5176 43134 5188
rect 43530 5176 43536 5188
rect 43588 5176 43594 5228
rect 44266 5176 44272 5228
rect 44324 5216 44330 5228
rect 44821 5219 44879 5225
rect 44821 5216 44833 5219
rect 44324 5188 44833 5216
rect 44324 5176 44330 5188
rect 44821 5185 44833 5188
rect 44867 5185 44879 5219
rect 44821 5179 44879 5185
rect 46934 5176 46940 5228
rect 46992 5176 46998 5228
rect 36909 5151 36967 5157
rect 36909 5117 36921 5151
rect 36955 5148 36967 5151
rect 37645 5151 37703 5157
rect 36955 5120 37596 5148
rect 36955 5117 36967 5120
rect 36909 5111 36967 5117
rect 34238 5080 34244 5092
rect 29420 5052 30696 5080
rect 32508 5052 34244 5080
rect 29420 5040 29426 5052
rect 23072 4984 23520 5012
rect 23072 4972 23078 4984
rect 23750 4972 23756 5024
rect 23808 5012 23814 5024
rect 24581 5015 24639 5021
rect 24581 5012 24593 5015
rect 23808 4984 24593 5012
rect 23808 4972 23814 4984
rect 24581 4981 24593 4984
rect 24627 4981 24639 5015
rect 24581 4975 24639 4981
rect 25406 4972 25412 5024
rect 25464 4972 25470 5024
rect 26973 5015 27031 5021
rect 26973 4981 26985 5015
rect 27019 5012 27031 5015
rect 30190 5012 30196 5024
rect 27019 4984 30196 5012
rect 27019 4981 27031 4984
rect 26973 4975 27031 4981
rect 30190 4972 30196 4984
rect 30248 5012 30254 5024
rect 30558 5012 30564 5024
rect 30248 4984 30564 5012
rect 30248 4972 30254 4984
rect 30558 4972 30564 4984
rect 30616 4972 30622 5024
rect 30668 5012 30696 5052
rect 34238 5040 34244 5052
rect 34296 5040 34302 5092
rect 34882 5040 34888 5092
rect 34940 5080 34946 5092
rect 36265 5083 36323 5089
rect 36265 5080 36277 5083
rect 34940 5052 36277 5080
rect 34940 5040 34946 5052
rect 36265 5049 36277 5052
rect 36311 5049 36323 5083
rect 36265 5043 36323 5049
rect 36538 5040 36544 5092
rect 36596 5080 36602 5092
rect 37001 5083 37059 5089
rect 37001 5080 37013 5083
rect 36596 5052 37013 5080
rect 36596 5040 36602 5052
rect 37001 5049 37013 5052
rect 37047 5049 37059 5083
rect 37568 5080 37596 5120
rect 37645 5117 37657 5151
rect 37691 5117 37703 5151
rect 37645 5111 37703 5117
rect 38289 5151 38347 5157
rect 38289 5117 38301 5151
rect 38335 5117 38347 5151
rect 38626 5120 38660 5160
rect 38289 5111 38347 5117
rect 37734 5080 37740 5092
rect 37568 5052 37740 5080
rect 37001 5043 37059 5049
rect 37734 5040 37740 5052
rect 37792 5040 37798 5092
rect 38304 5080 38332 5111
rect 38654 5108 38660 5120
rect 38712 5108 38718 5160
rect 39022 5108 39028 5160
rect 39080 5108 39086 5160
rect 40313 5151 40371 5157
rect 40313 5117 40325 5151
rect 40359 5148 40371 5151
rect 41141 5151 41199 5157
rect 41141 5148 41153 5151
rect 40359 5120 41153 5148
rect 40359 5117 40371 5120
rect 40313 5111 40371 5117
rect 41141 5117 41153 5120
rect 41187 5117 41199 5151
rect 41141 5111 41199 5117
rect 41598 5108 41604 5160
rect 41656 5148 41662 5160
rect 42058 5148 42064 5160
rect 41656 5120 42064 5148
rect 41656 5108 41662 5120
rect 42058 5108 42064 5120
rect 42116 5148 42122 5160
rect 42429 5151 42487 5157
rect 42429 5148 42441 5151
rect 42116 5120 42441 5148
rect 42116 5108 42122 5120
rect 42429 5117 42441 5120
rect 42475 5117 42487 5151
rect 42429 5111 42487 5117
rect 43993 5151 44051 5157
rect 43993 5117 44005 5151
rect 44039 5148 44051 5151
rect 44634 5148 44640 5160
rect 44039 5120 44640 5148
rect 44039 5117 44051 5120
rect 43993 5111 44051 5117
rect 44634 5108 44640 5120
rect 44692 5108 44698 5160
rect 44726 5108 44732 5160
rect 44784 5108 44790 5160
rect 45465 5151 45523 5157
rect 45465 5117 45477 5151
rect 45511 5148 45523 5151
rect 45557 5151 45615 5157
rect 45557 5148 45569 5151
rect 45511 5120 45569 5148
rect 45511 5117 45523 5120
rect 45465 5111 45523 5117
rect 45557 5117 45569 5120
rect 45603 5117 45615 5151
rect 45557 5111 45615 5117
rect 76926 5108 76932 5160
rect 76984 5148 76990 5160
rect 77481 5151 77539 5157
rect 77481 5148 77493 5151
rect 76984 5120 77493 5148
rect 76984 5108 76990 5120
rect 77481 5117 77493 5120
rect 77527 5117 77539 5151
rect 77481 5111 77539 5117
rect 41877 5083 41935 5089
rect 41877 5080 41889 5083
rect 38304 5052 38654 5080
rect 31846 5012 31852 5024
rect 30668 4984 31852 5012
rect 31846 4972 31852 4984
rect 31904 4972 31910 5024
rect 33226 4972 33232 5024
rect 33284 5012 33290 5024
rect 33321 5015 33379 5021
rect 33321 5012 33333 5015
rect 33284 4984 33333 5012
rect 33284 4972 33290 4984
rect 33321 4981 33333 4984
rect 33367 4981 33379 5015
rect 33321 4975 33379 4981
rect 34701 5015 34759 5021
rect 34701 4981 34713 5015
rect 34747 5012 34759 5015
rect 35158 5012 35164 5024
rect 34747 4984 35164 5012
rect 34747 4981 34759 4984
rect 34701 4975 34759 4981
rect 35158 4972 35164 4984
rect 35216 4972 35222 5024
rect 35437 5015 35495 5021
rect 35437 4981 35449 5015
rect 35483 5012 35495 5015
rect 37918 5012 37924 5024
rect 35483 4984 37924 5012
rect 35483 4981 35495 4984
rect 35437 4975 35495 4981
rect 37918 4972 37924 4984
rect 37976 4972 37982 5024
rect 38626 5012 38654 5052
rect 39500 5052 41889 5080
rect 39500 5012 39528 5052
rect 41877 5049 41889 5052
rect 41923 5049 41935 5083
rect 41877 5043 41935 5049
rect 42886 5040 42892 5092
rect 42944 5080 42950 5092
rect 43349 5083 43407 5089
rect 43349 5080 43361 5083
rect 42944 5052 43361 5080
rect 42944 5040 42950 5052
rect 43349 5049 43361 5052
rect 43395 5049 43407 5083
rect 43349 5043 43407 5049
rect 38626 4984 39528 5012
rect 39577 5015 39635 5021
rect 39577 4981 39589 5015
rect 39623 5012 39635 5015
rect 39942 5012 39948 5024
rect 39623 4984 39948 5012
rect 39623 4981 39635 4984
rect 39577 4975 39635 4981
rect 39942 4972 39948 4984
rect 40000 4972 40006 5024
rect 43070 4972 43076 5024
rect 43128 4972 43134 5024
rect 45830 4972 45836 5024
rect 45888 5012 45894 5024
rect 46201 5015 46259 5021
rect 46201 5012 46213 5015
rect 45888 4984 46213 5012
rect 45888 4972 45894 4984
rect 46201 4981 46213 4984
rect 46247 4981 46259 5015
rect 46201 4975 46259 4981
rect 46290 4972 46296 5024
rect 46348 4972 46354 5024
rect 76650 4972 76656 5024
rect 76708 5012 76714 5024
rect 76929 5015 76987 5021
rect 76929 5012 76941 5015
rect 76708 4984 76941 5012
rect 76708 4972 76714 4984
rect 76929 4981 76941 4984
rect 76975 4981 76987 5015
rect 76929 4975 76987 4981
rect 2024 4922 77924 4944
rect 2024 4870 5134 4922
rect 5186 4870 5198 4922
rect 5250 4870 5262 4922
rect 5314 4870 5326 4922
rect 5378 4870 5390 4922
rect 5442 4870 35854 4922
rect 35906 4870 35918 4922
rect 35970 4870 35982 4922
rect 36034 4870 36046 4922
rect 36098 4870 36110 4922
rect 36162 4870 66574 4922
rect 66626 4870 66638 4922
rect 66690 4870 66702 4922
rect 66754 4870 66766 4922
rect 66818 4870 66830 4922
rect 66882 4870 77924 4922
rect 2024 4848 77924 4870
rect 8938 4768 8944 4820
rect 8996 4768 9002 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 11054 4808 11060 4820
rect 9723 4780 11060 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 11054 4768 11060 4780
rect 11112 4768 11118 4820
rect 11885 4811 11943 4817
rect 11885 4777 11897 4811
rect 11931 4808 11943 4811
rect 11974 4808 11980 4820
rect 11931 4780 11980 4808
rect 11931 4777 11943 4780
rect 11885 4771 11943 4777
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 12618 4768 12624 4820
rect 12676 4768 12682 4820
rect 13357 4811 13415 4817
rect 13357 4777 13369 4811
rect 13403 4808 13415 4811
rect 13538 4808 13544 4820
rect 13403 4780 13544 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 14829 4811 14887 4817
rect 14829 4777 14841 4811
rect 14875 4808 14887 4811
rect 16574 4808 16580 4820
rect 14875 4780 16580 4808
rect 14875 4777 14887 4780
rect 14829 4771 14887 4777
rect 16574 4768 16580 4780
rect 16632 4768 16638 4820
rect 17034 4768 17040 4820
rect 17092 4768 17098 4820
rect 17236 4780 21864 4808
rect 8404 4712 11744 4740
rect 8404 4681 8432 4712
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4641 8447 4675
rect 8389 4635 8447 4641
rect 9125 4675 9183 4681
rect 9125 4641 9137 4675
rect 9171 4672 9183 4675
rect 9766 4672 9772 4684
rect 9171 4644 9772 4672
rect 9171 4641 9183 4644
rect 9125 4635 9183 4641
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 9950 4632 9956 4684
rect 10008 4672 10014 4684
rect 11238 4672 11244 4684
rect 10008 4644 11244 4672
rect 10008 4632 10014 4644
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4672 11391 4675
rect 11606 4672 11612 4684
rect 11379 4644 11612 4672
rect 11379 4641 11391 4644
rect 11333 4635 11391 4641
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 7374 4564 7380 4616
rect 7432 4564 7438 4616
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4604 10655 4607
rect 10686 4604 10692 4616
rect 10643 4576 10692 4604
rect 10643 4573 10655 4576
rect 10597 4567 10655 4573
rect 7668 4536 7696 4567
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 9950 4536 9956 4548
rect 7668 4508 9956 4536
rect 9950 4496 9956 4508
rect 10008 4496 10014 4548
rect 10042 4496 10048 4548
rect 10100 4496 10106 4548
rect 10413 4539 10471 4545
rect 10413 4505 10425 4539
rect 10459 4536 10471 4539
rect 11054 4536 11060 4548
rect 10459 4508 11060 4536
rect 10459 4505 10471 4508
rect 10413 4499 10471 4505
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 11716 4536 11744 4712
rect 12434 4700 12440 4752
rect 12492 4740 12498 4752
rect 13170 4740 13176 4752
rect 12492 4712 13176 4740
rect 12492 4700 12498 4712
rect 13170 4700 13176 4712
rect 13228 4700 13234 4752
rect 14182 4700 14188 4752
rect 14240 4740 14246 4752
rect 14240 4712 16436 4740
rect 14240 4700 14246 4712
rect 12069 4675 12127 4681
rect 12069 4641 12081 4675
rect 12115 4672 12127 4675
rect 12158 4672 12164 4684
rect 12115 4644 12164 4672
rect 12115 4641 12127 4644
rect 12069 4635 12127 4641
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 12805 4675 12863 4681
rect 12805 4641 12817 4675
rect 12851 4672 12863 4675
rect 14366 4672 14372 4684
rect 12851 4644 14372 4672
rect 12851 4641 12863 4644
rect 12805 4635 12863 4641
rect 14366 4632 14372 4644
rect 14424 4632 14430 4684
rect 14458 4632 14464 4684
rect 14516 4672 14522 4684
rect 16408 4681 16436 4712
rect 17236 4681 17264 4780
rect 17678 4700 17684 4752
rect 17736 4740 17742 4752
rect 17773 4743 17831 4749
rect 17773 4740 17785 4743
rect 17736 4712 17785 4740
rect 17736 4700 17742 4712
rect 17773 4709 17785 4712
rect 17819 4709 17831 4743
rect 17773 4703 17831 4709
rect 18506 4700 18512 4752
rect 18564 4700 18570 4752
rect 19242 4700 19248 4752
rect 19300 4700 19306 4752
rect 19610 4700 19616 4752
rect 19668 4740 19674 4752
rect 20438 4740 20444 4752
rect 19668 4712 20444 4740
rect 19668 4700 19674 4712
rect 20438 4700 20444 4712
rect 20496 4700 20502 4752
rect 21836 4740 21864 4780
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 22738 4808 22744 4820
rect 22152 4780 22744 4808
rect 22152 4768 22158 4780
rect 22738 4768 22744 4780
rect 22796 4768 22802 4820
rect 22922 4768 22928 4820
rect 22980 4768 22986 4820
rect 27801 4811 27859 4817
rect 23216 4780 27016 4808
rect 23216 4740 23244 4780
rect 21284 4712 21772 4740
rect 21836 4712 23244 4740
rect 23308 4712 24348 4740
rect 15197 4675 15255 4681
rect 15197 4672 15209 4675
rect 14516 4644 15209 4672
rect 14516 4632 14522 4644
rect 15197 4641 15209 4644
rect 15243 4641 15255 4675
rect 15197 4635 15255 4641
rect 15381 4675 15439 4681
rect 15381 4641 15393 4675
rect 15427 4672 15439 4675
rect 16393 4675 16451 4681
rect 15427 4644 16344 4672
rect 15427 4641 15439 4644
rect 15381 4635 15439 4641
rect 13446 4564 13452 4616
rect 13504 4564 13510 4616
rect 13538 4564 13544 4616
rect 13596 4604 13602 4616
rect 14185 4607 14243 4613
rect 14185 4604 14197 4607
rect 13596 4576 14197 4604
rect 13596 4564 13602 4576
rect 14185 4573 14197 4576
rect 14231 4573 14243 4607
rect 14185 4567 14243 4573
rect 15102 4564 15108 4616
rect 15160 4564 15166 4616
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4604 15347 4607
rect 15654 4604 15660 4616
rect 15335 4576 15660 4604
rect 15335 4573 15347 4576
rect 15289 4567 15347 4573
rect 15654 4564 15660 4576
rect 15712 4564 15718 4616
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4604 15807 4607
rect 15838 4604 15844 4616
rect 15795 4576 15844 4604
rect 15795 4573 15807 4576
rect 15749 4567 15807 4573
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 16316 4604 16344 4644
rect 16393 4641 16405 4675
rect 16439 4641 16451 4675
rect 16393 4635 16451 4641
rect 17221 4675 17279 4681
rect 17221 4641 17233 4675
rect 17267 4641 17279 4675
rect 17221 4635 17279 4641
rect 17865 4675 17923 4681
rect 17865 4641 17877 4675
rect 17911 4672 17923 4675
rect 20717 4675 20775 4681
rect 20717 4672 20729 4675
rect 17911 4644 20729 4672
rect 17911 4641 17923 4644
rect 17865 4635 17923 4641
rect 20717 4641 20729 4644
rect 20763 4641 20775 4675
rect 20717 4635 20775 4641
rect 18598 4604 18604 4616
rect 16316 4576 18604 4604
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 18690 4564 18696 4616
rect 18748 4564 18754 4616
rect 19426 4564 19432 4616
rect 19484 4564 19490 4616
rect 19610 4564 19616 4616
rect 19668 4604 19674 4616
rect 19978 4604 19984 4616
rect 19668 4576 19984 4604
rect 19668 4564 19674 4576
rect 19978 4564 19984 4576
rect 20036 4604 20042 4616
rect 20349 4607 20407 4613
rect 20349 4604 20361 4607
rect 20036 4576 20361 4604
rect 20036 4564 20042 4576
rect 20349 4573 20361 4576
rect 20395 4573 20407 4607
rect 20349 4567 20407 4573
rect 20625 4607 20683 4613
rect 20625 4573 20637 4607
rect 20671 4604 20683 4607
rect 21174 4604 21180 4616
rect 20671 4576 21180 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 21174 4564 21180 4576
rect 21232 4564 21238 4616
rect 21284 4604 21312 4712
rect 21361 4675 21419 4681
rect 21361 4641 21373 4675
rect 21407 4672 21419 4675
rect 21744 4672 21772 4712
rect 23014 4672 23020 4684
rect 21407 4644 21680 4672
rect 21744 4644 23020 4672
rect 21407 4641 21419 4644
rect 21361 4635 21419 4641
rect 21453 4607 21511 4613
rect 21453 4604 21465 4607
rect 21284 4576 21465 4604
rect 21453 4573 21465 4576
rect 21499 4573 21511 4607
rect 21652 4604 21680 4644
rect 23014 4632 23020 4644
rect 23072 4632 23078 4684
rect 23308 4672 23336 4712
rect 23124 4644 23336 4672
rect 23569 4675 23627 4681
rect 22094 4604 22100 4616
rect 21652 4576 22100 4604
rect 21453 4567 21511 4573
rect 22094 4564 22100 4576
rect 22152 4564 22158 4616
rect 22278 4564 22284 4616
rect 22336 4564 22342 4616
rect 14274 4536 14280 4548
rect 11716 4508 14280 4536
rect 14274 4496 14280 4508
rect 14332 4496 14338 4548
rect 20254 4536 20260 4548
rect 15488 4508 20260 4536
rect 6822 4428 6828 4480
rect 6880 4428 6886 4480
rect 8205 4471 8263 4477
rect 8205 4437 8217 4471
rect 8251 4468 8263 4471
rect 9398 4468 9404 4480
rect 8251 4440 9404 4468
rect 8251 4437 8263 4440
rect 8205 4431 8263 4437
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 11146 4428 11152 4480
rect 11204 4428 11210 4480
rect 11422 4428 11428 4480
rect 11480 4468 11486 4480
rect 12802 4468 12808 4480
rect 11480 4440 12808 4468
rect 11480 4428 11486 4440
rect 12802 4428 12808 4440
rect 12860 4428 12866 4480
rect 14093 4471 14151 4477
rect 14093 4437 14105 4471
rect 14139 4468 14151 4471
rect 15488 4468 15516 4508
rect 20254 4496 20260 4508
rect 20312 4496 20318 4548
rect 22833 4539 22891 4545
rect 22833 4505 22845 4539
rect 22879 4536 22891 4539
rect 23124 4536 23152 4644
rect 23569 4641 23581 4675
rect 23615 4672 23627 4675
rect 24118 4672 24124 4684
rect 23615 4644 24124 4672
rect 23615 4641 23627 4644
rect 23569 4635 23627 4641
rect 24118 4632 24124 4644
rect 24176 4632 24182 4684
rect 22879 4508 23152 4536
rect 23293 4539 23351 4545
rect 22879 4505 22891 4508
rect 22833 4499 22891 4505
rect 23293 4505 23305 4539
rect 23339 4536 23351 4539
rect 24320 4536 24348 4712
rect 24394 4700 24400 4752
rect 24452 4740 24458 4752
rect 24452 4712 24808 4740
rect 24452 4700 24458 4712
rect 24673 4675 24731 4681
rect 24673 4641 24685 4675
rect 24719 4641 24731 4675
rect 24780 4672 24808 4712
rect 25406 4700 25412 4752
rect 25464 4740 25470 4752
rect 26602 4740 26608 4752
rect 25464 4712 26608 4740
rect 25464 4700 25470 4712
rect 26602 4700 26608 4712
rect 26660 4700 26666 4752
rect 25501 4675 25559 4681
rect 25501 4672 25513 4675
rect 24780 4644 25513 4672
rect 24673 4635 24731 4641
rect 25501 4641 25513 4644
rect 25547 4641 25559 4675
rect 26988 4672 27016 4780
rect 27801 4777 27813 4811
rect 27847 4808 27859 4811
rect 29822 4808 29828 4820
rect 27847 4780 29828 4808
rect 27847 4777 27859 4780
rect 27801 4771 27859 4777
rect 29822 4768 29828 4780
rect 29880 4768 29886 4820
rect 31294 4768 31300 4820
rect 31352 4808 31358 4820
rect 31389 4811 31447 4817
rect 31389 4808 31401 4811
rect 31352 4780 31401 4808
rect 31352 4768 31358 4780
rect 31389 4777 31401 4780
rect 31435 4777 31447 4811
rect 31389 4771 31447 4777
rect 31570 4768 31576 4820
rect 31628 4808 31634 4820
rect 32766 4808 32772 4820
rect 31628 4780 32772 4808
rect 31628 4768 31634 4780
rect 32766 4768 32772 4780
rect 32824 4768 32830 4820
rect 33778 4768 33784 4820
rect 33836 4808 33842 4820
rect 36078 4808 36084 4820
rect 33836 4780 36084 4808
rect 33836 4768 33842 4780
rect 36078 4768 36084 4780
rect 36136 4768 36142 4820
rect 36173 4811 36231 4817
rect 36173 4777 36185 4811
rect 36219 4808 36231 4811
rect 36262 4808 36268 4820
rect 36219 4780 36268 4808
rect 36219 4777 36231 4780
rect 36173 4771 36231 4777
rect 36262 4768 36268 4780
rect 36320 4768 36326 4820
rect 36446 4768 36452 4820
rect 36504 4808 36510 4820
rect 37458 4808 37464 4820
rect 36504 4780 37464 4808
rect 36504 4768 36510 4780
rect 37458 4768 37464 4780
rect 37516 4768 37522 4820
rect 37918 4768 37924 4820
rect 37976 4808 37982 4820
rect 38086 4811 38144 4817
rect 38086 4808 38098 4811
rect 37976 4780 38098 4808
rect 37976 4768 37982 4780
rect 38086 4777 38098 4780
rect 38132 4777 38144 4811
rect 38086 4771 38144 4777
rect 44729 4811 44787 4817
rect 44729 4777 44741 4811
rect 44775 4808 44787 4811
rect 47026 4808 47032 4820
rect 44775 4780 47032 4808
rect 44775 4777 44787 4780
rect 44729 4771 44787 4777
rect 47026 4768 47032 4780
rect 47084 4768 47090 4820
rect 76926 4768 76932 4820
rect 76984 4768 76990 4820
rect 27065 4743 27123 4749
rect 27065 4709 27077 4743
rect 27111 4740 27123 4743
rect 29549 4743 29607 4749
rect 27111 4712 29408 4740
rect 27111 4709 27123 4712
rect 27065 4703 27123 4709
rect 28258 4672 28264 4684
rect 26988 4644 28264 4672
rect 25501 4635 25559 4641
rect 24688 4604 24716 4635
rect 28258 4632 28264 4644
rect 28316 4632 28322 4684
rect 28350 4632 28356 4684
rect 28408 4632 28414 4684
rect 28445 4675 28503 4681
rect 28445 4641 28457 4675
rect 28491 4641 28503 4675
rect 28445 4635 28503 4641
rect 24762 4604 24768 4616
rect 24688 4576 24768 4604
rect 24762 4564 24768 4576
rect 24820 4564 24826 4616
rect 25133 4607 25191 4613
rect 25133 4573 25145 4607
rect 25179 4604 25191 4607
rect 25222 4604 25228 4616
rect 25179 4576 25228 4604
rect 25179 4573 25191 4576
rect 25133 4567 25191 4573
rect 25222 4564 25228 4576
rect 25280 4564 25286 4616
rect 25961 4607 26019 4613
rect 25961 4573 25973 4607
rect 26007 4573 26019 4607
rect 25961 4567 26019 4573
rect 25976 4536 26004 4567
rect 26510 4564 26516 4616
rect 26568 4564 26574 4616
rect 27249 4607 27307 4613
rect 27249 4573 27261 4607
rect 27295 4604 27307 4607
rect 27522 4604 27528 4616
rect 27295 4576 27528 4604
rect 27295 4573 27307 4576
rect 27249 4567 27307 4573
rect 27522 4564 27528 4576
rect 27580 4564 27586 4616
rect 27614 4564 27620 4616
rect 27672 4604 27678 4616
rect 28460 4604 28488 4635
rect 28902 4632 28908 4684
rect 28960 4632 28966 4684
rect 29086 4632 29092 4684
rect 29144 4672 29150 4684
rect 29270 4672 29276 4684
rect 29144 4644 29276 4672
rect 29144 4632 29150 4644
rect 29270 4632 29276 4644
rect 29328 4632 29334 4684
rect 27672 4576 28488 4604
rect 29380 4604 29408 4712
rect 29549 4709 29561 4743
rect 29595 4740 29607 4743
rect 29595 4712 31616 4740
rect 29595 4709 29607 4712
rect 29549 4703 29607 4709
rect 29733 4675 29791 4681
rect 29733 4641 29745 4675
rect 29779 4672 29791 4675
rect 30745 4675 30803 4681
rect 29779 4644 30696 4672
rect 29779 4641 29791 4644
rect 29733 4635 29791 4641
rect 30466 4604 30472 4616
rect 29380 4576 30472 4604
rect 27672 4564 27678 4576
rect 30466 4564 30472 4576
rect 30524 4564 30530 4616
rect 30668 4604 30696 4644
rect 30745 4641 30757 4675
rect 30791 4672 30803 4675
rect 30834 4672 30840 4684
rect 30791 4644 30840 4672
rect 30791 4641 30803 4644
rect 30745 4635 30803 4641
rect 30834 4632 30840 4644
rect 30892 4632 30898 4684
rect 30668 4576 31064 4604
rect 28810 4536 28816 4548
rect 23339 4508 24256 4536
rect 24320 4508 25912 4536
rect 25976 4508 28816 4536
rect 23339 4505 23351 4508
rect 23293 4499 23351 4505
rect 14139 4440 15516 4468
rect 15565 4471 15623 4477
rect 14139 4437 14151 4440
rect 14093 4431 14151 4437
rect 15565 4437 15577 4471
rect 15611 4468 15623 4471
rect 16114 4468 16120 4480
rect 15611 4440 16120 4468
rect 15611 4437 15623 4440
rect 15565 4431 15623 4437
rect 16114 4428 16120 4440
rect 16172 4428 16178 4480
rect 16298 4428 16304 4480
rect 16356 4428 16362 4480
rect 16666 4428 16672 4480
rect 16724 4468 16730 4480
rect 19518 4468 19524 4480
rect 16724 4440 19524 4468
rect 16724 4428 16730 4440
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 19978 4428 19984 4480
rect 20036 4428 20042 4480
rect 22094 4428 22100 4480
rect 22152 4428 22158 4480
rect 23385 4471 23443 4477
rect 23385 4437 23397 4471
rect 23431 4468 23443 4471
rect 23658 4468 23664 4480
rect 23431 4440 23664 4468
rect 23431 4437 23443 4440
rect 23385 4431 23443 4437
rect 23658 4428 23664 4440
rect 23716 4428 23722 4480
rect 24228 4468 24256 4508
rect 25406 4468 25412 4480
rect 24228 4440 25412 4468
rect 25406 4428 25412 4440
rect 25464 4428 25470 4480
rect 25884 4468 25912 4508
rect 28810 4496 28816 4508
rect 28868 4496 28874 4548
rect 27062 4468 27068 4480
rect 25884 4440 27068 4468
rect 27062 4428 27068 4440
rect 27120 4428 27126 4480
rect 27893 4471 27951 4477
rect 27893 4437 27905 4471
rect 27939 4468 27951 4471
rect 28074 4468 28080 4480
rect 27939 4440 28080 4468
rect 27939 4437 27951 4440
rect 27893 4431 27951 4437
rect 28074 4428 28080 4440
rect 28132 4428 28138 4480
rect 28261 4471 28319 4477
rect 28261 4437 28273 4471
rect 28307 4468 28319 4471
rect 28442 4468 28448 4480
rect 28307 4440 28448 4468
rect 28307 4437 28319 4440
rect 28261 4431 28319 4437
rect 28442 4428 28448 4440
rect 28500 4428 28506 4480
rect 30282 4428 30288 4480
rect 30340 4428 30346 4480
rect 31036 4468 31064 4576
rect 31202 4564 31208 4616
rect 31260 4604 31266 4616
rect 31297 4607 31355 4613
rect 31297 4604 31309 4607
rect 31260 4576 31309 4604
rect 31260 4564 31266 4576
rect 31297 4573 31309 4576
rect 31343 4573 31355 4607
rect 31588 4604 31616 4712
rect 31662 4700 31668 4752
rect 31720 4740 31726 4752
rect 33321 4743 33379 4749
rect 33321 4740 33333 4743
rect 31720 4712 33333 4740
rect 31720 4700 31726 4712
rect 33321 4709 33333 4712
rect 33367 4709 33379 4743
rect 34974 4740 34980 4752
rect 33321 4703 33379 4709
rect 33980 4712 34980 4740
rect 31846 4632 31852 4684
rect 31904 4632 31910 4684
rect 32033 4675 32091 4681
rect 32033 4641 32045 4675
rect 32079 4672 32091 4675
rect 32214 4672 32220 4684
rect 32079 4644 32220 4672
rect 32079 4641 32091 4644
rect 32033 4635 32091 4641
rect 32214 4632 32220 4644
rect 32272 4632 32278 4684
rect 32950 4632 32956 4684
rect 33008 4632 33014 4684
rect 33980 4681 34008 4712
rect 34974 4700 34980 4712
rect 35032 4700 35038 4752
rect 40589 4743 40647 4749
rect 40589 4709 40601 4743
rect 40635 4740 40647 4743
rect 41322 4740 41328 4752
rect 40635 4712 41328 4740
rect 40635 4709 40647 4712
rect 40589 4703 40647 4709
rect 41322 4700 41328 4712
rect 41380 4700 41386 4752
rect 43070 4740 43076 4752
rect 41524 4712 43076 4740
rect 33965 4675 34023 4681
rect 33965 4641 33977 4675
rect 34011 4641 34023 4675
rect 33965 4635 34023 4641
rect 34882 4632 34888 4684
rect 34940 4632 34946 4684
rect 36817 4675 36875 4681
rect 36817 4641 36829 4675
rect 36863 4672 36875 4675
rect 36906 4672 36912 4684
rect 36863 4644 36912 4672
rect 36863 4641 36875 4644
rect 36817 4635 36875 4641
rect 36906 4632 36912 4644
rect 36964 4632 36970 4684
rect 37461 4675 37519 4681
rect 37461 4641 37473 4675
rect 37507 4672 37519 4675
rect 37507 4644 39804 4672
rect 37507 4641 37519 4644
rect 37461 4635 37519 4641
rect 34149 4607 34207 4613
rect 31588 4576 34100 4604
rect 31297 4567 31355 4573
rect 31570 4496 31576 4548
rect 31628 4536 31634 4548
rect 31757 4539 31815 4545
rect 31757 4536 31769 4539
rect 31628 4508 31769 4536
rect 31628 4496 31634 4508
rect 31757 4505 31769 4508
rect 31803 4505 31815 4539
rect 32401 4539 32459 4545
rect 32401 4536 32413 4539
rect 31757 4499 31815 4505
rect 31864 4508 32413 4536
rect 31864 4468 31892 4508
rect 32401 4505 32413 4508
rect 32447 4505 32459 4539
rect 34072 4536 34100 4576
rect 34149 4573 34161 4607
rect 34195 4604 34207 4607
rect 34606 4604 34612 4616
rect 34195 4576 34612 4604
rect 34195 4573 34207 4576
rect 34149 4567 34207 4573
rect 34606 4564 34612 4576
rect 34664 4564 34670 4616
rect 34701 4607 34759 4613
rect 34701 4573 34713 4607
rect 34747 4604 34759 4607
rect 34747 4576 37688 4604
rect 34747 4573 34759 4576
rect 34701 4567 34759 4573
rect 36078 4536 36084 4548
rect 34072 4508 36084 4536
rect 32401 4499 32459 4505
rect 36078 4496 36084 4508
rect 36136 4496 36142 4548
rect 37660 4536 37688 4576
rect 37734 4564 37740 4616
rect 37792 4564 37798 4616
rect 37826 4564 37832 4616
rect 37884 4564 37890 4616
rect 39776 4604 39804 4644
rect 39850 4632 39856 4684
rect 39908 4632 39914 4684
rect 39942 4632 39948 4684
rect 40000 4632 40006 4684
rect 41524 4681 41552 4712
rect 43070 4700 43076 4712
rect 43128 4700 43134 4752
rect 41509 4675 41567 4681
rect 41509 4641 41521 4675
rect 41555 4641 41567 4675
rect 41509 4635 41567 4641
rect 41708 4644 43116 4672
rect 39776 4600 41644 4604
rect 41708 4600 41736 4644
rect 43088 4616 43116 4644
rect 43346 4632 43352 4684
rect 43404 4672 43410 4684
rect 43441 4675 43499 4681
rect 43441 4672 43453 4675
rect 43404 4644 43453 4672
rect 43404 4632 43410 4644
rect 43441 4641 43453 4644
rect 43487 4641 43499 4675
rect 43441 4635 43499 4641
rect 44082 4632 44088 4684
rect 44140 4672 44146 4684
rect 45097 4675 45155 4681
rect 45097 4672 45109 4675
rect 44140 4644 45109 4672
rect 44140 4632 44146 4644
rect 45097 4641 45109 4644
rect 45143 4641 45155 4675
rect 45097 4635 45155 4641
rect 45186 4632 45192 4684
rect 45244 4672 45250 4684
rect 45649 4675 45707 4681
rect 45649 4672 45661 4675
rect 45244 4644 45661 4672
rect 45244 4632 45250 4644
rect 45649 4641 45661 4644
rect 45695 4641 45707 4675
rect 45649 4635 45707 4641
rect 46569 4675 46627 4681
rect 46569 4641 46581 4675
rect 46615 4672 46627 4675
rect 47210 4672 47216 4684
rect 46615 4644 47216 4672
rect 46615 4641 46627 4644
rect 46569 4635 46627 4641
rect 47210 4632 47216 4644
rect 47268 4632 47274 4684
rect 47305 4675 47363 4681
rect 47305 4641 47317 4675
rect 47351 4672 47363 4675
rect 48133 4675 48191 4681
rect 48133 4672 48145 4675
rect 47351 4644 48145 4672
rect 47351 4641 47363 4644
rect 47305 4635 47363 4641
rect 48133 4641 48145 4644
rect 48179 4641 48191 4675
rect 48133 4635 48191 4641
rect 39776 4576 41736 4600
rect 41616 4572 41736 4576
rect 41782 4564 41788 4616
rect 41840 4564 41846 4616
rect 42061 4607 42119 4613
rect 42061 4573 42073 4607
rect 42107 4604 42119 4607
rect 42610 4604 42616 4616
rect 42107 4576 42616 4604
rect 42107 4573 42119 4576
rect 42061 4567 42119 4573
rect 42610 4564 42616 4576
rect 42668 4564 42674 4616
rect 42797 4607 42855 4613
rect 42797 4573 42809 4607
rect 42843 4573 42855 4607
rect 42797 4567 42855 4573
rect 38378 4536 38384 4548
rect 37660 4508 38384 4536
rect 38378 4496 38384 4508
rect 38436 4496 38442 4548
rect 39482 4536 39488 4548
rect 39330 4508 39488 4536
rect 31036 4440 31892 4468
rect 32122 4428 32128 4480
rect 32180 4468 32186 4480
rect 33229 4471 33287 4477
rect 33229 4468 33241 4471
rect 32180 4440 33241 4468
rect 32180 4428 32186 4440
rect 33229 4437 33241 4440
rect 33275 4468 33287 4471
rect 33778 4468 33784 4480
rect 33275 4440 33784 4468
rect 33275 4437 33287 4440
rect 33229 4431 33287 4437
rect 33778 4428 33784 4440
rect 33836 4428 33842 4480
rect 35434 4428 35440 4480
rect 35492 4428 35498 4480
rect 37550 4428 37556 4480
rect 37608 4468 37614 4480
rect 39408 4468 39436 4508
rect 39482 4496 39488 4508
rect 39540 4536 39546 4548
rect 40034 4536 40040 4548
rect 39540 4508 40040 4536
rect 39540 4496 39546 4508
rect 40034 4496 40040 4508
rect 40092 4496 40098 4548
rect 40126 4496 40132 4548
rect 40184 4536 40190 4548
rect 40865 4539 40923 4545
rect 40865 4536 40877 4539
rect 40184 4508 40877 4536
rect 40184 4496 40190 4508
rect 40865 4505 40877 4508
rect 40911 4505 40923 4539
rect 40865 4499 40923 4505
rect 40954 4496 40960 4548
rect 41012 4536 41018 4548
rect 42812 4536 42840 4567
rect 43070 4564 43076 4616
rect 43128 4564 43134 4616
rect 43993 4607 44051 4613
rect 43993 4573 44005 4607
rect 44039 4604 44051 4607
rect 44039 4576 44128 4604
rect 44039 4573 44051 4576
rect 43993 4567 44051 4573
rect 41012 4508 42840 4536
rect 44100 4536 44128 4576
rect 44174 4564 44180 4616
rect 44232 4564 44238 4616
rect 46753 4607 46811 4613
rect 46753 4573 46765 4607
rect 46799 4604 46811 4607
rect 46799 4576 47992 4604
rect 46799 4573 46811 4576
rect 46753 4567 46811 4573
rect 45462 4536 45468 4548
rect 44100 4508 45468 4536
rect 41012 4496 41018 4508
rect 45462 4496 45468 4508
rect 45520 4496 45526 4548
rect 45646 4496 45652 4548
rect 45704 4536 45710 4548
rect 47397 4539 47455 4545
rect 47397 4536 47409 4539
rect 45704 4508 47409 4536
rect 45704 4496 45710 4508
rect 47397 4505 47409 4508
rect 47443 4505 47455 4539
rect 47964 4536 47992 4576
rect 48038 4564 48044 4616
rect 48096 4564 48102 4616
rect 48866 4564 48872 4616
rect 48924 4564 48930 4616
rect 77570 4564 77576 4616
rect 77628 4564 77634 4616
rect 49970 4536 49976 4548
rect 47964 4508 49976 4536
rect 47397 4499 47455 4505
rect 49970 4496 49976 4508
rect 50028 4496 50034 4548
rect 37608 4440 39436 4468
rect 41601 4471 41659 4477
rect 37608 4428 37614 4440
rect 41601 4437 41613 4471
rect 41647 4468 41659 4471
rect 42242 4468 42248 4480
rect 41647 4440 42248 4468
rect 41647 4437 41659 4440
rect 41601 4431 41659 4437
rect 42242 4428 42248 4440
rect 42300 4428 42306 4480
rect 42613 4471 42671 4477
rect 42613 4437 42625 4471
rect 42659 4468 42671 4471
rect 43254 4468 43260 4480
rect 42659 4440 43260 4468
rect 42659 4437 42671 4440
rect 42613 4431 42671 4437
rect 43254 4428 43260 4440
rect 43312 4428 43318 4480
rect 43346 4428 43352 4480
rect 43404 4428 43410 4480
rect 45554 4428 45560 4480
rect 45612 4468 45618 4480
rect 45925 4471 45983 4477
rect 45925 4468 45937 4471
rect 45612 4440 45937 4468
rect 45612 4428 45618 4440
rect 45925 4437 45937 4440
rect 45971 4437 45983 4471
rect 45925 4431 45983 4437
rect 48314 4428 48320 4480
rect 48372 4468 48378 4480
rect 48777 4471 48835 4477
rect 48777 4468 48789 4471
rect 48372 4440 48789 4468
rect 48372 4428 48378 4440
rect 48777 4437 48789 4440
rect 48823 4437 48835 4471
rect 48777 4431 48835 4437
rect 49513 4471 49571 4477
rect 49513 4437 49525 4471
rect 49559 4468 49571 4471
rect 50522 4468 50528 4480
rect 49559 4440 50528 4468
rect 49559 4437 49571 4440
rect 49513 4431 49571 4437
rect 50522 4428 50528 4440
rect 50580 4428 50586 4480
rect 2024 4378 77924 4400
rect 2024 4326 5794 4378
rect 5846 4326 5858 4378
rect 5910 4326 5922 4378
rect 5974 4326 5986 4378
rect 6038 4326 6050 4378
rect 6102 4326 36514 4378
rect 36566 4326 36578 4378
rect 36630 4326 36642 4378
rect 36694 4326 36706 4378
rect 36758 4326 36770 4378
rect 36822 4326 67234 4378
rect 67286 4326 67298 4378
rect 67350 4326 67362 4378
rect 67414 4326 67426 4378
rect 67478 4326 67490 4378
rect 67542 4326 77924 4378
rect 2024 4304 77924 4326
rect 7374 4224 7380 4276
rect 7432 4264 7438 4276
rect 9766 4264 9772 4276
rect 7432 4236 9772 4264
rect 7432 4224 7438 4236
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 11238 4264 11244 4276
rect 10008 4236 11244 4264
rect 10008 4224 10014 4236
rect 11238 4224 11244 4236
rect 11296 4224 11302 4276
rect 13446 4224 13452 4276
rect 13504 4264 13510 4276
rect 14458 4264 14464 4276
rect 13504 4236 14464 4264
rect 13504 4224 13510 4236
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 15102 4224 15108 4276
rect 15160 4264 15166 4276
rect 16666 4264 16672 4276
rect 15160 4236 16672 4264
rect 15160 4224 15166 4236
rect 16666 4224 16672 4236
rect 16724 4224 16730 4276
rect 19886 4224 19892 4276
rect 19944 4224 19950 4276
rect 26418 4264 26424 4276
rect 25884 4236 26424 4264
rect 25884 4208 25912 4236
rect 26418 4224 26424 4236
rect 26476 4224 26482 4276
rect 26513 4267 26571 4273
rect 26513 4233 26525 4267
rect 26559 4264 26571 4267
rect 26694 4264 26700 4276
rect 26559 4236 26700 4264
rect 26559 4233 26571 4236
rect 26513 4227 26571 4233
rect 26694 4224 26700 4236
rect 26752 4224 26758 4276
rect 28810 4224 28816 4276
rect 28868 4264 28874 4276
rect 30650 4264 30656 4276
rect 28868 4236 30656 4264
rect 28868 4224 28874 4236
rect 30650 4224 30656 4236
rect 30708 4224 30714 4276
rect 31110 4224 31116 4276
rect 31168 4264 31174 4276
rect 32214 4264 32220 4276
rect 31168 4236 32220 4264
rect 31168 4224 31174 4236
rect 32214 4224 32220 4236
rect 32272 4224 32278 4276
rect 32490 4224 32496 4276
rect 32548 4264 32554 4276
rect 32950 4264 32956 4276
rect 32548 4236 32956 4264
rect 32548 4224 32554 4236
rect 32950 4224 32956 4236
rect 33008 4224 33014 4276
rect 34054 4224 34060 4276
rect 34112 4264 34118 4276
rect 38197 4267 38255 4273
rect 38197 4264 38209 4267
rect 34112 4236 38209 4264
rect 34112 4224 34118 4236
rect 38197 4233 38209 4236
rect 38243 4233 38255 4267
rect 38197 4227 38255 4233
rect 40221 4267 40279 4273
rect 40221 4233 40233 4267
rect 40267 4264 40279 4267
rect 40954 4264 40960 4276
rect 40267 4236 40960 4264
rect 40267 4233 40279 4236
rect 40221 4227 40279 4233
rect 40954 4224 40960 4236
rect 41012 4224 41018 4276
rect 41322 4224 41328 4276
rect 41380 4264 41386 4276
rect 44174 4264 44180 4276
rect 41380 4236 44180 4264
rect 41380 4224 41386 4236
rect 44174 4224 44180 4236
rect 44232 4224 44238 4276
rect 6362 4156 6368 4208
rect 6420 4196 6426 4208
rect 6914 4196 6920 4208
rect 6420 4168 6920 4196
rect 6420 4156 6426 4168
rect 6914 4156 6920 4168
rect 6972 4156 6978 4208
rect 7469 4199 7527 4205
rect 7469 4165 7481 4199
rect 7515 4196 7527 4199
rect 10226 4196 10232 4208
rect 7515 4168 10232 4196
rect 7515 4165 7527 4168
rect 7469 4159 7527 4165
rect 10226 4156 10232 4168
rect 10284 4156 10290 4208
rect 16758 4196 16764 4208
rect 10796 4168 16764 4196
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 6052 4100 6745 4128
rect 6052 4088 6058 4100
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4128 7895 4131
rect 9309 4131 9367 4137
rect 7883 4100 8800 4128
rect 7883 4097 7895 4100
rect 7837 4091 7895 4097
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 8570 4060 8576 4072
rect 8067 4032 8576 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 8772 4069 8800 4100
rect 9309 4097 9321 4131
rect 9355 4128 9367 4131
rect 10318 4128 10324 4140
rect 9355 4100 10324 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 10796 4137 10824 4168
rect 16758 4156 16764 4168
rect 16816 4156 16822 4208
rect 16868 4168 17356 4196
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 12437 4131 12495 4137
rect 12437 4128 12449 4131
rect 11204 4100 12449 4128
rect 11204 4088 11210 4100
rect 12437 4097 12449 4100
rect 12483 4097 12495 4131
rect 12437 4091 12495 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 12618 4128 12624 4140
rect 12575 4100 12624 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4128 13415 4131
rect 13722 4128 13728 4140
rect 13403 4100 13728 4128
rect 13403 4097 13415 4100
rect 13357 4091 13415 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14642 4088 14648 4140
rect 14700 4128 14706 4140
rect 14700 4100 14780 4128
rect 14700 4088 14706 4100
rect 8757 4063 8815 4069
rect 8757 4029 8769 4063
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4060 9551 4063
rect 10134 4060 10140 4072
rect 9539 4032 10140 4060
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 4890 3952 4896 4004
rect 4948 3992 4954 4004
rect 8110 3992 8116 4004
rect 4948 3964 8116 3992
rect 4948 3952 4954 3964
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 8772 3992 8800 4023
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 10410 4060 10416 4072
rect 10275 4032 10416 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 10870 4020 10876 4072
rect 10928 4020 10934 4072
rect 11517 4063 11575 4069
rect 11517 4029 11529 4063
rect 11563 4060 11575 4063
rect 11606 4060 11612 4072
rect 11563 4032 11612 4060
rect 11563 4029 11575 4032
rect 11517 4023 11575 4029
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 11698 4020 11704 4072
rect 11756 4020 11762 4072
rect 11882 4020 11888 4072
rect 11940 4060 11946 4072
rect 12713 4063 12771 4069
rect 12713 4060 12725 4063
rect 11940 4032 12725 4060
rect 11940 4020 11946 4032
rect 12713 4029 12725 4032
rect 12759 4029 12771 4063
rect 12713 4023 12771 4029
rect 14369 4063 14427 4069
rect 14369 4029 14381 4063
rect 14415 4060 14427 4063
rect 14415 4032 14688 4060
rect 14415 4029 14427 4032
rect 14369 4023 14427 4029
rect 14660 4004 14688 4032
rect 9950 3992 9956 4004
rect 8772 3964 9956 3992
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 10045 3995 10103 4001
rect 10045 3961 10057 3995
rect 10091 3992 10103 3995
rect 11974 3992 11980 4004
rect 10091 3964 11980 3992
rect 10091 3961 10103 3964
rect 10045 3955 10103 3961
rect 11974 3952 11980 3964
rect 12032 3952 12038 4004
rect 13814 3992 13820 4004
rect 12084 3964 13820 3992
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 5592 3896 6561 3924
rect 5592 3884 5598 3896
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 8573 3927 8631 3933
rect 8573 3893 8585 3927
rect 8619 3924 8631 3927
rect 12084 3924 12112 3964
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 14642 3952 14648 4004
rect 14700 3952 14706 4004
rect 14752 3992 14780 4100
rect 14826 4088 14832 4140
rect 14884 4088 14890 4140
rect 15010 4088 15016 4140
rect 15068 4088 15074 4140
rect 16390 4128 16396 4140
rect 16040 4100 16396 4128
rect 15102 4020 15108 4072
rect 15160 4060 15166 4072
rect 15197 4063 15255 4069
rect 15197 4060 15209 4063
rect 15160 4032 15209 4060
rect 15160 4020 15166 4032
rect 15197 4029 15209 4032
rect 15243 4029 15255 4063
rect 15197 4023 15255 4029
rect 15381 4063 15439 4069
rect 15381 4029 15393 4063
rect 15427 4060 15439 4063
rect 16040 4060 16068 4100
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 16574 4088 16580 4140
rect 16632 4128 16638 4140
rect 16868 4128 16896 4168
rect 16632 4100 16896 4128
rect 16632 4088 16638 4100
rect 17218 4088 17224 4140
rect 17276 4088 17282 4140
rect 17328 4128 17356 4168
rect 17586 4156 17592 4208
rect 17644 4196 17650 4208
rect 19334 4196 19340 4208
rect 17644 4168 19340 4196
rect 17644 4156 17650 4168
rect 19334 4156 19340 4168
rect 19392 4156 19398 4208
rect 19429 4199 19487 4205
rect 19429 4165 19441 4199
rect 19475 4196 19487 4199
rect 19518 4196 19524 4208
rect 19475 4168 19524 4196
rect 19475 4165 19487 4168
rect 19429 4159 19487 4165
rect 19518 4156 19524 4168
rect 19576 4156 19582 4208
rect 19812 4168 20024 4196
rect 17328 4100 18368 4128
rect 15427 4032 16068 4060
rect 16945 4063 17003 4069
rect 15427 4029 15439 4032
rect 15381 4023 15439 4029
rect 16945 4029 16957 4063
rect 16991 4060 17003 4063
rect 18230 4060 18236 4072
rect 16991 4032 18236 4060
rect 16991 4029 17003 4032
rect 16945 4023 17003 4029
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 15933 3995 15991 4001
rect 15933 3992 15945 3995
rect 14752 3964 15945 3992
rect 15933 3961 15945 3964
rect 15979 3961 15991 3995
rect 15933 3955 15991 3961
rect 18138 3952 18144 4004
rect 18196 3952 18202 4004
rect 18340 3992 18368 4100
rect 19150 4088 19156 4140
rect 19208 4128 19214 4140
rect 19812 4128 19840 4168
rect 19208 4118 19334 4128
rect 19628 4118 19840 4128
rect 19208 4100 19840 4118
rect 19996 4128 20024 4168
rect 20438 4156 20444 4208
rect 20496 4156 20502 4208
rect 20622 4156 20628 4208
rect 20680 4205 20686 4208
rect 20680 4199 20699 4205
rect 20687 4165 20699 4199
rect 20680 4159 20699 4165
rect 20680 4156 20686 4159
rect 21082 4156 21088 4208
rect 21140 4196 21146 4208
rect 21269 4199 21327 4205
rect 21269 4196 21281 4199
rect 21140 4168 21281 4196
rect 21140 4156 21146 4168
rect 21269 4165 21281 4168
rect 21315 4165 21327 4199
rect 24118 4196 24124 4208
rect 21269 4159 21327 4165
rect 21657 4168 24124 4196
rect 21361 4131 21419 4137
rect 21361 4128 21373 4131
rect 19996 4100 21373 4128
rect 19208 4088 19214 4100
rect 19306 4090 19656 4100
rect 21361 4097 21373 4100
rect 21407 4097 21419 4131
rect 21361 4091 21419 4097
rect 18782 4020 18788 4072
rect 18840 4060 18846 4072
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 18840 4032 19993 4060
rect 18840 4020 18846 4032
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 20165 4063 20223 4069
rect 20165 4029 20177 4063
rect 20211 4060 20223 4063
rect 20254 4060 20260 4072
rect 20211 4032 20260 4060
rect 20211 4029 20223 4032
rect 20165 4023 20223 4029
rect 20254 4020 20260 4032
rect 20312 4060 20318 4072
rect 21545 4063 21603 4069
rect 21545 4060 21557 4063
rect 20312 4032 21557 4060
rect 20312 4020 20318 4032
rect 21545 4029 21557 4032
rect 21591 4060 21603 4063
rect 21657 4060 21685 4168
rect 24118 4156 24124 4168
rect 24176 4156 24182 4208
rect 25866 4196 25872 4208
rect 25806 4168 25872 4196
rect 25866 4156 25872 4168
rect 25924 4156 25930 4208
rect 27709 4199 27767 4205
rect 26344 4168 26832 4196
rect 22830 4088 22836 4140
rect 22888 4088 22894 4140
rect 23566 4088 23572 4140
rect 23624 4128 23630 4140
rect 24026 4128 24032 4140
rect 23624 4100 24032 4128
rect 23624 4088 23630 4100
rect 24026 4088 24032 4100
rect 24084 4128 24090 4140
rect 24305 4131 24363 4137
rect 24305 4128 24317 4131
rect 24084 4100 24317 4128
rect 24084 4088 24090 4100
rect 24305 4097 24317 4100
rect 24351 4097 24363 4131
rect 24305 4091 24363 4097
rect 26050 4088 26056 4140
rect 26108 4128 26114 4140
rect 26344 4128 26372 4168
rect 26108 4100 26372 4128
rect 26108 4088 26114 4100
rect 26418 4088 26424 4140
rect 26476 4088 26482 4140
rect 26697 4131 26755 4137
rect 26697 4097 26709 4131
rect 26743 4097 26755 4131
rect 26804 4128 26832 4168
rect 27709 4165 27721 4199
rect 27755 4196 27767 4199
rect 27982 4196 27988 4208
rect 27755 4168 27988 4196
rect 27755 4165 27767 4168
rect 27709 4159 27767 4165
rect 27982 4156 27988 4168
rect 28040 4156 28046 4208
rect 28258 4156 28264 4208
rect 28316 4196 28322 4208
rect 30285 4199 30343 4205
rect 30285 4196 30297 4199
rect 28316 4168 30297 4196
rect 28316 4156 28322 4168
rect 30285 4165 30297 4168
rect 30331 4165 30343 4199
rect 30285 4159 30343 4165
rect 30484 4168 31616 4196
rect 26804 4100 28396 4128
rect 26697 4091 26755 4097
rect 21591 4032 21685 4060
rect 21729 4063 21787 4069
rect 21591 4029 21603 4032
rect 21545 4023 21603 4029
rect 21729 4029 21741 4063
rect 21775 4060 21787 4063
rect 21818 4060 21824 4072
rect 21775 4032 21824 4060
rect 21775 4029 21787 4032
rect 21729 4023 21787 4029
rect 21818 4020 21824 4032
rect 21876 4020 21882 4072
rect 22373 4063 22431 4069
rect 22373 4029 22385 4063
rect 22419 4060 22431 4063
rect 22646 4060 22652 4072
rect 22419 4032 22652 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 22646 4020 22652 4032
rect 22704 4020 22710 4072
rect 23658 4020 23664 4072
rect 23716 4020 23722 4072
rect 24581 4063 24639 4069
rect 24581 4060 24593 4063
rect 23768 4032 24593 4060
rect 23768 3992 23796 4032
rect 24581 4029 24593 4032
rect 24627 4029 24639 4063
rect 24581 4023 24639 4029
rect 25958 4020 25964 4072
rect 26016 4060 26022 4072
rect 26329 4063 26387 4069
rect 26329 4060 26341 4063
rect 26016 4032 26341 4060
rect 26016 4020 26022 4032
rect 26329 4029 26341 4032
rect 26375 4060 26387 4063
rect 26712 4060 26740 4091
rect 26375 4032 26740 4060
rect 26375 4029 26387 4032
rect 26329 4023 26387 4029
rect 27062 4020 27068 4072
rect 27120 4060 27126 4072
rect 27341 4063 27399 4069
rect 27341 4060 27353 4063
rect 27120 4032 27353 4060
rect 27120 4020 27126 4032
rect 27341 4029 27353 4032
rect 27387 4029 27399 4063
rect 27341 4023 27399 4029
rect 27562 4063 27620 4069
rect 27562 4029 27574 4063
rect 27608 4060 27620 4063
rect 28368 4060 28396 4100
rect 28442 4088 28448 4140
rect 28500 4088 28506 4140
rect 30484 4128 30512 4168
rect 31110 4128 31116 4140
rect 28920 4100 30512 4128
rect 30576 4100 31116 4128
rect 28920 4060 28948 4100
rect 27608 4032 28304 4060
rect 28368 4032 28948 4060
rect 27608 4029 27620 4032
rect 27562 4023 27620 4029
rect 18340 3964 23796 3992
rect 26694 3952 26700 4004
rect 26752 3952 26758 4004
rect 27249 3995 27307 4001
rect 27249 3961 27261 3995
rect 27295 3992 27307 3995
rect 28276 3992 28304 4032
rect 29086 4020 29092 4072
rect 29144 4020 29150 4072
rect 29638 4020 29644 4072
rect 29696 4060 29702 4072
rect 30576 4069 30604 4100
rect 31110 4088 31116 4100
rect 31168 4088 31174 4140
rect 31588 4128 31616 4168
rect 33428 4168 34560 4196
rect 31588 4100 32628 4128
rect 30377 4063 30435 4069
rect 30377 4060 30389 4063
rect 29696 4032 30389 4060
rect 29696 4020 29702 4032
rect 30377 4029 30389 4032
rect 30423 4029 30435 4063
rect 30377 4023 30435 4029
rect 30561 4063 30619 4069
rect 30561 4029 30573 4063
rect 30607 4029 30619 4063
rect 30561 4023 30619 4029
rect 30837 4063 30895 4069
rect 30837 4029 30849 4063
rect 30883 4060 30895 4063
rect 32401 4063 32459 4069
rect 30883 4032 31708 4060
rect 30883 4029 30895 4032
rect 30837 4023 30895 4029
rect 31680 4004 31708 4032
rect 32401 4029 32413 4063
rect 32447 4060 32459 4063
rect 32490 4060 32496 4072
rect 32447 4032 32496 4060
rect 32447 4029 32459 4032
rect 32401 4023 32459 4029
rect 32490 4020 32496 4032
rect 32548 4020 32554 4072
rect 29178 3992 29184 4004
rect 27295 3964 28212 3992
rect 28276 3964 29184 3992
rect 27295 3961 27307 3964
rect 27249 3955 27307 3961
rect 8619 3896 12112 3924
rect 12253 3927 12311 3933
rect 8619 3893 8631 3896
rect 8573 3887 8631 3893
rect 12253 3893 12265 3927
rect 12299 3924 12311 3927
rect 13262 3924 13268 3936
rect 12299 3896 13268 3924
rect 12299 3893 12311 3896
rect 12253 3887 12311 3893
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 14458 3884 14464 3936
rect 14516 3924 14522 3936
rect 19426 3924 19432 3936
rect 14516 3896 19432 3924
rect 14516 3884 14522 3896
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 19518 3884 19524 3936
rect 19576 3884 19582 3936
rect 20070 3884 20076 3936
rect 20128 3924 20134 3936
rect 20625 3927 20683 3933
rect 20625 3924 20637 3927
rect 20128 3896 20637 3924
rect 20128 3884 20134 3896
rect 20625 3893 20637 3896
rect 20671 3893 20683 3927
rect 20625 3887 20683 3893
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 20809 3927 20867 3933
rect 20809 3924 20821 3927
rect 20772 3896 20821 3924
rect 20772 3884 20778 3896
rect 20809 3893 20821 3896
rect 20855 3893 20867 3927
rect 20809 3887 20867 3893
rect 20898 3884 20904 3936
rect 20956 3884 20962 3936
rect 20990 3884 20996 3936
rect 21048 3924 21054 3936
rect 26418 3924 26424 3936
rect 21048 3896 26424 3924
rect 21048 3884 21054 3896
rect 26418 3884 26424 3896
rect 26476 3884 26482 3936
rect 27430 3884 27436 3936
rect 27488 3884 27494 3936
rect 28184 3924 28212 3964
rect 29178 3952 29184 3964
rect 29236 3952 29242 4004
rect 29454 3952 29460 4004
rect 29512 3992 29518 4004
rect 29917 3995 29975 4001
rect 29917 3992 29929 3995
rect 29512 3964 29929 3992
rect 29512 3952 29518 3964
rect 29917 3961 29929 3964
rect 29963 3961 29975 3995
rect 31570 3992 31576 4004
rect 29917 3955 29975 3961
rect 31312 3964 31576 3992
rect 31312 3924 31340 3964
rect 31570 3952 31576 3964
rect 31628 3952 31634 4004
rect 31662 3952 31668 4004
rect 31720 3952 31726 4004
rect 32600 3992 32628 4100
rect 32674 4088 32680 4140
rect 32732 4088 32738 4140
rect 33042 4088 33048 4140
rect 33100 4088 33106 4140
rect 33226 4088 33232 4140
rect 33284 4088 33290 4140
rect 33428 4137 33456 4168
rect 33413 4131 33471 4137
rect 33413 4097 33425 4131
rect 33459 4097 33471 4131
rect 33413 4091 33471 4097
rect 34057 4131 34115 4137
rect 34057 4097 34069 4131
rect 34103 4097 34115 4131
rect 34532 4128 34560 4168
rect 34606 4156 34612 4208
rect 34664 4196 34670 4208
rect 39942 4196 39948 4208
rect 34664 4168 39948 4196
rect 34664 4156 34670 4168
rect 39942 4156 39948 4168
rect 40000 4156 40006 4208
rect 40034 4156 40040 4208
rect 40092 4196 40098 4208
rect 40092 4168 40526 4196
rect 40092 4156 40098 4168
rect 41598 4156 41604 4208
rect 41656 4196 41662 4208
rect 42242 4196 42248 4208
rect 41656 4168 42248 4196
rect 41656 4156 41662 4168
rect 42242 4156 42248 4168
rect 42300 4156 42306 4208
rect 42610 4156 42616 4208
rect 42668 4196 42674 4208
rect 45370 4196 45376 4208
rect 42668 4168 45376 4196
rect 42668 4156 42674 4168
rect 45370 4156 45376 4168
rect 45428 4156 45434 4208
rect 52638 4156 52644 4208
rect 52696 4156 52702 4208
rect 34532 4100 36032 4128
rect 34057 4091 34115 4097
rect 33962 4020 33968 4072
rect 34020 4020 34026 4072
rect 34072 3992 34100 4091
rect 34514 4020 34520 4072
rect 34572 4060 34578 4072
rect 34882 4060 34888 4072
rect 34572 4032 34888 4060
rect 34572 4020 34578 4032
rect 34882 4020 34888 4032
rect 34940 4020 34946 4072
rect 35069 4063 35127 4069
rect 35069 4029 35081 4063
rect 35115 4029 35127 4063
rect 35069 4023 35127 4029
rect 32600 3964 34100 3992
rect 35084 3992 35112 4023
rect 35158 4020 35164 4072
rect 35216 4060 35222 4072
rect 35897 4063 35955 4069
rect 35897 4060 35909 4063
rect 35216 4032 35909 4060
rect 35216 4020 35222 4032
rect 35897 4029 35909 4032
rect 35943 4029 35955 4063
rect 35897 4023 35955 4029
rect 35250 3992 35256 4004
rect 35084 3964 35256 3992
rect 35250 3952 35256 3964
rect 35308 3952 35314 4004
rect 28184 3896 31340 3924
rect 31389 3927 31447 3933
rect 31389 3893 31401 3927
rect 31435 3924 31447 3927
rect 32766 3924 32772 3936
rect 31435 3896 32772 3924
rect 31435 3893 31447 3896
rect 31389 3887 31447 3893
rect 32766 3884 32772 3896
rect 32824 3884 32830 3936
rect 33045 3927 33103 3933
rect 33045 3893 33057 3927
rect 33091 3924 33103 3927
rect 35526 3924 35532 3936
rect 33091 3896 35532 3924
rect 33091 3893 33103 3896
rect 33045 3887 33103 3893
rect 35526 3884 35532 3896
rect 35584 3884 35590 3936
rect 35912 3924 35940 4023
rect 36004 3992 36032 4100
rect 36078 4088 36084 4140
rect 36136 4088 36142 4140
rect 36170 4088 36176 4140
rect 36228 4088 36234 4140
rect 36814 4088 36820 4140
rect 36872 4088 36878 4140
rect 38194 4088 38200 4140
rect 38252 4088 38258 4140
rect 38381 4131 38439 4137
rect 38381 4097 38393 4131
rect 38427 4128 38439 4131
rect 38562 4128 38568 4140
rect 38427 4100 38568 4128
rect 38427 4097 38439 4100
rect 38381 4091 38439 4097
rect 38562 4088 38568 4100
rect 38620 4088 38626 4140
rect 38654 4088 38660 4140
rect 38712 4088 38718 4140
rect 42705 4131 42763 4137
rect 42705 4097 42717 4131
rect 42751 4128 42763 4131
rect 45649 4131 45707 4137
rect 45649 4128 45661 4131
rect 42751 4100 45661 4128
rect 42751 4097 42763 4100
rect 42705 4091 42763 4097
rect 45649 4097 45661 4100
rect 45695 4097 45707 4131
rect 47857 4131 47915 4137
rect 47857 4128 47869 4131
rect 45649 4091 45707 4097
rect 45756 4100 47869 4128
rect 37274 4020 37280 4072
rect 37332 4020 37338 4072
rect 38102 4020 38108 4072
rect 38160 4060 38166 4072
rect 39025 4063 39083 4069
rect 39025 4060 39037 4063
rect 38160 4032 39037 4060
rect 38160 4020 38166 4032
rect 39025 4029 39037 4032
rect 39071 4029 39083 4063
rect 41598 4060 41604 4072
rect 39025 4023 39083 4029
rect 39132 4032 41604 4060
rect 39132 3992 39160 4032
rect 41598 4020 41604 4032
rect 41656 4020 41662 4072
rect 41690 4020 41696 4072
rect 41748 4020 41754 4072
rect 41969 4063 42027 4069
rect 41969 4029 41981 4063
rect 42015 4029 42027 4063
rect 41969 4023 42027 4029
rect 42153 4063 42211 4069
rect 42153 4029 42165 4063
rect 42199 4060 42211 4063
rect 42794 4060 42800 4072
rect 42199 4032 42800 4060
rect 42199 4029 42211 4032
rect 42153 4023 42211 4029
rect 36004 3964 39160 3992
rect 41984 3992 42012 4023
rect 42794 4020 42800 4032
rect 42852 4020 42858 4072
rect 43070 4020 43076 4072
rect 43128 4060 43134 4072
rect 43441 4063 43499 4069
rect 43441 4060 43453 4063
rect 43128 4032 43453 4060
rect 43128 4020 43134 4032
rect 43441 4029 43453 4032
rect 43487 4029 43499 4063
rect 43441 4023 43499 4029
rect 43806 4020 43812 4072
rect 43864 4060 43870 4072
rect 44177 4063 44235 4069
rect 44177 4060 44189 4063
rect 43864 4032 44189 4060
rect 43864 4020 43870 4032
rect 44177 4029 44189 4032
rect 44223 4029 44235 4063
rect 44177 4023 44235 4029
rect 44818 4020 44824 4072
rect 44876 4020 44882 4072
rect 44910 4020 44916 4072
rect 44968 4020 44974 4072
rect 45557 4063 45615 4069
rect 45557 4029 45569 4063
rect 45603 4029 45615 4063
rect 45557 4023 45615 4029
rect 42242 3992 42248 4004
rect 41984 3964 42248 3992
rect 42242 3952 42248 3964
rect 42300 3952 42306 4004
rect 43254 3952 43260 4004
rect 43312 3992 43318 4004
rect 45572 3992 45600 4023
rect 43312 3964 45600 3992
rect 43312 3952 43318 3964
rect 36446 3924 36452 3936
rect 35912 3896 36452 3924
rect 36446 3884 36452 3896
rect 36504 3884 36510 3936
rect 36541 3927 36599 3933
rect 36541 3893 36553 3927
rect 36587 3924 36599 3927
rect 37182 3924 37188 3936
rect 36587 3896 37188 3924
rect 36587 3893 36599 3896
rect 36541 3887 36599 3893
rect 37182 3884 37188 3896
rect 37240 3884 37246 3936
rect 38930 3884 38936 3936
rect 38988 3924 38994 3936
rect 42886 3924 42892 3936
rect 38988 3896 42892 3924
rect 38988 3884 38994 3896
rect 42886 3884 42892 3896
rect 42944 3884 42950 3936
rect 43530 3884 43536 3936
rect 43588 3924 43594 3936
rect 44085 3927 44143 3933
rect 44085 3924 44097 3927
rect 43588 3896 44097 3924
rect 43588 3884 43594 3896
rect 44085 3893 44097 3896
rect 44131 3924 44143 3927
rect 45756 3924 45784 4100
rect 47857 4097 47869 4100
rect 47903 4097 47915 4131
rect 47857 4091 47915 4097
rect 50522 4088 50528 4140
rect 50580 4088 50586 4140
rect 74626 4088 74632 4140
rect 74684 4128 74690 4140
rect 74721 4131 74779 4137
rect 74721 4128 74733 4131
rect 74684 4100 74733 4128
rect 74684 4088 74690 4100
rect 74721 4097 74733 4100
rect 74767 4097 74779 4131
rect 76193 4131 76251 4137
rect 76193 4128 76205 4131
rect 74721 4091 74779 4097
rect 75288 4100 76205 4128
rect 46934 4020 46940 4072
rect 46992 4020 46998 4072
rect 47118 4020 47124 4072
rect 47176 4020 47182 4072
rect 47210 4020 47216 4072
rect 47268 4060 47274 4072
rect 48501 4063 48559 4069
rect 48501 4060 48513 4063
rect 47268 4032 48513 4060
rect 47268 4020 47274 4032
rect 48501 4029 48513 4032
rect 48547 4029 48559 4063
rect 48501 4023 48559 4029
rect 48590 4020 48596 4072
rect 48648 4060 48654 4072
rect 49053 4063 49111 4069
rect 49053 4060 49065 4063
rect 48648 4032 49065 4060
rect 48648 4020 48654 4032
rect 49053 4029 49065 4032
rect 49099 4029 49111 4063
rect 49053 4023 49111 4029
rect 49881 4063 49939 4069
rect 49881 4029 49893 4063
rect 49927 4060 49939 4063
rect 50062 4060 50068 4072
rect 49927 4032 50068 4060
rect 49927 4029 49939 4032
rect 49881 4023 49939 4029
rect 50062 4020 50068 4032
rect 50120 4020 50126 4072
rect 65426 4020 65432 4072
rect 65484 4060 65490 4072
rect 65521 4063 65579 4069
rect 65521 4060 65533 4063
rect 65484 4032 65533 4060
rect 65484 4020 65490 4032
rect 65521 4029 65533 4032
rect 65567 4029 65579 4063
rect 65521 4023 65579 4029
rect 67637 4063 67695 4069
rect 67637 4029 67649 4063
rect 67683 4060 67695 4063
rect 67910 4060 67916 4072
rect 67683 4032 67916 4060
rect 67683 4029 67695 4032
rect 67637 4023 67695 4029
rect 67910 4020 67916 4032
rect 67968 4020 67974 4072
rect 71501 4063 71559 4069
rect 71501 4029 71513 4063
rect 71547 4060 71559 4063
rect 71682 4060 71688 4072
rect 71547 4032 71688 4060
rect 71547 4029 71559 4032
rect 71501 4023 71559 4029
rect 71682 4020 71688 4032
rect 71740 4020 71746 4072
rect 74074 4020 74080 4072
rect 74132 4060 74138 4072
rect 75288 4060 75316 4100
rect 76193 4097 76205 4100
rect 76239 4097 76251 4131
rect 76193 4091 76251 4097
rect 74132 4032 75316 4060
rect 75917 4063 75975 4069
rect 74132 4020 74138 4032
rect 75917 4029 75929 4063
rect 75963 4060 75975 4063
rect 76558 4060 76564 4072
rect 75963 4032 76564 4060
rect 75963 4029 75975 4032
rect 75917 4023 75975 4029
rect 76558 4020 76564 4032
rect 76616 4020 76622 4072
rect 77018 4020 77024 4072
rect 77076 4020 77082 4072
rect 48041 3995 48099 4001
rect 48041 3961 48053 3995
rect 48087 3992 48099 3995
rect 48866 3992 48872 4004
rect 48087 3964 48872 3992
rect 48087 3961 48099 3964
rect 48041 3955 48099 3961
rect 48866 3952 48872 3964
rect 48924 3952 48930 4004
rect 44131 3896 45784 3924
rect 44131 3893 44143 3896
rect 44085 3887 44143 3893
rect 46106 3884 46112 3936
rect 46164 3924 46170 3936
rect 46293 3927 46351 3933
rect 46293 3924 46305 3927
rect 46164 3896 46305 3924
rect 46164 3884 46170 3896
rect 46293 3893 46305 3896
rect 46339 3893 46351 3927
rect 46293 3887 46351 3893
rect 46382 3884 46388 3936
rect 46440 3884 46446 3936
rect 47486 3884 47492 3936
rect 47544 3924 47550 3936
rect 47765 3927 47823 3933
rect 47765 3924 47777 3927
rect 47544 3896 47777 3924
rect 47544 3884 47550 3896
rect 47765 3893 47777 3896
rect 47811 3893 47823 3927
rect 47765 3887 47823 3893
rect 49234 3884 49240 3936
rect 49292 3884 49298 3936
rect 49878 3884 49884 3936
rect 49936 3924 49942 3936
rect 49973 3927 50031 3933
rect 49973 3924 49985 3927
rect 49936 3896 49985 3924
rect 49936 3884 49942 3896
rect 49973 3893 49985 3896
rect 50019 3893 50031 3927
rect 49973 3887 50031 3893
rect 51074 3884 51080 3936
rect 51132 3924 51138 3936
rect 52362 3924 52368 3936
rect 51132 3896 52368 3924
rect 51132 3884 51138 3896
rect 52362 3884 52368 3896
rect 52420 3924 52426 3936
rect 52733 3927 52791 3933
rect 52733 3924 52745 3927
rect 52420 3896 52745 3924
rect 52420 3884 52426 3896
rect 52733 3893 52745 3896
rect 52779 3893 52791 3927
rect 52733 3887 52791 3893
rect 66165 3927 66223 3933
rect 66165 3893 66177 3927
rect 66211 3924 66223 3927
rect 66254 3924 66260 3936
rect 66211 3896 66260 3924
rect 66211 3893 66223 3896
rect 66165 3887 66223 3893
rect 66254 3884 66260 3896
rect 66312 3884 66318 3936
rect 68189 3927 68247 3933
rect 68189 3893 68201 3927
rect 68235 3924 68247 3927
rect 68278 3924 68284 3936
rect 68235 3896 68284 3924
rect 68235 3893 68247 3896
rect 68189 3887 68247 3893
rect 68278 3884 68284 3896
rect 68336 3884 68342 3936
rect 72053 3927 72111 3933
rect 72053 3893 72065 3927
rect 72099 3924 72111 3927
rect 72418 3924 72424 3936
rect 72099 3896 72424 3924
rect 72099 3893 72111 3896
rect 72053 3887 72111 3893
rect 72418 3884 72424 3896
rect 72476 3884 72482 3936
rect 2024 3834 77924 3856
rect 2024 3782 5134 3834
rect 5186 3782 5198 3834
rect 5250 3782 5262 3834
rect 5314 3782 5326 3834
rect 5378 3782 5390 3834
rect 5442 3782 35854 3834
rect 35906 3782 35918 3834
rect 35970 3782 35982 3834
rect 36034 3782 36046 3834
rect 36098 3782 36110 3834
rect 36162 3782 66574 3834
rect 66626 3782 66638 3834
rect 66690 3782 66702 3834
rect 66754 3782 66766 3834
rect 66818 3782 66830 3834
rect 66882 3782 77924 3834
rect 2024 3760 77924 3782
rect 4893 3723 4951 3729
rect 4893 3689 4905 3723
rect 4939 3720 4951 3723
rect 5718 3720 5724 3732
rect 4939 3692 5724 3720
rect 4939 3689 4951 3692
rect 4893 3683 4951 3689
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 5994 3680 6000 3732
rect 6052 3680 6058 3732
rect 6886 3692 9812 3720
rect 6886 3652 6914 3692
rect 5460 3624 6914 3652
rect 7469 3655 7527 3661
rect 5460 3593 5488 3624
rect 7469 3621 7481 3655
rect 7515 3652 7527 3655
rect 8294 3652 8300 3664
rect 7515 3624 8300 3652
rect 7515 3621 7527 3624
rect 7469 3615 7527 3621
rect 8294 3612 8300 3624
rect 8352 3612 8358 3664
rect 9784 3652 9812 3692
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 9916 3692 10885 3720
rect 9916 3680 9922 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 10873 3683 10931 3689
rect 11882 3680 11888 3732
rect 11940 3680 11946 3732
rect 14829 3723 14887 3729
rect 12084 3692 14780 3720
rect 10686 3652 10692 3664
rect 9784 3624 10692 3652
rect 10686 3612 10692 3624
rect 10744 3612 10750 3664
rect 10781 3655 10839 3661
rect 10781 3621 10793 3655
rect 10827 3652 10839 3655
rect 12084 3652 12112 3692
rect 10827 3624 12112 3652
rect 10827 3621 10839 3624
rect 10781 3615 10839 3621
rect 14090 3612 14096 3664
rect 14148 3612 14154 3664
rect 14752 3652 14780 3692
rect 14829 3689 14841 3723
rect 14875 3720 14887 3723
rect 16574 3720 16580 3732
rect 14875 3692 16580 3720
rect 14875 3689 14887 3692
rect 14829 3683 14887 3689
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 16758 3680 16764 3732
rect 16816 3720 16822 3732
rect 22094 3720 22100 3732
rect 16816 3692 18736 3720
rect 16816 3680 16822 3692
rect 16482 3652 16488 3664
rect 14752 3624 16488 3652
rect 16482 3612 16488 3624
rect 16540 3612 16546 3664
rect 5445 3587 5503 3593
rect 4724 3556 5396 3584
rect 4724 3525 4752 3556
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 5074 3476 5080 3528
rect 5132 3476 5138 3528
rect 5368 3516 5396 3556
rect 5445 3553 5457 3587
rect 5491 3553 5503 3587
rect 6270 3584 6276 3596
rect 5445 3547 5503 3553
rect 5552 3556 6276 3584
rect 5552 3516 5580 3556
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 6822 3544 6828 3596
rect 6880 3544 6886 3596
rect 9033 3587 9091 3593
rect 9033 3584 9045 3587
rect 7024 3556 9045 3584
rect 5368 3488 5580 3516
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 5684 3488 6101 3516
rect 5684 3476 5690 3488
rect 6089 3485 6101 3488
rect 6135 3485 6147 3519
rect 6089 3479 6147 3485
rect 6178 3476 6184 3528
rect 6236 3516 6242 3528
rect 7024 3516 7052 3556
rect 9033 3553 9045 3556
rect 9079 3553 9091 3587
rect 9033 3547 9091 3553
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 12253 3587 12311 3593
rect 12253 3584 12265 3587
rect 9180 3556 12265 3584
rect 9180 3544 9186 3556
rect 12253 3553 12265 3556
rect 12299 3553 12311 3587
rect 12253 3547 12311 3553
rect 12802 3544 12808 3596
rect 12860 3584 12866 3596
rect 13725 3587 13783 3593
rect 13725 3584 13737 3587
rect 12860 3556 13737 3584
rect 12860 3544 12866 3556
rect 13725 3553 13737 3556
rect 13771 3553 13783 3587
rect 13725 3547 13783 3553
rect 14274 3544 14280 3596
rect 14332 3544 14338 3596
rect 15470 3544 15476 3596
rect 15528 3544 15534 3596
rect 15657 3587 15715 3593
rect 15657 3553 15669 3587
rect 15703 3584 15715 3587
rect 15746 3584 15752 3596
rect 15703 3556 15752 3584
rect 15703 3553 15715 3556
rect 15657 3547 15715 3553
rect 15746 3544 15752 3556
rect 15804 3544 15810 3596
rect 17310 3544 17316 3596
rect 17368 3584 17374 3596
rect 18708 3593 18736 3692
rect 19996 3692 22100 3720
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 19797 3655 19855 3661
rect 19797 3652 19809 3655
rect 19484 3624 19809 3652
rect 19484 3612 19490 3624
rect 19797 3621 19809 3624
rect 19843 3621 19855 3655
rect 19797 3615 19855 3621
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 17368 3556 17877 3584
rect 17368 3544 17374 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 18693 3587 18751 3593
rect 18693 3553 18705 3587
rect 18739 3553 18751 3587
rect 18693 3547 18751 3553
rect 6236 3488 7052 3516
rect 6236 3476 6242 3488
rect 7650 3476 7656 3528
rect 7708 3476 7714 3528
rect 8202 3476 8208 3528
rect 8260 3476 8266 3528
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3516 9735 3519
rect 9766 3516 9772 3528
rect 9723 3488 9772 3516
rect 9723 3485 9735 3488
rect 9677 3479 9735 3485
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 10226 3476 10232 3528
rect 10284 3476 10290 3528
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3485 11483 3519
rect 11425 3479 11483 3485
rect 7466 3448 7472 3460
rect 5276 3420 7472 3448
rect 5276 3389 5304 3420
rect 7466 3408 7472 3420
rect 7524 3408 7530 3460
rect 8941 3451 8999 3457
rect 8941 3417 8953 3451
rect 8987 3448 8999 3451
rect 11440 3448 11468 3479
rect 11698 3476 11704 3528
rect 11756 3476 11762 3528
rect 11977 3519 12035 3525
rect 11977 3485 11989 3519
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3516 13967 3519
rect 13998 3516 14004 3528
rect 13955 3488 14004 3516
rect 13955 3485 13967 3488
rect 13909 3479 13967 3485
rect 8987 3420 11468 3448
rect 11992 3448 12020 3479
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 15286 3476 15292 3528
rect 15344 3516 15350 3528
rect 15381 3519 15439 3525
rect 15381 3516 15393 3519
rect 15344 3488 15393 3516
rect 15344 3476 15350 3488
rect 15381 3485 15393 3488
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 15488 3488 16528 3516
rect 12158 3448 12164 3460
rect 11992 3420 12164 3448
rect 8987 3417 8999 3420
rect 8941 3411 8999 3417
rect 12158 3408 12164 3420
rect 12216 3408 12222 3460
rect 12710 3408 12716 3460
rect 12768 3408 12774 3460
rect 15488 3448 15516 3488
rect 13556 3420 15516 3448
rect 5261 3383 5319 3389
rect 5261 3349 5273 3383
rect 5307 3349 5319 3383
rect 5261 3343 5319 3349
rect 6730 3340 6736 3392
rect 6788 3340 6794 3392
rect 10045 3383 10103 3389
rect 10045 3349 10057 3383
rect 10091 3380 10103 3383
rect 10134 3380 10140 3392
rect 10091 3352 10140 3380
rect 10091 3349 10103 3352
rect 10045 3343 10103 3349
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 11422 3340 11428 3392
rect 11480 3380 11486 3392
rect 13556 3380 13584 3420
rect 15930 3408 15936 3460
rect 15988 3408 15994 3460
rect 11480 3352 13584 3380
rect 11480 3340 11486 3352
rect 13722 3340 13728 3392
rect 13780 3380 13786 3392
rect 15013 3383 15071 3389
rect 15013 3380 15025 3383
rect 13780 3352 15025 3380
rect 13780 3340 13786 3352
rect 15013 3349 15025 3352
rect 15059 3349 15071 3383
rect 15013 3343 15071 3349
rect 16206 3340 16212 3392
rect 16264 3340 16270 3392
rect 16390 3340 16396 3392
rect 16448 3340 16454 3392
rect 16500 3380 16528 3488
rect 18138 3476 18144 3528
rect 18196 3476 18202 3528
rect 18230 3476 18236 3528
rect 18288 3476 18294 3528
rect 16850 3408 16856 3460
rect 16908 3408 16914 3460
rect 17954 3408 17960 3460
rect 18012 3448 18018 3460
rect 19812 3448 19840 3615
rect 19996 3525 20024 3692
rect 22094 3680 22100 3692
rect 22152 3720 22158 3732
rect 22152 3692 28212 3720
rect 22152 3680 22158 3692
rect 20070 3612 20076 3664
rect 20128 3652 20134 3664
rect 21450 3652 21456 3664
rect 20128 3624 21456 3652
rect 20128 3612 20134 3624
rect 21450 3612 21456 3624
rect 21508 3612 21514 3664
rect 24210 3612 24216 3664
rect 24268 3652 24274 3664
rect 24268 3624 25360 3652
rect 24268 3612 24274 3624
rect 20806 3544 20812 3596
rect 20864 3544 20870 3596
rect 22830 3544 22836 3596
rect 22888 3544 22894 3596
rect 19981 3519 20039 3525
rect 19981 3485 19993 3519
rect 20027 3485 20039 3519
rect 19981 3479 20039 3485
rect 20346 3476 20352 3528
rect 20404 3476 20410 3528
rect 20438 3476 20444 3528
rect 20496 3516 20502 3528
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 20496 3488 21925 3516
rect 20496 3476 20502 3488
rect 21913 3485 21925 3488
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 23198 3476 23204 3528
rect 23256 3516 23262 3528
rect 24394 3516 24400 3528
rect 23256 3488 24400 3516
rect 23256 3476 23262 3488
rect 24394 3476 24400 3488
rect 24452 3476 24458 3528
rect 24670 3476 24676 3528
rect 24728 3516 24734 3528
rect 25332 3525 25360 3624
rect 25590 3612 25596 3664
rect 25648 3612 25654 3664
rect 26142 3544 26148 3596
rect 26200 3544 26206 3596
rect 26329 3587 26387 3593
rect 26329 3553 26341 3587
rect 26375 3584 26387 3587
rect 27614 3584 27620 3596
rect 26375 3556 27620 3584
rect 26375 3553 26387 3556
rect 26329 3547 26387 3553
rect 25133 3519 25191 3525
rect 25133 3516 25145 3519
rect 24728 3488 25145 3516
rect 24728 3476 24734 3488
rect 25133 3485 25145 3488
rect 25179 3485 25191 3519
rect 25133 3479 25191 3485
rect 25317 3519 25375 3525
rect 25317 3485 25329 3519
rect 25363 3485 25375 3519
rect 26344 3516 26372 3547
rect 27614 3544 27620 3556
rect 27672 3544 27678 3596
rect 25317 3479 25375 3485
rect 25424 3488 26372 3516
rect 18012 3420 19748 3448
rect 19812 3420 21956 3448
rect 18012 3408 18018 3420
rect 18598 3380 18604 3392
rect 16500 3352 18604 3380
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 19720 3380 19748 3420
rect 20070 3380 20076 3392
rect 19720 3352 20076 3380
rect 20070 3340 20076 3352
rect 20128 3340 20134 3392
rect 20257 3383 20315 3389
rect 20257 3349 20269 3383
rect 20303 3380 20315 3383
rect 21818 3380 21824 3392
rect 20303 3352 21824 3380
rect 20303 3349 20315 3352
rect 20257 3343 20315 3349
rect 21818 3340 21824 3352
rect 21876 3340 21882 3392
rect 21928 3380 21956 3420
rect 22094 3408 22100 3460
rect 22152 3448 22158 3460
rect 22462 3448 22468 3460
rect 22152 3420 22468 3448
rect 22152 3408 22158 3420
rect 22462 3408 22468 3420
rect 22520 3408 22526 3460
rect 24118 3408 24124 3460
rect 24176 3448 24182 3460
rect 25424 3448 25452 3488
rect 26602 3476 26608 3528
rect 26660 3516 26666 3528
rect 26697 3519 26755 3525
rect 26697 3516 26709 3519
rect 26660 3488 26709 3516
rect 26660 3476 26666 3488
rect 26697 3485 26709 3488
rect 26743 3485 26755 3519
rect 28184 3516 28212 3692
rect 28350 3680 28356 3732
rect 28408 3720 28414 3732
rect 28445 3723 28503 3729
rect 28445 3720 28457 3723
rect 28408 3692 28457 3720
rect 28408 3680 28414 3692
rect 28445 3689 28457 3692
rect 28491 3689 28503 3723
rect 28445 3683 28503 3689
rect 28718 3680 28724 3732
rect 28776 3680 28782 3732
rect 30282 3680 30288 3732
rect 30340 3720 30346 3732
rect 32125 3723 32183 3729
rect 32125 3720 32137 3723
rect 30340 3692 32137 3720
rect 30340 3680 30346 3692
rect 32125 3689 32137 3692
rect 32171 3689 32183 3723
rect 32125 3683 32183 3689
rect 33318 3680 33324 3732
rect 33376 3720 33382 3732
rect 34149 3723 34207 3729
rect 34149 3720 34161 3723
rect 33376 3692 34161 3720
rect 33376 3680 33382 3692
rect 34149 3689 34161 3692
rect 34195 3689 34207 3723
rect 34149 3683 34207 3689
rect 34238 3680 34244 3732
rect 34296 3680 34302 3732
rect 34701 3723 34759 3729
rect 34701 3689 34713 3723
rect 34747 3720 34759 3723
rect 34790 3720 34796 3732
rect 34747 3692 34796 3720
rect 34747 3689 34759 3692
rect 34701 3683 34759 3689
rect 34790 3680 34796 3692
rect 34848 3680 34854 3732
rect 35710 3680 35716 3732
rect 35768 3720 35774 3732
rect 35805 3723 35863 3729
rect 35805 3720 35817 3723
rect 35768 3692 35817 3720
rect 35768 3680 35774 3692
rect 35805 3689 35817 3692
rect 35851 3689 35863 3723
rect 35805 3683 35863 3689
rect 36446 3680 36452 3732
rect 36504 3720 36510 3732
rect 40310 3720 40316 3732
rect 36504 3692 40316 3720
rect 36504 3680 36510 3692
rect 40310 3680 40316 3692
rect 40368 3680 40374 3732
rect 44821 3723 44879 3729
rect 40420 3692 41920 3720
rect 28736 3652 28764 3680
rect 31846 3652 31852 3664
rect 28736 3624 31852 3652
rect 31846 3612 31852 3624
rect 31904 3612 31910 3664
rect 31941 3655 31999 3661
rect 31941 3621 31953 3655
rect 31987 3652 31999 3655
rect 32030 3652 32036 3664
rect 31987 3624 32036 3652
rect 31987 3621 31999 3624
rect 31941 3615 31999 3621
rect 32030 3612 32036 3624
rect 32088 3612 32094 3664
rect 38930 3652 38936 3664
rect 34624 3624 38936 3652
rect 28350 3544 28356 3596
rect 28408 3584 28414 3596
rect 29365 3587 29423 3593
rect 29365 3584 29377 3587
rect 28408 3556 29377 3584
rect 28408 3544 28414 3556
rect 29365 3553 29377 3556
rect 29411 3553 29423 3587
rect 29365 3547 29423 3553
rect 30374 3544 30380 3596
rect 30432 3584 30438 3596
rect 31294 3584 31300 3596
rect 30432 3556 31300 3584
rect 30432 3544 30438 3556
rect 31294 3544 31300 3556
rect 31352 3584 31358 3596
rect 32401 3587 32459 3593
rect 32401 3584 32413 3587
rect 31352 3556 32413 3584
rect 31352 3544 31358 3556
rect 32401 3553 32413 3556
rect 32447 3553 32459 3587
rect 32401 3547 32459 3553
rect 32766 3544 32772 3596
rect 32824 3584 32830 3596
rect 34624 3593 34652 3624
rect 38930 3612 38936 3624
rect 38988 3612 38994 3664
rect 40420 3652 40448 3692
rect 41601 3655 41659 3661
rect 41601 3652 41613 3655
rect 39316 3624 40448 3652
rect 40696 3624 41613 3652
rect 34609 3587 34667 3593
rect 32824 3556 34560 3584
rect 32824 3544 32830 3556
rect 28629 3519 28687 3525
rect 28629 3516 28641 3519
rect 28184 3488 28641 3516
rect 26697 3479 26755 3485
rect 28629 3485 28641 3488
rect 28675 3485 28687 3519
rect 28629 3479 28687 3485
rect 29086 3476 29092 3528
rect 29144 3476 29150 3528
rect 30282 3476 30288 3528
rect 30340 3516 30346 3528
rect 30469 3519 30527 3525
rect 30469 3516 30481 3519
rect 30340 3488 30481 3516
rect 30340 3476 30346 3488
rect 30469 3485 30481 3488
rect 30515 3485 30527 3519
rect 30469 3479 30527 3485
rect 30742 3476 30748 3528
rect 30800 3516 30806 3528
rect 31202 3516 31208 3528
rect 30800 3488 31208 3516
rect 30800 3476 30806 3488
rect 31202 3476 31208 3488
rect 31260 3476 31266 3528
rect 34422 3476 34428 3528
rect 34480 3476 34486 3528
rect 34532 3516 34560 3556
rect 34609 3553 34621 3587
rect 34655 3553 34667 3587
rect 34609 3547 34667 3553
rect 35158 3544 35164 3596
rect 35216 3584 35222 3596
rect 35253 3587 35311 3593
rect 35253 3584 35265 3587
rect 35216 3556 35265 3584
rect 35216 3544 35222 3556
rect 35253 3553 35265 3556
rect 35299 3553 35311 3587
rect 35253 3547 35311 3553
rect 35434 3544 35440 3596
rect 35492 3584 35498 3596
rect 35492 3556 36768 3584
rect 35492 3544 35498 3556
rect 36357 3519 36415 3525
rect 34532 3488 35848 3516
rect 24176 3420 25452 3448
rect 25593 3451 25651 3457
rect 24176 3408 24182 3420
rect 25593 3417 25605 3451
rect 25639 3448 25651 3451
rect 26053 3451 26111 3457
rect 25639 3420 25820 3448
rect 25639 3417 25651 3420
rect 25593 3411 25651 3417
rect 22738 3380 22744 3392
rect 21928 3352 22744 3380
rect 22738 3340 22744 3352
rect 22796 3380 22802 3392
rect 23382 3380 23388 3392
rect 22796 3352 23388 3380
rect 22796 3340 22802 3352
rect 23382 3340 23388 3352
rect 23440 3340 23446 3392
rect 23845 3383 23903 3389
rect 23845 3349 23857 3383
rect 23891 3380 23903 3383
rect 24486 3380 24492 3392
rect 23891 3352 24492 3380
rect 23891 3349 23903 3352
rect 23845 3343 23903 3349
rect 24486 3340 24492 3352
rect 24544 3340 24550 3392
rect 25406 3340 25412 3392
rect 25464 3340 25470 3392
rect 25682 3340 25688 3392
rect 25740 3340 25746 3392
rect 25792 3380 25820 3420
rect 26053 3417 26065 3451
rect 26099 3448 26111 3451
rect 26878 3448 26884 3460
rect 26099 3420 26884 3448
rect 26099 3417 26111 3420
rect 26053 3411 26111 3417
rect 26878 3408 26884 3420
rect 26936 3408 26942 3460
rect 26973 3451 27031 3457
rect 26973 3417 26985 3451
rect 27019 3417 27031 3451
rect 28534 3448 28540 3460
rect 28198 3420 28540 3448
rect 26973 3411 27031 3417
rect 26142 3380 26148 3392
rect 25792 3352 26148 3380
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 26326 3340 26332 3392
rect 26384 3380 26390 3392
rect 26605 3383 26663 3389
rect 26605 3380 26617 3383
rect 26384 3352 26617 3380
rect 26384 3340 26390 3352
rect 26605 3349 26617 3352
rect 26651 3380 26663 3383
rect 26694 3380 26700 3392
rect 26651 3352 26700 3380
rect 26651 3349 26663 3352
rect 26605 3343 26663 3349
rect 26694 3340 26700 3352
rect 26752 3340 26758 3392
rect 26786 3340 26792 3392
rect 26844 3380 26850 3392
rect 26988 3380 27016 3411
rect 28534 3408 28540 3420
rect 28592 3408 28598 3460
rect 30190 3408 30196 3460
rect 30248 3448 30254 3460
rect 30374 3448 30380 3460
rect 30248 3420 30380 3448
rect 30248 3408 30254 3420
rect 30374 3408 30380 3420
rect 30432 3408 30438 3460
rect 30558 3408 30564 3460
rect 30616 3448 30622 3460
rect 31389 3451 31447 3457
rect 31389 3448 31401 3451
rect 30616 3420 31401 3448
rect 30616 3408 30622 3420
rect 31389 3417 31401 3420
rect 31435 3417 31447 3451
rect 31389 3411 31447 3417
rect 31846 3408 31852 3460
rect 31904 3448 31910 3460
rect 32309 3451 32367 3457
rect 32309 3448 32321 3451
rect 31904 3420 32321 3448
rect 31904 3408 31910 3420
rect 32309 3417 32321 3420
rect 32355 3417 32367 3451
rect 32309 3411 32367 3417
rect 32398 3408 32404 3460
rect 32456 3448 32462 3460
rect 32677 3451 32735 3457
rect 32677 3448 32689 3451
rect 32456 3420 32689 3448
rect 32456 3408 32462 3420
rect 32677 3417 32689 3420
rect 32723 3417 32735 3451
rect 32677 3411 32735 3417
rect 32950 3408 32956 3460
rect 33008 3448 33014 3460
rect 34974 3448 34980 3460
rect 33008 3420 33166 3448
rect 33980 3420 34980 3448
rect 33008 3408 33014 3420
rect 26844 3352 27016 3380
rect 26844 3340 26850 3352
rect 27982 3340 27988 3392
rect 28040 3380 28046 3392
rect 30466 3380 30472 3392
rect 28040 3352 30472 3380
rect 28040 3340 28046 3352
rect 30466 3340 30472 3352
rect 30524 3340 30530 3392
rect 30650 3340 30656 3392
rect 30708 3380 30714 3392
rect 32109 3383 32167 3389
rect 32109 3380 32121 3383
rect 30708 3352 32121 3380
rect 30708 3340 30714 3352
rect 32109 3349 32121 3352
rect 32155 3380 32167 3383
rect 33980 3380 34008 3420
rect 34974 3408 34980 3420
rect 35032 3408 35038 3460
rect 35066 3408 35072 3460
rect 35124 3408 35130 3460
rect 35710 3408 35716 3460
rect 35768 3408 35774 3460
rect 35820 3448 35848 3488
rect 36357 3485 36369 3519
rect 36403 3516 36415 3519
rect 36630 3516 36636 3528
rect 36403 3488 36636 3516
rect 36403 3485 36415 3488
rect 36357 3479 36415 3485
rect 36630 3476 36636 3488
rect 36688 3476 36694 3528
rect 36740 3516 36768 3556
rect 36814 3544 36820 3596
rect 36872 3544 36878 3596
rect 37660 3556 37872 3584
rect 37660 3516 37688 3556
rect 36740 3488 37688 3516
rect 37737 3519 37795 3525
rect 37737 3485 37749 3519
rect 37783 3485 37795 3519
rect 37844 3516 37872 3556
rect 38654 3544 38660 3596
rect 38712 3544 38718 3596
rect 39209 3519 39267 3525
rect 39209 3516 39221 3519
rect 37844 3488 39221 3516
rect 37737 3479 37795 3485
rect 39209 3485 39221 3488
rect 39255 3485 39267 3519
rect 39209 3479 39267 3485
rect 37752 3448 37780 3479
rect 35820 3420 37780 3448
rect 37918 3408 37924 3460
rect 37976 3448 37982 3460
rect 39316 3448 39344 3624
rect 39669 3587 39727 3593
rect 39669 3553 39681 3587
rect 39715 3553 39727 3587
rect 39669 3547 39727 3553
rect 37976 3420 39344 3448
rect 37976 3408 37982 3420
rect 32155 3352 34008 3380
rect 32155 3349 32167 3352
rect 32109 3343 32167 3349
rect 34606 3340 34612 3392
rect 34664 3380 34670 3392
rect 35084 3380 35112 3408
rect 34664 3352 35112 3380
rect 35161 3383 35219 3389
rect 34664 3340 34670 3352
rect 35161 3349 35173 3383
rect 35207 3380 35219 3383
rect 37090 3380 37096 3392
rect 35207 3352 37096 3380
rect 35207 3349 35219 3352
rect 35161 3343 35219 3349
rect 37090 3340 37096 3352
rect 37148 3340 37154 3392
rect 38746 3340 38752 3392
rect 38804 3380 38810 3392
rect 39684 3380 39712 3547
rect 39758 3544 39764 3596
rect 39816 3584 39822 3596
rect 40696 3584 40724 3624
rect 41601 3621 41613 3624
rect 41647 3621 41659 3655
rect 41601 3615 41659 3621
rect 41892 3593 41920 3692
rect 44821 3689 44833 3723
rect 44867 3720 44879 3723
rect 46934 3720 46940 3732
rect 44867 3692 46940 3720
rect 44867 3689 44879 3692
rect 44821 3683 44879 3689
rect 46934 3680 46940 3692
rect 46992 3680 46998 3732
rect 48774 3680 48780 3732
rect 48832 3720 48838 3732
rect 48869 3723 48927 3729
rect 48869 3720 48881 3723
rect 48832 3692 48881 3720
rect 48832 3680 48838 3692
rect 48869 3689 48881 3692
rect 48915 3689 48927 3723
rect 48869 3683 48927 3689
rect 67910 3680 67916 3732
rect 67968 3680 67974 3732
rect 71682 3680 71688 3732
rect 71740 3680 71746 3732
rect 77570 3680 77576 3732
rect 77628 3680 77634 3732
rect 46382 3652 46388 3664
rect 43916 3624 46388 3652
rect 39816 3556 40724 3584
rect 41325 3587 41383 3593
rect 39816 3544 39822 3556
rect 41325 3553 41337 3587
rect 41371 3553 41383 3587
rect 41325 3547 41383 3553
rect 41877 3587 41935 3593
rect 41877 3553 41889 3587
rect 41923 3553 41935 3587
rect 41877 3547 41935 3553
rect 40310 3476 40316 3528
rect 40368 3516 40374 3528
rect 41340 3516 41368 3547
rect 42242 3544 42248 3596
rect 42300 3544 42306 3596
rect 42521 3587 42579 3593
rect 42521 3553 42533 3587
rect 42567 3584 42579 3587
rect 43916 3584 43944 3624
rect 46382 3612 46388 3624
rect 46440 3612 46446 3664
rect 42567 3556 43944 3584
rect 43993 3587 44051 3593
rect 42567 3553 42579 3556
rect 42521 3547 42579 3553
rect 43993 3553 44005 3587
rect 44039 3553 44051 3587
rect 43993 3547 44051 3553
rect 41969 3519 42027 3525
rect 40368 3488 41414 3516
rect 40368 3476 40374 3488
rect 38804 3352 39712 3380
rect 38804 3340 38810 3352
rect 39942 3340 39948 3392
rect 40000 3380 40006 3392
rect 40773 3383 40831 3389
rect 40773 3380 40785 3383
rect 40000 3352 40785 3380
rect 40000 3340 40006 3352
rect 40773 3349 40785 3352
rect 40819 3349 40831 3383
rect 40773 3343 40831 3349
rect 41138 3340 41144 3392
rect 41196 3340 41202 3392
rect 41230 3340 41236 3392
rect 41288 3340 41294 3392
rect 41386 3380 41414 3488
rect 41969 3485 41981 3519
rect 42015 3516 42027 3519
rect 42058 3516 42064 3528
rect 42015 3488 42064 3516
rect 42015 3485 42027 3488
rect 41969 3479 42027 3485
rect 42058 3476 42064 3488
rect 42116 3476 42122 3528
rect 44008 3516 44036 3547
rect 44266 3544 44272 3596
rect 44324 3544 44330 3596
rect 44361 3587 44419 3593
rect 44361 3553 44373 3587
rect 44407 3584 44419 3587
rect 45554 3584 45560 3596
rect 44407 3556 45560 3584
rect 44407 3553 44419 3556
rect 44361 3547 44419 3553
rect 45554 3544 45560 3556
rect 45612 3544 45618 3596
rect 45738 3544 45744 3596
rect 45796 3584 45802 3596
rect 46753 3587 46811 3593
rect 46753 3584 46765 3587
rect 45796 3556 46765 3584
rect 45796 3544 45802 3556
rect 46753 3553 46765 3556
rect 46799 3553 46811 3587
rect 49973 3587 50031 3593
rect 49973 3584 49985 3587
rect 46753 3547 46811 3553
rect 46860 3556 49985 3584
rect 44453 3519 44511 3525
rect 44453 3516 44465 3519
rect 44008 3488 44465 3516
rect 44453 3485 44465 3488
rect 44499 3516 44511 3519
rect 45465 3519 45523 3525
rect 45465 3516 45477 3519
rect 44499 3488 45477 3516
rect 44499 3485 44511 3488
rect 44453 3479 44511 3485
rect 45465 3485 45477 3488
rect 45511 3485 45523 3519
rect 45465 3479 45523 3485
rect 45925 3519 45983 3525
rect 45925 3485 45937 3519
rect 45971 3516 45983 3519
rect 46290 3516 46296 3528
rect 45971 3488 46296 3516
rect 45971 3485 45983 3488
rect 45925 3479 45983 3485
rect 46290 3476 46296 3488
rect 46348 3476 46354 3528
rect 46474 3476 46480 3528
rect 46532 3476 46538 3528
rect 46658 3476 46664 3528
rect 46716 3516 46722 3528
rect 46860 3516 46888 3556
rect 49973 3553 49985 3556
rect 50019 3553 50031 3587
rect 49973 3547 50031 3553
rect 72418 3544 72424 3596
rect 72476 3544 72482 3596
rect 77018 3544 77024 3596
rect 77076 3544 77082 3596
rect 46716 3488 46888 3516
rect 46716 3476 46722 3488
rect 46934 3476 46940 3528
rect 46992 3516 46998 3528
rect 48317 3519 48375 3525
rect 48317 3516 48329 3519
rect 46992 3488 48329 3516
rect 46992 3476 46998 3488
rect 48317 3485 48329 3488
rect 48363 3485 48375 3519
rect 48317 3479 48375 3485
rect 49786 3476 49792 3528
rect 49844 3476 49850 3528
rect 51258 3476 51264 3528
rect 51316 3516 51322 3528
rect 52273 3519 52331 3525
rect 52273 3516 52285 3519
rect 51316 3488 52285 3516
rect 51316 3476 51322 3488
rect 52273 3485 52285 3488
rect 52319 3485 52331 3519
rect 52273 3479 52331 3485
rect 52454 3476 52460 3528
rect 52512 3476 52518 3528
rect 53650 3476 53656 3528
rect 53708 3476 53714 3528
rect 54297 3519 54355 3525
rect 54297 3485 54309 3519
rect 54343 3516 54355 3519
rect 54389 3519 54447 3525
rect 54389 3516 54401 3519
rect 54343 3488 54401 3516
rect 54343 3485 54355 3488
rect 54297 3479 54355 3485
rect 54389 3485 54401 3488
rect 54435 3485 54447 3519
rect 54389 3479 54447 3485
rect 57330 3476 57336 3528
rect 57388 3516 57394 3528
rect 57977 3519 58035 3525
rect 57977 3516 57989 3519
rect 57388 3488 57989 3516
rect 57388 3476 57394 3488
rect 57977 3485 57989 3488
rect 58023 3485 58035 3519
rect 57977 3479 58035 3485
rect 58066 3476 58072 3528
rect 58124 3516 58130 3528
rect 58161 3519 58219 3525
rect 58161 3516 58173 3519
rect 58124 3488 58173 3516
rect 58124 3476 58130 3488
rect 58161 3485 58173 3488
rect 58207 3485 58219 3519
rect 58161 3479 58219 3485
rect 60918 3476 60924 3528
rect 60976 3516 60982 3528
rect 61933 3519 61991 3525
rect 61933 3516 61945 3519
rect 60976 3488 61945 3516
rect 60976 3476 60982 3488
rect 61933 3485 61945 3488
rect 61979 3485 61991 3519
rect 61933 3479 61991 3485
rect 62114 3476 62120 3528
rect 62172 3476 62178 3528
rect 64690 3476 64696 3528
rect 64748 3516 64754 3528
rect 65705 3519 65763 3525
rect 65705 3516 65717 3519
rect 64748 3488 65717 3516
rect 64748 3476 64754 3488
rect 65705 3485 65717 3488
rect 65751 3485 65763 3519
rect 65705 3479 65763 3485
rect 67082 3476 67088 3528
rect 67140 3516 67146 3528
rect 67177 3519 67235 3525
rect 67177 3516 67189 3519
rect 67140 3488 67189 3516
rect 67140 3476 67146 3488
rect 67177 3485 67189 3488
rect 67223 3485 67235 3519
rect 67177 3479 67235 3485
rect 67821 3519 67879 3525
rect 67821 3485 67833 3519
rect 67867 3516 67879 3519
rect 68465 3519 68523 3525
rect 68465 3516 68477 3519
rect 67867 3488 68477 3516
rect 67867 3485 67879 3488
rect 67821 3479 67879 3485
rect 68465 3485 68477 3488
rect 68511 3485 68523 3519
rect 68465 3479 68523 3485
rect 69106 3476 69112 3528
rect 69164 3476 69170 3528
rect 69753 3519 69811 3525
rect 69753 3485 69765 3519
rect 69799 3516 69811 3519
rect 69845 3519 69903 3525
rect 69845 3516 69857 3519
rect 69799 3488 69857 3516
rect 69799 3485 69811 3488
rect 69753 3479 69811 3485
rect 69845 3485 69857 3488
rect 69891 3485 69903 3519
rect 69845 3479 69903 3485
rect 72234 3476 72240 3528
rect 72292 3476 72298 3528
rect 74442 3476 74448 3528
rect 74500 3516 74506 3528
rect 75089 3519 75147 3525
rect 75089 3516 75101 3519
rect 74500 3488 75101 3516
rect 74500 3476 74506 3488
rect 75089 3485 75101 3488
rect 75135 3485 75147 3519
rect 75089 3479 75147 3485
rect 76650 3476 76656 3528
rect 76708 3476 76714 3528
rect 41690 3408 41696 3460
rect 41748 3448 41754 3460
rect 42794 3448 42800 3460
rect 41748 3420 42800 3448
rect 41748 3408 41754 3420
rect 42794 3408 42800 3420
rect 42852 3408 42858 3460
rect 42978 3408 42984 3460
rect 43036 3408 43042 3460
rect 46842 3408 46848 3460
rect 46900 3448 46906 3460
rect 49237 3451 49295 3457
rect 49237 3448 49249 3451
rect 46900 3420 49249 3448
rect 46900 3408 46906 3420
rect 49237 3417 49249 3420
rect 49283 3417 49295 3451
rect 49237 3411 49295 3417
rect 75454 3408 75460 3460
rect 75512 3408 75518 3460
rect 44266 3380 44272 3392
rect 41386 3352 44272 3380
rect 44266 3340 44272 3352
rect 44324 3340 44330 3392
rect 44910 3340 44916 3392
rect 44968 3340 44974 3392
rect 46109 3383 46167 3389
rect 46109 3349 46121 3383
rect 46155 3380 46167 3383
rect 48590 3380 48596 3392
rect 46155 3352 48596 3380
rect 46155 3349 46167 3352
rect 46109 3343 46167 3349
rect 48590 3340 48596 3352
rect 48648 3340 48654 3392
rect 50614 3340 50620 3392
rect 50672 3340 50678 3392
rect 51442 3340 51448 3392
rect 51500 3380 51506 3392
rect 51721 3383 51779 3389
rect 51721 3380 51733 3383
rect 51500 3352 51733 3380
rect 51500 3340 51506 3352
rect 51721 3349 51733 3352
rect 51767 3349 51779 3383
rect 51721 3343 51779 3349
rect 53006 3340 53012 3392
rect 53064 3380 53070 3392
rect 53101 3383 53159 3389
rect 53101 3380 53113 3383
rect 53064 3352 53113 3380
rect 53064 3340 53070 3352
rect 53101 3349 53113 3352
rect 53147 3349 53159 3383
rect 53101 3343 53159 3349
rect 55033 3383 55091 3389
rect 55033 3349 55045 3383
rect 55079 3380 55091 3383
rect 56042 3380 56048 3392
rect 55079 3352 56048 3380
rect 55079 3349 55091 3352
rect 55033 3343 55091 3349
rect 56042 3340 56048 3352
rect 56100 3340 56106 3392
rect 57422 3340 57428 3392
rect 57480 3340 57486 3392
rect 58618 3340 58624 3392
rect 58676 3380 58682 3392
rect 58805 3383 58863 3389
rect 58805 3380 58817 3383
rect 58676 3352 58817 3380
rect 58676 3340 58682 3352
rect 58805 3349 58817 3352
rect 58851 3349 58863 3383
rect 58805 3343 58863 3349
rect 61102 3340 61108 3392
rect 61160 3380 61166 3392
rect 61381 3383 61439 3389
rect 61381 3380 61393 3383
rect 61160 3352 61393 3380
rect 61160 3340 61166 3352
rect 61381 3349 61393 3352
rect 61427 3349 61439 3383
rect 61381 3343 61439 3349
rect 62758 3340 62764 3392
rect 62816 3340 62822 3392
rect 64874 3340 64880 3392
rect 64932 3380 64938 3392
rect 65153 3383 65211 3389
rect 65153 3380 65165 3383
rect 64932 3352 65165 3380
rect 64932 3340 64938 3352
rect 65153 3349 65165 3352
rect 65199 3349 65211 3383
rect 65153 3343 65211 3349
rect 70489 3383 70547 3389
rect 70489 3349 70501 3383
rect 70535 3380 70547 3383
rect 71498 3380 71504 3392
rect 70535 3352 71504 3380
rect 70535 3349 70547 3352
rect 70489 3343 70547 3349
rect 71498 3340 71504 3352
rect 71556 3340 71562 3392
rect 73062 3340 73068 3392
rect 73120 3340 73126 3392
rect 74534 3340 74540 3392
rect 74592 3340 74598 3392
rect 2024 3290 77924 3312
rect 2024 3238 5794 3290
rect 5846 3238 5858 3290
rect 5910 3238 5922 3290
rect 5974 3238 5986 3290
rect 6038 3238 6050 3290
rect 6102 3238 36514 3290
rect 36566 3238 36578 3290
rect 36630 3238 36642 3290
rect 36694 3238 36706 3290
rect 36758 3238 36770 3290
rect 36822 3238 67234 3290
rect 67286 3238 67298 3290
rect 67350 3238 67362 3290
rect 67414 3238 67426 3290
rect 67478 3238 67490 3290
rect 67542 3238 77924 3290
rect 2024 3216 77924 3238
rect 4890 3136 4896 3188
rect 4948 3136 4954 3188
rect 6365 3179 6423 3185
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 7834 3176 7840 3188
rect 6411 3148 7840 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8205 3179 8263 3185
rect 8205 3145 8217 3179
rect 8251 3176 8263 3179
rect 9122 3176 9128 3188
rect 8251 3148 9128 3176
rect 8251 3145 8263 3148
rect 8205 3139 8263 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 9456 3148 10548 3176
rect 9456 3136 9462 3148
rect 6730 3068 6736 3120
rect 6788 3108 6794 3120
rect 10520 3108 10548 3148
rect 10594 3136 10600 3188
rect 10652 3176 10658 3188
rect 12158 3176 12164 3188
rect 10652 3148 12164 3176
rect 10652 3136 10658 3148
rect 12158 3136 12164 3148
rect 12216 3176 12222 3188
rect 12529 3179 12587 3185
rect 12216 3148 12434 3176
rect 12216 3136 12222 3148
rect 10781 3111 10839 3117
rect 10781 3108 10793 3111
rect 6788 3080 9904 3108
rect 10520 3080 10793 3108
rect 6788 3068 6794 3080
rect 4338 3000 4344 3052
rect 4396 3000 4402 3052
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 5534 3040 5540 3052
rect 5123 3012 5540 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 7006 3040 7012 3052
rect 6595 3012 7012 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 7101 3043 7159 3049
rect 7101 3009 7113 3043
rect 7147 3040 7159 3043
rect 8294 3040 8300 3052
rect 7147 3012 8300 3040
rect 7147 3009 7159 3012
rect 7101 3003 7159 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8386 3000 8392 3052
rect 8444 3000 8450 3052
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 9769 3043 9827 3049
rect 9769 3040 9781 3043
rect 9732 3012 9781 3040
rect 9732 3000 9738 3012
rect 9769 3009 9781 3012
rect 9815 3009 9827 3043
rect 9876 3040 9904 3080
rect 10781 3077 10793 3080
rect 10827 3077 10839 3111
rect 10781 3071 10839 3077
rect 11330 3068 11336 3120
rect 11388 3068 11394 3120
rect 12406 3108 12434 3148
rect 12529 3145 12541 3179
rect 12575 3176 12587 3179
rect 12894 3176 12900 3188
rect 12575 3148 12900 3176
rect 12575 3145 12587 3148
rect 12529 3139 12587 3145
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 15378 3176 15384 3188
rect 13096 3148 15384 3176
rect 13096 3108 13124 3148
rect 12406 3080 13124 3108
rect 10410 3040 10416 3052
rect 9876 3012 10416 3040
rect 9769 3003 9827 3009
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 10502 3000 10508 3052
rect 10560 3000 10566 3052
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 12897 3043 12955 3049
rect 12759 3012 12848 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 5813 2975 5871 2981
rect 5813 2941 5825 2975
rect 5859 2972 5871 2975
rect 7558 2972 7564 2984
rect 5859 2944 7564 2972
rect 5859 2941 5871 2944
rect 5813 2935 5871 2941
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 7653 2975 7711 2981
rect 7653 2941 7665 2975
rect 7699 2972 7711 2975
rect 8846 2972 8852 2984
rect 7699 2944 8852 2972
rect 7699 2941 7711 2944
rect 7653 2935 7711 2941
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 8941 2975 8999 2981
rect 8941 2941 8953 2975
rect 8987 2972 8999 2975
rect 11422 2972 11428 2984
rect 8987 2944 11428 2972
rect 8987 2941 8999 2944
rect 8941 2935 8999 2941
rect 11422 2932 11428 2944
rect 11480 2932 11486 2984
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 12253 2975 12311 2981
rect 12253 2972 12265 2975
rect 11572 2944 12265 2972
rect 11572 2932 11578 2944
rect 12253 2941 12265 2944
rect 12299 2941 12311 2975
rect 12253 2935 12311 2941
rect 5629 2907 5687 2913
rect 5629 2873 5641 2907
rect 5675 2904 5687 2907
rect 8018 2904 8024 2916
rect 5675 2876 8024 2904
rect 5675 2873 5687 2876
rect 5629 2867 5687 2873
rect 8018 2864 8024 2876
rect 8076 2864 8082 2916
rect 9677 2907 9735 2913
rect 9677 2873 9689 2907
rect 9723 2904 9735 2907
rect 10502 2904 10508 2916
rect 9723 2876 10508 2904
rect 9723 2873 9735 2876
rect 9677 2867 9735 2873
rect 10502 2864 10508 2876
rect 10560 2864 10566 2916
rect 7469 2839 7527 2845
rect 7469 2805 7481 2839
rect 7515 2836 7527 2839
rect 7650 2836 7656 2848
rect 7515 2808 7656 2836
rect 7515 2805 7527 2808
rect 7469 2799 7527 2805
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 10413 2839 10471 2845
rect 10413 2805 10425 2839
rect 10459 2836 10471 2839
rect 12710 2836 12716 2848
rect 10459 2808 12716 2836
rect 10459 2805 10471 2808
rect 10413 2799 10471 2805
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 12820 2836 12848 3012
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 12912 2972 12940 3003
rect 12986 3000 12992 3052
rect 13044 3000 13050 3052
rect 13096 3049 13124 3080
rect 13354 3068 13360 3120
rect 13412 3068 13418 3120
rect 13630 3068 13636 3120
rect 13688 3108 13694 3120
rect 13688 3080 13846 3108
rect 13688 3068 13694 3080
rect 14936 3049 14964 3148
rect 15378 3136 15384 3148
rect 15436 3176 15442 3188
rect 18138 3176 18144 3188
rect 15436 3148 18144 3176
rect 15436 3136 15442 3148
rect 18138 3136 18144 3148
rect 18196 3176 18202 3188
rect 19886 3176 19892 3188
rect 18196 3148 18368 3176
rect 18196 3136 18202 3148
rect 15654 3068 15660 3120
rect 15712 3068 15718 3120
rect 17405 3111 17463 3117
rect 17405 3077 17417 3111
rect 17451 3108 17463 3111
rect 17770 3108 17776 3120
rect 17451 3080 17776 3108
rect 17451 3077 17463 3080
rect 17405 3071 17463 3077
rect 17770 3068 17776 3080
rect 17828 3068 17834 3120
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3009 13139 3043
rect 13081 3003 13139 3009
rect 14921 3043 14979 3049
rect 14921 3009 14933 3043
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 16482 3000 16488 3052
rect 16540 3040 16546 3052
rect 18340 3049 18368 3148
rect 18984 3148 19892 3176
rect 18598 3068 18604 3120
rect 18656 3068 18662 3120
rect 18984 3108 19012 3148
rect 19886 3136 19892 3148
rect 19944 3136 19950 3188
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 20073 3179 20131 3185
rect 20073 3176 20085 3179
rect 20036 3148 20085 3176
rect 20036 3136 20042 3148
rect 20073 3145 20085 3148
rect 20119 3145 20131 3179
rect 20073 3139 20131 3145
rect 20162 3136 20168 3188
rect 20220 3176 20226 3188
rect 22951 3179 23009 3185
rect 20220 3148 22876 3176
rect 20220 3136 20226 3148
rect 19058 3108 19064 3120
rect 18984 3080 19064 3108
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 20180 3049 20208 3136
rect 21726 3108 21732 3120
rect 21666 3080 21732 3108
rect 21726 3068 21732 3080
rect 21784 3068 21790 3120
rect 22002 3068 22008 3120
rect 22060 3068 22066 3120
rect 22094 3068 22100 3120
rect 22152 3108 22158 3120
rect 22189 3111 22247 3117
rect 22189 3108 22201 3111
rect 22152 3080 22201 3108
rect 22152 3068 22158 3080
rect 22189 3077 22201 3080
rect 22235 3077 22247 3111
rect 22189 3071 22247 3077
rect 22370 3068 22376 3120
rect 22428 3068 22434 3120
rect 22738 3068 22744 3120
rect 22796 3068 22802 3120
rect 22848 3108 22876 3148
rect 22951 3145 22963 3179
rect 22997 3176 23009 3179
rect 23198 3176 23204 3188
rect 22997 3148 23204 3176
rect 22997 3145 23009 3148
rect 22951 3139 23009 3145
rect 23198 3136 23204 3148
rect 23256 3136 23262 3188
rect 25222 3176 25228 3188
rect 23584 3148 25228 3176
rect 23584 3120 23612 3148
rect 25222 3136 25228 3148
rect 25280 3176 25286 3188
rect 26602 3176 26608 3188
rect 25280 3148 26608 3176
rect 25280 3136 25286 3148
rect 26602 3136 26608 3148
rect 26660 3136 26666 3188
rect 26878 3136 26884 3188
rect 26936 3176 26942 3188
rect 27065 3179 27123 3185
rect 27065 3176 27077 3179
rect 26936 3148 27077 3176
rect 26936 3136 26942 3148
rect 27065 3145 27077 3148
rect 27111 3176 27123 3179
rect 27338 3176 27344 3188
rect 27111 3148 27344 3176
rect 27111 3145 27123 3148
rect 27065 3139 27123 3145
rect 27338 3136 27344 3148
rect 27396 3136 27402 3188
rect 28077 3179 28135 3185
rect 28077 3145 28089 3179
rect 28123 3176 28135 3179
rect 28166 3176 28172 3188
rect 28123 3148 28172 3176
rect 28123 3145 28135 3148
rect 28077 3139 28135 3145
rect 28166 3136 28172 3148
rect 28224 3136 28230 3188
rect 28258 3136 28264 3188
rect 28316 3176 28322 3188
rect 28537 3179 28595 3185
rect 28537 3176 28549 3179
rect 28316 3148 28549 3176
rect 28316 3136 28322 3148
rect 28537 3145 28549 3148
rect 28583 3145 28595 3179
rect 28537 3139 28595 3145
rect 30466 3136 30472 3188
rect 30524 3136 30530 3188
rect 32674 3136 32680 3188
rect 32732 3136 32738 3188
rect 33318 3136 33324 3188
rect 33376 3176 33382 3188
rect 33413 3179 33471 3185
rect 33413 3176 33425 3179
rect 33376 3148 33425 3176
rect 33376 3136 33382 3148
rect 33413 3145 33425 3148
rect 33459 3145 33471 3179
rect 33413 3139 33471 3145
rect 33502 3136 33508 3188
rect 33560 3136 33566 3188
rect 34054 3136 34060 3188
rect 34112 3136 34118 3188
rect 34149 3179 34207 3185
rect 34149 3145 34161 3179
rect 34195 3176 34207 3179
rect 34606 3176 34612 3188
rect 34195 3148 34612 3176
rect 34195 3145 34207 3148
rect 34149 3139 34207 3145
rect 34606 3136 34612 3148
rect 34664 3136 34670 3188
rect 35802 3176 35808 3188
rect 35544 3148 35808 3176
rect 23566 3108 23572 3120
rect 22848 3080 23572 3108
rect 18325 3043 18383 3049
rect 16540 3012 17724 3040
rect 16540 3000 16546 3012
rect 13446 2972 13452 2984
rect 12912 2944 13452 2972
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 15197 2975 15255 2981
rect 15197 2972 15209 2975
rect 13872 2944 15209 2972
rect 13872 2932 13878 2944
rect 15197 2941 15209 2944
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 16669 2975 16727 2981
rect 16669 2972 16681 2975
rect 15620 2944 16681 2972
rect 15620 2932 15626 2944
rect 16669 2941 16681 2944
rect 16715 2941 16727 2975
rect 16669 2935 16727 2941
rect 16853 2975 16911 2981
rect 16853 2941 16865 2975
rect 16899 2972 16911 2975
rect 16942 2972 16948 2984
rect 16899 2944 16948 2972
rect 16899 2941 16911 2944
rect 16853 2935 16911 2941
rect 16942 2932 16948 2944
rect 17000 2932 17006 2984
rect 17494 2932 17500 2984
rect 17552 2972 17558 2984
rect 17589 2975 17647 2981
rect 17589 2972 17601 2975
rect 17552 2944 17601 2972
rect 17552 2932 17558 2944
rect 17589 2941 17601 2944
rect 17635 2941 17647 2975
rect 17696 2972 17724 3012
rect 18325 3009 18337 3043
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3009 20223 3043
rect 20165 3003 20223 3009
rect 22278 3000 22284 3052
rect 22336 3000 22342 3052
rect 22557 3043 22615 3049
rect 22557 3009 22569 3043
rect 22603 3040 22615 3043
rect 23106 3040 23112 3052
rect 22603 3012 23112 3040
rect 22603 3009 22615 3012
rect 22557 3003 22615 3009
rect 23106 3000 23112 3012
rect 23164 3000 23170 3052
rect 23216 3049 23244 3080
rect 23566 3068 23572 3080
rect 23624 3068 23630 3120
rect 25866 3108 25872 3120
rect 24702 3094 25872 3108
rect 24688 3080 25872 3094
rect 24688 3074 24716 3080
rect 24596 3052 24716 3074
rect 25866 3068 25872 3080
rect 25924 3108 25930 3120
rect 25924 3080 26082 3108
rect 25924 3068 25930 3080
rect 27798 3068 27804 3120
rect 27856 3108 27862 3120
rect 28718 3108 28724 3120
rect 27856 3080 28724 3108
rect 27856 3068 27862 3080
rect 23201 3043 23259 3049
rect 23201 3009 23213 3043
rect 23247 3009 23259 3043
rect 23201 3003 23259 3009
rect 24578 3000 24584 3052
rect 24636 3046 24716 3052
rect 24636 3000 24642 3046
rect 25038 3000 25044 3052
rect 25096 3000 25102 3052
rect 25222 3000 25228 3052
rect 25280 3040 25286 3052
rect 25317 3043 25375 3049
rect 25317 3040 25329 3043
rect 25280 3012 25329 3040
rect 25280 3000 25286 3012
rect 25317 3009 25329 3012
rect 25363 3009 25375 3043
rect 25317 3003 25375 3009
rect 27246 3000 27252 3052
rect 27304 3000 27310 3052
rect 27338 3000 27344 3052
rect 27396 3000 27402 3052
rect 27525 3043 27583 3049
rect 27525 3009 27537 3043
rect 27571 3040 27583 3043
rect 27982 3040 27988 3052
rect 27571 3012 27988 3040
rect 27571 3009 27583 3012
rect 27525 3003 27583 3009
rect 27982 3000 27988 3012
rect 28040 3000 28046 3052
rect 28276 3049 28304 3080
rect 28718 3068 28724 3080
rect 28776 3068 28782 3120
rect 30006 3068 30012 3120
rect 30064 3068 30070 3120
rect 31110 3108 31116 3120
rect 30300 3080 30512 3108
rect 28169 3043 28227 3049
rect 28169 3009 28181 3043
rect 28215 3009 28227 3043
rect 28169 3003 28227 3009
rect 28261 3043 28319 3049
rect 28261 3009 28273 3043
rect 28307 3009 28319 3043
rect 28261 3003 28319 3009
rect 20441 2975 20499 2981
rect 20441 2972 20453 2975
rect 17696 2944 20453 2972
rect 17589 2935 17647 2941
rect 20441 2941 20453 2944
rect 20487 2941 20499 2975
rect 23477 2975 23535 2981
rect 23477 2972 23489 2975
rect 20441 2935 20499 2941
rect 22756 2944 23489 2972
rect 14550 2836 14556 2848
rect 12820 2808 14556 2836
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 14829 2839 14887 2845
rect 14829 2805 14841 2839
rect 14875 2836 14887 2839
rect 15286 2836 15292 2848
rect 14875 2808 15292 2836
rect 14875 2805 14887 2808
rect 14829 2799 14887 2805
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 16850 2796 16856 2848
rect 16908 2836 16914 2848
rect 17512 2836 17540 2932
rect 21450 2864 21456 2916
rect 21508 2904 21514 2916
rect 22756 2904 22784 2944
rect 23477 2941 23489 2944
rect 23523 2941 23535 2975
rect 23477 2935 23535 2941
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 25593 2975 25651 2981
rect 25593 2972 25605 2975
rect 23624 2944 25605 2972
rect 23624 2932 23630 2944
rect 25593 2941 25605 2944
rect 25639 2941 25651 2975
rect 25593 2935 25651 2941
rect 27154 2932 27160 2984
rect 27212 2972 27218 2984
rect 27433 2975 27491 2981
rect 27433 2972 27445 2975
rect 27212 2944 27445 2972
rect 27212 2932 27218 2944
rect 27433 2941 27445 2944
rect 27479 2941 27491 2975
rect 27433 2935 27491 2941
rect 27893 2975 27951 2981
rect 27893 2941 27905 2975
rect 27939 2972 27951 2975
rect 28074 2972 28080 2984
rect 27939 2944 28080 2972
rect 27939 2941 27951 2944
rect 27893 2935 27951 2941
rect 28074 2932 28080 2944
rect 28132 2932 28138 2984
rect 28184 2972 28212 3003
rect 28534 3000 28540 3052
rect 28592 3040 28598 3052
rect 30300 3049 30328 3080
rect 30285 3043 30343 3049
rect 28592 3012 28934 3040
rect 28592 3000 28598 3012
rect 30285 3009 30297 3043
rect 30331 3009 30343 3043
rect 30285 3003 30343 3009
rect 30377 3043 30435 3049
rect 30377 3009 30389 3043
rect 30423 3009 30435 3043
rect 30377 3003 30435 3009
rect 29270 2972 29276 2984
rect 28184 2944 29276 2972
rect 29270 2932 29276 2944
rect 29328 2932 29334 2984
rect 21508 2876 22784 2904
rect 21508 2864 21514 2876
rect 24670 2864 24676 2916
rect 24728 2904 24734 2916
rect 27709 2907 27767 2913
rect 27709 2904 27721 2907
rect 24728 2876 25452 2904
rect 24728 2864 24734 2876
rect 16908 2808 17540 2836
rect 18233 2839 18291 2845
rect 16908 2796 16914 2808
rect 18233 2805 18245 2839
rect 18279 2836 18291 2839
rect 20530 2836 20536 2848
rect 18279 2808 20536 2836
rect 18279 2805 18291 2808
rect 18233 2799 18291 2805
rect 20530 2796 20536 2808
rect 20588 2796 20594 2848
rect 21082 2796 21088 2848
rect 21140 2836 21146 2848
rect 21913 2839 21971 2845
rect 21913 2836 21925 2839
rect 21140 2808 21925 2836
rect 21140 2796 21146 2808
rect 21913 2805 21925 2808
rect 21959 2805 21971 2839
rect 21913 2799 21971 2805
rect 22922 2796 22928 2848
rect 22980 2796 22986 2848
rect 23109 2839 23167 2845
rect 23109 2805 23121 2839
rect 23155 2836 23167 2839
rect 24854 2836 24860 2848
rect 23155 2808 24860 2836
rect 23155 2805 23167 2808
rect 23109 2799 23167 2805
rect 24854 2796 24860 2808
rect 24912 2796 24918 2848
rect 24949 2839 25007 2845
rect 24949 2805 24961 2839
rect 24995 2836 25007 2839
rect 25130 2836 25136 2848
rect 24995 2808 25136 2836
rect 24995 2805 25007 2808
rect 24949 2799 25007 2805
rect 25130 2796 25136 2808
rect 25188 2796 25194 2848
rect 25222 2796 25228 2848
rect 25280 2796 25286 2848
rect 25424 2836 25452 2876
rect 26620 2876 27721 2904
rect 26620 2836 26648 2876
rect 27709 2873 27721 2876
rect 27755 2873 27767 2907
rect 30392 2904 30420 3003
rect 30484 2972 30512 3080
rect 30668 3080 31116 3108
rect 30668 3049 30696 3080
rect 31110 3068 31116 3080
rect 31168 3068 31174 3120
rect 31202 3068 31208 3120
rect 31260 3068 31266 3120
rect 32950 3108 32956 3120
rect 32430 3080 32956 3108
rect 32950 3068 32956 3080
rect 33008 3068 33014 3120
rect 33134 3068 33140 3120
rect 33192 3108 33198 3120
rect 35544 3108 35572 3148
rect 35802 3136 35808 3148
rect 35860 3136 35866 3188
rect 37826 3176 37832 3188
rect 35912 3148 37832 3176
rect 33192 3080 34100 3108
rect 35190 3080 35572 3108
rect 33192 3068 33198 3080
rect 30653 3043 30711 3049
rect 30653 3009 30665 3043
rect 30699 3009 30711 3043
rect 33778 3040 33784 3052
rect 30653 3003 30711 3009
rect 32508 3012 33784 3040
rect 30929 2975 30987 2981
rect 30929 2972 30941 2975
rect 30484 2944 30941 2972
rect 30929 2941 30941 2944
rect 30975 2972 30987 2975
rect 31294 2972 31300 2984
rect 30975 2944 31300 2972
rect 30975 2941 30987 2944
rect 30929 2935 30987 2941
rect 31294 2932 31300 2944
rect 31352 2932 31358 2984
rect 32214 2932 32220 2984
rect 32272 2972 32278 2984
rect 32508 2972 32536 3012
rect 33612 2981 33640 3012
rect 33778 3000 33784 3012
rect 33836 3000 33842 3052
rect 33870 3000 33876 3052
rect 33928 3000 33934 3052
rect 34072 3049 34100 3080
rect 35618 3068 35624 3120
rect 35676 3068 35682 3120
rect 35912 3049 35940 3148
rect 37826 3136 37832 3148
rect 37884 3176 37890 3188
rect 38381 3179 38439 3185
rect 37884 3148 37964 3176
rect 37884 3136 37890 3148
rect 37550 3108 37556 3120
rect 37214 3080 37556 3108
rect 37550 3068 37556 3080
rect 37608 3068 37614 3120
rect 37642 3068 37648 3120
rect 37700 3068 37706 3120
rect 37936 3108 37964 3148
rect 38381 3145 38393 3179
rect 38427 3176 38439 3179
rect 38470 3176 38476 3188
rect 38427 3148 38476 3176
rect 38427 3145 38439 3148
rect 38381 3139 38439 3145
rect 38470 3136 38476 3148
rect 38528 3136 38534 3188
rect 40405 3179 40463 3185
rect 38672 3148 40264 3176
rect 38672 3108 38700 3148
rect 37936 3080 38700 3108
rect 40236 3108 40264 3148
rect 40405 3145 40417 3179
rect 40451 3176 40463 3179
rect 41138 3176 41144 3188
rect 40451 3148 41144 3176
rect 40451 3145 40463 3148
rect 40405 3139 40463 3145
rect 41138 3136 41144 3148
rect 41196 3136 41202 3188
rect 41325 3179 41383 3185
rect 41325 3145 41337 3179
rect 41371 3176 41383 3179
rect 41690 3176 41696 3188
rect 41371 3148 41696 3176
rect 41371 3145 41383 3148
rect 41325 3139 41383 3145
rect 41690 3136 41696 3148
rect 41748 3136 41754 3188
rect 42334 3176 42340 3188
rect 41800 3148 42340 3176
rect 41800 3108 41828 3148
rect 42334 3136 42340 3148
rect 42392 3136 42398 3188
rect 43165 3179 43223 3185
rect 43165 3145 43177 3179
rect 43211 3176 43223 3179
rect 44818 3176 44824 3188
rect 43211 3148 44824 3176
rect 43211 3145 43223 3148
rect 43165 3139 43223 3145
rect 44818 3136 44824 3148
rect 44876 3136 44882 3188
rect 45370 3136 45376 3188
rect 45428 3136 45434 3188
rect 45649 3179 45707 3185
rect 45649 3145 45661 3179
rect 45695 3176 45707 3179
rect 45922 3176 45928 3188
rect 45695 3148 45928 3176
rect 45695 3145 45707 3148
rect 45649 3139 45707 3145
rect 45922 3136 45928 3148
rect 45980 3136 45986 3188
rect 48038 3136 48044 3188
rect 48096 3136 48102 3188
rect 50062 3136 50068 3188
rect 50120 3136 50126 3188
rect 51258 3136 51264 3188
rect 51316 3136 51322 3188
rect 51997 3179 52055 3185
rect 51997 3145 52009 3179
rect 52043 3176 52055 3179
rect 52454 3176 52460 3188
rect 52043 3148 52460 3176
rect 52043 3145 52055 3148
rect 51997 3139 52055 3145
rect 52454 3136 52460 3148
rect 52512 3136 52518 3188
rect 53650 3136 53656 3188
rect 53708 3136 53714 3188
rect 57330 3136 57336 3188
rect 57388 3136 57394 3188
rect 58066 3136 58072 3188
rect 58124 3136 58130 3188
rect 60918 3136 60924 3188
rect 60976 3136 60982 3188
rect 61657 3179 61715 3185
rect 61657 3145 61669 3179
rect 61703 3176 61715 3179
rect 62114 3176 62120 3188
rect 61703 3148 62120 3176
rect 61703 3145 61715 3148
rect 61657 3139 61715 3145
rect 62114 3136 62120 3148
rect 62172 3136 62178 3188
rect 64690 3136 64696 3188
rect 64748 3136 64754 3188
rect 65426 3136 65432 3188
rect 65484 3136 65490 3188
rect 67082 3136 67088 3188
rect 67140 3176 67146 3188
rect 67177 3179 67235 3185
rect 67177 3176 67189 3179
rect 67140 3148 67189 3176
rect 67140 3136 67146 3148
rect 67177 3145 67189 3148
rect 67223 3145 67235 3179
rect 67177 3139 67235 3145
rect 69106 3136 69112 3188
rect 69164 3136 69170 3188
rect 74442 3136 74448 3188
rect 74500 3136 74506 3188
rect 42978 3108 42984 3120
rect 40236 3080 41828 3108
rect 42918 3080 42984 3108
rect 34057 3043 34115 3049
rect 34057 3009 34069 3043
rect 34103 3009 34115 3043
rect 34057 3003 34115 3009
rect 35897 3043 35955 3049
rect 35897 3009 35909 3043
rect 35943 3009 35955 3043
rect 35897 3003 35955 3009
rect 35986 3000 35992 3052
rect 36044 3040 36050 3052
rect 36081 3043 36139 3049
rect 36081 3040 36093 3043
rect 36044 3012 36093 3040
rect 36044 3000 36050 3012
rect 36081 3009 36093 3012
rect 36127 3040 36139 3043
rect 36262 3040 36268 3052
rect 36127 3012 36268 3040
rect 36127 3009 36139 3012
rect 36081 3003 36139 3009
rect 36262 3000 36268 3012
rect 36320 3000 36326 3052
rect 37936 3049 37964 3080
rect 38672 3049 38700 3080
rect 37921 3043 37979 3049
rect 37921 3009 37933 3043
rect 37967 3009 37979 3043
rect 37921 3003 37979 3009
rect 38197 3043 38255 3049
rect 38197 3009 38209 3043
rect 38243 3009 38255 3043
rect 38197 3003 38255 3009
rect 38657 3043 38715 3049
rect 38657 3009 38669 3043
rect 38703 3009 38715 3043
rect 38657 3003 38715 3009
rect 33597 2975 33655 2981
rect 32272 2944 32536 2972
rect 32600 2944 33180 2972
rect 32272 2932 32278 2944
rect 30392 2876 31064 2904
rect 27709 2867 27767 2873
rect 25424 2808 26648 2836
rect 28445 2839 28503 2845
rect 28445 2805 28457 2839
rect 28491 2836 28503 2839
rect 29914 2836 29920 2848
rect 28491 2808 29920 2836
rect 28491 2805 28503 2808
rect 28445 2799 28503 2805
rect 29914 2796 29920 2808
rect 29972 2796 29978 2848
rect 30374 2796 30380 2848
rect 30432 2836 30438 2848
rect 30558 2836 30564 2848
rect 30432 2808 30564 2836
rect 30432 2796 30438 2808
rect 30558 2796 30564 2808
rect 30616 2796 30622 2848
rect 30834 2796 30840 2848
rect 30892 2796 30898 2848
rect 31036 2836 31064 2876
rect 32600 2836 32628 2944
rect 33042 2864 33048 2916
rect 33100 2864 33106 2916
rect 33152 2904 33180 2944
rect 33597 2941 33609 2975
rect 33643 2941 33655 2975
rect 33597 2935 33655 2941
rect 34606 2932 34612 2984
rect 34664 2972 34670 2984
rect 38212 2972 38240 3003
rect 40034 3000 40040 3052
rect 40092 3000 40098 3052
rect 40954 3000 40960 3052
rect 41012 3000 41018 3052
rect 41432 3049 41460 3080
rect 42978 3068 42984 3080
rect 43036 3068 43042 3120
rect 43806 3068 43812 3120
rect 43864 3068 43870 3120
rect 45094 3068 45100 3120
rect 45152 3108 45158 3120
rect 46934 3108 46940 3120
rect 45152 3080 46940 3108
rect 45152 3068 45158 3080
rect 46934 3068 46940 3080
rect 46992 3068 46998 3120
rect 70302 3108 70308 3120
rect 53852 3080 70308 3108
rect 41406 3043 41464 3049
rect 41406 3009 41418 3043
rect 41452 3009 41464 3043
rect 41406 3003 41464 3009
rect 43346 3000 43352 3052
rect 43404 3040 43410 3052
rect 43533 3043 43591 3049
rect 43533 3040 43545 3043
rect 43404 3012 43545 3040
rect 43404 3000 43410 3012
rect 43533 3009 43545 3012
rect 43579 3009 43591 3043
rect 43901 3043 43959 3049
rect 43901 3040 43913 3043
rect 43533 3003 43591 3009
rect 43640 3012 43913 3040
rect 34664 2944 38240 2972
rect 34664 2932 34670 2944
rect 38378 2932 38384 2984
rect 38436 2972 38442 2984
rect 38933 2975 38991 2981
rect 38933 2972 38945 2975
rect 38436 2944 38945 2972
rect 38436 2932 38442 2944
rect 38933 2941 38945 2944
rect 38979 2941 38991 2975
rect 38933 2935 38991 2941
rect 40310 2932 40316 2984
rect 40368 2972 40374 2984
rect 40681 2975 40739 2981
rect 40681 2972 40693 2975
rect 40368 2944 40693 2972
rect 40368 2932 40374 2944
rect 40681 2941 40693 2944
rect 40727 2941 40739 2975
rect 40681 2935 40739 2941
rect 40865 2975 40923 2981
rect 40865 2941 40877 2975
rect 40911 2972 40923 2975
rect 41693 2975 41751 2981
rect 40911 2944 41414 2972
rect 40911 2941 40923 2944
rect 40865 2935 40923 2941
rect 41386 2916 41414 2944
rect 41693 2941 41705 2975
rect 41739 2972 41751 2975
rect 42150 2972 42156 2984
rect 41739 2944 42156 2972
rect 41739 2941 41751 2944
rect 41693 2935 41751 2941
rect 42150 2932 42156 2944
rect 42208 2932 42214 2984
rect 43640 2972 43668 3012
rect 43901 3009 43913 3012
rect 43947 3009 43959 3043
rect 43901 3003 43959 3009
rect 45557 3043 45615 3049
rect 45557 3009 45569 3043
rect 45603 3040 45615 3043
rect 45646 3040 45652 3052
rect 45603 3012 45652 3040
rect 45603 3009 45615 3012
rect 45557 3003 45615 3009
rect 45646 3000 45652 3012
rect 45704 3000 45710 3052
rect 45830 3000 45836 3052
rect 45888 3000 45894 3052
rect 46106 3000 46112 3052
rect 46164 3000 46170 3052
rect 47486 3000 47492 3052
rect 47544 3000 47550 3052
rect 48317 3043 48375 3049
rect 48317 3009 48329 3043
rect 48363 3040 48375 3043
rect 49234 3040 49240 3052
rect 48363 3012 49240 3040
rect 48363 3009 48375 3012
rect 48317 3003 48375 3009
rect 49234 3000 49240 3012
rect 49292 3000 49298 3052
rect 49786 3000 49792 3052
rect 49844 3000 49850 3052
rect 50614 3000 50620 3052
rect 50672 3000 50678 3052
rect 51074 3000 51080 3052
rect 51132 3000 51138 3052
rect 51442 3000 51448 3052
rect 51500 3000 51506 3052
rect 52086 3000 52092 3052
rect 52144 3000 52150 3052
rect 52362 3000 52368 3052
rect 52420 3040 52426 3052
rect 53852 3049 53880 3080
rect 53837 3043 53895 3049
rect 53837 3040 53849 3043
rect 52420 3012 53849 3040
rect 52420 3000 52426 3012
rect 53837 3009 53849 3012
rect 53883 3009 53895 3043
rect 53837 3003 53895 3009
rect 54018 3000 54024 3052
rect 54076 3000 54082 3052
rect 56042 3000 56048 3052
rect 56100 3000 56106 3052
rect 57164 3049 57192 3080
rect 57149 3043 57207 3049
rect 57149 3009 57161 3043
rect 57195 3009 57207 3043
rect 57149 3003 57207 3009
rect 57422 3000 57428 3052
rect 57480 3000 57486 3052
rect 60752 3049 60780 3080
rect 60737 3043 60795 3049
rect 60737 3009 60749 3043
rect 60783 3009 60795 3043
rect 60737 3003 60795 3009
rect 61102 3000 61108 3052
rect 61160 3000 61166 3052
rect 61746 3000 61752 3052
rect 61804 3000 61810 3052
rect 64524 3049 64552 3080
rect 64509 3043 64567 3049
rect 64509 3009 64521 3043
rect 64555 3009 64567 3043
rect 64509 3003 64567 3009
rect 64874 3000 64880 3052
rect 64932 3000 64938 3052
rect 65518 3000 65524 3052
rect 65576 3000 65582 3052
rect 67008 3049 67036 3080
rect 66993 3043 67051 3049
rect 66993 3009 67005 3043
rect 67039 3009 67051 3043
rect 66993 3003 67051 3009
rect 67634 3000 67640 3052
rect 67692 3000 67698 3052
rect 69308 3049 69336 3080
rect 70302 3068 70308 3080
rect 70360 3068 70366 3120
rect 69293 3043 69351 3049
rect 69293 3009 69305 3043
rect 69339 3009 69351 3043
rect 69293 3003 69351 3009
rect 69474 3000 69480 3052
rect 69532 3000 69538 3052
rect 71498 3000 71504 3052
rect 71556 3000 71562 3052
rect 72602 3000 72608 3052
rect 72660 3040 72666 3052
rect 72973 3043 73031 3049
rect 72973 3040 72985 3043
rect 72660 3012 72985 3040
rect 72660 3000 72666 3012
rect 72973 3009 72985 3012
rect 73019 3009 73031 3043
rect 72973 3003 73031 3009
rect 74074 3000 74080 3052
rect 74132 3040 74138 3052
rect 74261 3043 74319 3049
rect 74261 3040 74273 3043
rect 74132 3012 74273 3040
rect 74132 3000 74138 3012
rect 74261 3009 74273 3012
rect 74307 3009 74319 3043
rect 74261 3003 74319 3009
rect 74534 3000 74540 3052
rect 74592 3000 74598 3052
rect 76650 3000 76656 3052
rect 76708 3000 76714 3052
rect 42720 2944 43668 2972
rect 43717 2975 43775 2981
rect 34422 2904 34428 2916
rect 33152 2876 34428 2904
rect 34422 2864 34428 2876
rect 34480 2864 34486 2916
rect 35912 2876 36676 2904
rect 41386 2876 41420 2916
rect 31036 2808 32628 2836
rect 34882 2796 34888 2848
rect 34940 2836 34946 2848
rect 35066 2836 35072 2848
rect 34940 2808 35072 2836
rect 34940 2796 34946 2808
rect 35066 2796 35072 2808
rect 35124 2796 35130 2848
rect 35526 2796 35532 2848
rect 35584 2836 35590 2848
rect 35912 2836 35940 2876
rect 35584 2808 35940 2836
rect 35584 2796 35590 2808
rect 36170 2796 36176 2848
rect 36228 2796 36234 2848
rect 36648 2836 36676 2876
rect 41414 2864 41420 2876
rect 41472 2864 41478 2916
rect 42720 2836 42748 2944
rect 43717 2941 43729 2975
rect 43763 2972 43775 2975
rect 44910 2972 44916 2984
rect 43763 2944 44916 2972
rect 43763 2941 43775 2944
rect 43717 2935 43775 2941
rect 44910 2932 44916 2944
rect 44968 2932 44974 2984
rect 45097 2975 45155 2981
rect 45097 2941 45109 2975
rect 45143 2972 45155 2975
rect 45922 2972 45928 2984
rect 45143 2944 45928 2972
rect 45143 2941 45155 2944
rect 45097 2935 45155 2941
rect 45922 2932 45928 2944
rect 45980 2932 45986 2984
rect 46474 2932 46480 2984
rect 46532 2932 46538 2984
rect 47670 2932 47676 2984
rect 47728 2972 47734 2984
rect 48777 2975 48835 2981
rect 48777 2972 48789 2975
rect 47728 2944 48789 2972
rect 47728 2932 47734 2944
rect 48777 2941 48789 2944
rect 48823 2941 48835 2975
rect 48777 2935 48835 2941
rect 51534 2932 51540 2984
rect 51592 2972 51598 2984
rect 52549 2975 52607 2981
rect 52549 2972 52561 2975
rect 51592 2944 52561 2972
rect 51592 2932 51598 2944
rect 52549 2941 52561 2944
rect 52595 2941 52607 2975
rect 52549 2935 52607 2941
rect 53466 2932 53472 2984
rect 53524 2972 53530 2984
rect 54481 2975 54539 2981
rect 54481 2972 54493 2975
rect 53524 2944 54493 2972
rect 53524 2932 53530 2944
rect 54481 2941 54493 2944
rect 54527 2941 54539 2975
rect 54481 2935 54539 2941
rect 61194 2932 61200 2984
rect 61252 2972 61258 2984
rect 62209 2975 62267 2981
rect 62209 2972 62221 2975
rect 61252 2944 62221 2972
rect 61252 2932 61258 2944
rect 62209 2941 62221 2944
rect 62255 2941 62267 2975
rect 62209 2935 62267 2941
rect 65058 2932 65064 2984
rect 65116 2972 65122 2984
rect 65981 2975 66039 2981
rect 65981 2972 65993 2975
rect 65116 2944 65993 2972
rect 65116 2932 65122 2944
rect 65981 2941 65993 2944
rect 66027 2941 66039 2975
rect 68005 2975 68063 2981
rect 68005 2972 68017 2975
rect 65981 2935 66039 2941
rect 67008 2944 68017 2972
rect 67008 2916 67036 2944
rect 68005 2941 68017 2944
rect 68051 2941 68063 2975
rect 68005 2935 68063 2941
rect 68922 2932 68928 2984
rect 68980 2972 68986 2984
rect 69937 2975 69995 2981
rect 69937 2972 69949 2975
rect 68980 2944 69949 2972
rect 68980 2932 68986 2944
rect 69937 2941 69949 2944
rect 69983 2941 69995 2975
rect 69937 2935 69995 2941
rect 70854 2932 70860 2984
rect 70912 2972 70918 2984
rect 71961 2975 72019 2981
rect 71961 2972 71973 2975
rect 70912 2944 71973 2972
rect 70912 2932 70918 2944
rect 71961 2941 71973 2944
rect 72007 2941 72019 2975
rect 71961 2935 72019 2941
rect 74718 2932 74724 2984
rect 74776 2972 74782 2984
rect 75457 2975 75515 2981
rect 75457 2972 75469 2975
rect 74776 2944 75469 2972
rect 74776 2932 74782 2944
rect 75457 2941 75469 2944
rect 75503 2941 75515 2975
rect 75457 2935 75515 2941
rect 77297 2975 77355 2981
rect 77297 2941 77309 2975
rect 77343 2941 77355 2975
rect 77297 2935 77355 2941
rect 45462 2864 45468 2916
rect 45520 2904 45526 2916
rect 48133 2907 48191 2913
rect 48133 2904 48145 2907
rect 45520 2876 48145 2904
rect 45520 2864 45526 2876
rect 48133 2873 48145 2876
rect 48179 2873 48191 2907
rect 48133 2867 48191 2873
rect 66990 2864 66996 2916
rect 67048 2864 67054 2916
rect 75181 2907 75239 2913
rect 75181 2873 75193 2907
rect 75227 2904 75239 2907
rect 77312 2904 77340 2935
rect 75227 2876 77340 2904
rect 75227 2873 75239 2876
rect 75181 2867 75239 2873
rect 36648 2808 42748 2836
rect 42794 2796 42800 2848
rect 42852 2836 42858 2848
rect 43349 2839 43407 2845
rect 43349 2836 43361 2839
rect 42852 2808 43361 2836
rect 42852 2796 42858 2808
rect 43349 2805 43361 2808
rect 43395 2805 43407 2839
rect 43349 2799 43407 2805
rect 43530 2796 43536 2848
rect 43588 2796 43594 2848
rect 55306 2796 55312 2848
rect 55364 2836 55370 2848
rect 55493 2839 55551 2845
rect 55493 2836 55505 2839
rect 55364 2808 55505 2836
rect 55364 2796 55370 2808
rect 55493 2805 55505 2808
rect 55539 2805 55551 2839
rect 55493 2799 55551 2805
rect 59262 2796 59268 2848
rect 59320 2836 59326 2848
rect 59357 2839 59415 2845
rect 59357 2836 59369 2839
rect 59320 2808 59369 2836
rect 59320 2796 59326 2808
rect 59357 2805 59369 2808
rect 59403 2805 59415 2839
rect 59357 2799 59415 2805
rect 70486 2796 70492 2848
rect 70544 2836 70550 2848
rect 70949 2839 71007 2845
rect 70949 2836 70961 2839
rect 70544 2808 70961 2836
rect 70544 2796 70550 2808
rect 70949 2805 70961 2808
rect 70995 2805 71007 2839
rect 70949 2799 71007 2805
rect 76190 2796 76196 2848
rect 76248 2836 76254 2848
rect 76745 2839 76803 2845
rect 76745 2836 76757 2839
rect 76248 2808 76757 2836
rect 76248 2796 76254 2808
rect 76745 2805 76757 2808
rect 76791 2805 76803 2839
rect 76745 2799 76803 2805
rect 2024 2746 77924 2768
rect 2024 2694 5134 2746
rect 5186 2694 5198 2746
rect 5250 2694 5262 2746
rect 5314 2694 5326 2746
rect 5378 2694 5390 2746
rect 5442 2694 35854 2746
rect 35906 2694 35918 2746
rect 35970 2694 35982 2746
rect 36034 2694 36046 2746
rect 36098 2694 36110 2746
rect 36162 2694 66574 2746
rect 66626 2694 66638 2746
rect 66690 2694 66702 2746
rect 66754 2694 66766 2746
rect 66818 2694 66830 2746
rect 66882 2694 77924 2746
rect 2024 2672 77924 2694
rect 3786 2592 3792 2644
rect 3844 2592 3850 2644
rect 4522 2592 4528 2644
rect 4580 2592 4586 2644
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5626 2632 5632 2644
rect 4939 2604 5632 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6362 2592 6368 2644
rect 6420 2592 6426 2644
rect 8205 2635 8263 2641
rect 8205 2601 8217 2635
rect 8251 2632 8263 2635
rect 9766 2632 9772 2644
rect 8251 2604 9772 2632
rect 8251 2601 8263 2604
rect 8205 2595 8263 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10042 2592 10048 2644
rect 10100 2592 10106 2644
rect 12437 2635 12495 2641
rect 12437 2632 12449 2635
rect 10152 2604 12449 2632
rect 8846 2524 8852 2576
rect 8904 2564 8910 2576
rect 10152 2564 10180 2604
rect 12437 2601 12449 2604
rect 12483 2601 12495 2635
rect 12437 2595 12495 2601
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 15105 2635 15163 2641
rect 12768 2604 15056 2632
rect 12768 2592 12774 2604
rect 8904 2536 10180 2564
rect 8904 2524 8910 2536
rect 11238 2524 11244 2576
rect 11296 2524 11302 2576
rect 13906 2564 13912 2576
rect 12544 2536 13912 2564
rect 3970 2456 3976 2508
rect 4028 2456 4034 2508
rect 5810 2456 5816 2508
rect 5868 2456 5874 2508
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 7926 2496 7932 2508
rect 6595 2468 7932 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 9677 2499 9735 2505
rect 9677 2465 9689 2499
rect 9723 2496 9735 2499
rect 10778 2496 10784 2508
rect 9723 2468 10784 2496
rect 9723 2465 9735 2468
rect 9677 2459 9735 2465
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 11790 2496 11796 2508
rect 11112 2468 11796 2496
rect 11112 2456 11118 2468
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 3602 2388 3608 2440
rect 3660 2388 3666 2440
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 6178 2428 6184 2440
rect 5123 2400 6184 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 6178 2388 6184 2400
rect 6236 2388 6242 2440
rect 7650 2388 7656 2440
rect 7708 2388 7714 2440
rect 8386 2388 8392 2440
rect 8444 2388 8450 2440
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2428 10379 2431
rect 10410 2428 10416 2440
rect 10367 2400 10416 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 10594 2388 10600 2440
rect 10652 2388 10658 2440
rect 11514 2388 11520 2440
rect 11572 2428 11578 2440
rect 11609 2431 11667 2437
rect 11609 2428 11621 2431
rect 11572 2400 11621 2428
rect 11572 2388 11578 2400
rect 11609 2397 11621 2400
rect 11655 2397 11667 2431
rect 11609 2391 11667 2397
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2428 12311 2431
rect 12544 2428 12572 2536
rect 13906 2524 13912 2536
rect 13964 2524 13970 2576
rect 15028 2564 15056 2604
rect 15105 2601 15117 2635
rect 15151 2632 15163 2635
rect 16850 2632 16856 2644
rect 15151 2604 16856 2632
rect 15151 2601 15163 2604
rect 15105 2595 15163 2601
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17126 2592 17132 2644
rect 17184 2632 17190 2644
rect 17589 2635 17647 2641
rect 17589 2632 17601 2635
rect 17184 2604 17601 2632
rect 17184 2592 17190 2604
rect 17589 2601 17601 2604
rect 17635 2601 17647 2635
rect 20254 2632 20260 2644
rect 17589 2595 17647 2601
rect 18156 2604 20260 2632
rect 15028 2536 15976 2564
rect 12618 2456 12624 2508
rect 12676 2496 12682 2508
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12676 2468 12909 2496
rect 12676 2456 12682 2468
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2496 13139 2499
rect 13127 2468 14780 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 12299 2400 12572 2428
rect 12299 2397 12311 2400
rect 12253 2391 12311 2397
rect 12802 2388 12808 2440
rect 12860 2388 12866 2440
rect 5626 2320 5632 2372
rect 5684 2320 5690 2372
rect 7469 2363 7527 2369
rect 7469 2329 7481 2363
rect 7515 2360 7527 2363
rect 8404 2360 8432 2388
rect 10962 2360 10968 2372
rect 7515 2332 8432 2360
rect 8864 2332 10968 2360
rect 7515 2329 7527 2332
rect 7469 2323 7527 2329
rect 7101 2295 7159 2301
rect 7101 2261 7113 2295
rect 7147 2292 7159 2295
rect 8864 2292 8892 2332
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 11149 2363 11207 2369
rect 11149 2329 11161 2363
rect 11195 2360 11207 2363
rect 12986 2360 12992 2372
rect 11195 2332 12992 2360
rect 11195 2329 11207 2332
rect 11149 2323 11207 2329
rect 12986 2320 12992 2332
rect 13044 2320 13050 2372
rect 7147 2264 8892 2292
rect 7147 2261 7159 2264
rect 7101 2255 7159 2261
rect 8938 2252 8944 2304
rect 8996 2252 9002 2304
rect 11698 2252 11704 2304
rect 11756 2252 11762 2304
rect 11790 2252 11796 2304
rect 11848 2292 11854 2304
rect 13096 2292 13124 2459
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2428 13415 2431
rect 13403 2400 14596 2428
rect 13403 2397 13415 2400
rect 13357 2391 13415 2397
rect 13538 2320 13544 2372
rect 13596 2360 13602 2372
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 13596 2332 13645 2360
rect 13596 2320 13602 2332
rect 13633 2329 13645 2332
rect 13679 2329 13691 2363
rect 14568 2360 14596 2400
rect 14642 2388 14648 2440
rect 14700 2388 14706 2440
rect 14752 2428 14780 2468
rect 14826 2456 14832 2508
rect 14884 2496 14890 2508
rect 15657 2499 15715 2505
rect 15657 2496 15669 2499
rect 14884 2468 15669 2496
rect 14884 2456 14890 2468
rect 15657 2465 15669 2468
rect 15703 2465 15715 2499
rect 15657 2459 15715 2465
rect 15841 2499 15899 2505
rect 15841 2465 15853 2499
rect 15887 2465 15899 2499
rect 15948 2496 15976 2536
rect 16022 2524 16028 2576
rect 16080 2564 16086 2576
rect 18156 2564 18184 2604
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 21361 2635 21419 2641
rect 21361 2601 21373 2635
rect 21407 2632 21419 2635
rect 24302 2632 24308 2644
rect 21407 2604 24308 2632
rect 21407 2601 21419 2604
rect 21361 2595 21419 2601
rect 24302 2592 24308 2604
rect 24360 2592 24366 2644
rect 26510 2632 26516 2644
rect 25056 2604 26516 2632
rect 16080 2536 18184 2564
rect 16080 2524 16086 2536
rect 18156 2505 18184 2536
rect 18509 2567 18567 2573
rect 18509 2533 18521 2567
rect 18555 2564 18567 2567
rect 23661 2567 23719 2573
rect 18555 2536 20760 2564
rect 18555 2533 18567 2536
rect 18509 2527 18567 2533
rect 20732 2508 20760 2536
rect 23661 2533 23673 2567
rect 23707 2564 23719 2567
rect 25056 2564 25084 2604
rect 26510 2592 26516 2604
rect 26568 2592 26574 2644
rect 33965 2635 34023 2641
rect 33965 2601 33977 2635
rect 34011 2632 34023 2635
rect 34606 2632 34612 2644
rect 34011 2604 34612 2632
rect 34011 2601 34023 2604
rect 33965 2595 34023 2601
rect 34606 2592 34612 2604
rect 34664 2592 34670 2644
rect 41598 2632 41604 2644
rect 36464 2604 41604 2632
rect 23707 2536 25084 2564
rect 25501 2567 25559 2573
rect 23707 2533 23719 2536
rect 23661 2527 23719 2533
rect 25501 2533 25513 2567
rect 25547 2564 25559 2567
rect 30653 2567 30711 2573
rect 30653 2564 30665 2567
rect 25547 2536 25636 2564
rect 25547 2533 25559 2536
rect 25501 2527 25559 2533
rect 18141 2499 18199 2505
rect 15948 2468 16068 2496
rect 15841 2459 15899 2465
rect 14752 2424 15700 2428
rect 15746 2424 15752 2440
rect 14752 2400 15752 2424
rect 15672 2396 15752 2400
rect 15746 2388 15752 2396
rect 15804 2428 15810 2440
rect 15856 2428 15884 2459
rect 16040 2437 16068 2468
rect 18141 2465 18153 2499
rect 18187 2465 18199 2499
rect 18141 2459 18199 2465
rect 19334 2456 19340 2508
rect 19392 2456 19398 2508
rect 20714 2456 20720 2508
rect 20772 2456 20778 2508
rect 22186 2456 22192 2508
rect 22244 2496 22250 2508
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 22244 2468 22753 2496
rect 22244 2456 22250 2468
rect 22741 2465 22753 2468
rect 22787 2465 22799 2499
rect 22741 2459 22799 2465
rect 22830 2456 22836 2508
rect 22888 2496 22894 2508
rect 23934 2496 23940 2508
rect 22888 2468 23940 2496
rect 22888 2456 22894 2468
rect 23934 2456 23940 2468
rect 23992 2456 23998 2508
rect 24394 2456 24400 2508
rect 24452 2456 24458 2508
rect 24762 2456 24768 2508
rect 24820 2496 24826 2508
rect 25608 2505 25636 2536
rect 28276 2536 30665 2564
rect 25593 2499 25651 2505
rect 24820 2468 25544 2496
rect 24820 2456 24826 2468
rect 15804 2400 15884 2428
rect 16025 2431 16083 2437
rect 15804 2388 15810 2400
rect 16025 2397 16037 2431
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 17862 2388 17868 2440
rect 17920 2428 17926 2440
rect 18601 2431 18659 2437
rect 18601 2428 18613 2431
rect 17920 2400 18613 2428
rect 17920 2388 17926 2400
rect 18601 2397 18613 2400
rect 18647 2397 18659 2431
rect 18601 2391 18659 2397
rect 20162 2388 20168 2440
rect 20220 2388 20226 2440
rect 20346 2388 20352 2440
rect 20404 2388 20410 2440
rect 20441 2431 20499 2437
rect 20441 2397 20453 2431
rect 20487 2397 20499 2431
rect 20441 2391 20499 2397
rect 16942 2360 16948 2372
rect 14568 2332 16948 2360
rect 13633 2323 13691 2329
rect 16942 2320 16948 2332
rect 17000 2320 17006 2372
rect 17221 2363 17279 2369
rect 17221 2329 17233 2363
rect 17267 2360 17279 2363
rect 20364 2360 20392 2388
rect 17267 2332 20392 2360
rect 20456 2360 20484 2391
rect 21542 2388 21548 2440
rect 21600 2388 21606 2440
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 22373 2431 22431 2437
rect 22373 2428 22385 2431
rect 22336 2400 22385 2428
rect 22336 2388 22342 2400
rect 22373 2397 22385 2400
rect 22419 2397 22431 2431
rect 22373 2391 22431 2397
rect 22554 2388 22560 2440
rect 22612 2388 22618 2440
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2428 23535 2431
rect 23523 2400 24532 2428
rect 23523 2397 23535 2400
rect 23477 2391 23535 2397
rect 23753 2363 23811 2369
rect 23753 2360 23765 2363
rect 20456 2332 23765 2360
rect 17267 2329 17279 2332
rect 17221 2323 17279 2329
rect 23753 2329 23765 2332
rect 23799 2329 23811 2363
rect 24504 2360 24532 2400
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 25314 2388 25320 2440
rect 25372 2388 25378 2440
rect 25516 2428 25544 2468
rect 25593 2465 25605 2499
rect 25639 2465 25651 2499
rect 25593 2459 25651 2465
rect 26234 2456 26240 2508
rect 26292 2456 26298 2508
rect 26418 2456 26424 2508
rect 26476 2496 26482 2508
rect 28276 2505 28304 2536
rect 30653 2533 30665 2536
rect 30699 2564 30711 2567
rect 34146 2564 34152 2576
rect 30699 2536 34152 2564
rect 30699 2533 30711 2536
rect 30653 2527 30711 2533
rect 34146 2524 34152 2536
rect 34204 2524 34210 2576
rect 35802 2524 35808 2576
rect 35860 2524 35866 2576
rect 26789 2499 26847 2505
rect 26789 2496 26801 2499
rect 26476 2468 26801 2496
rect 26476 2456 26482 2468
rect 26789 2465 26801 2468
rect 26835 2465 26847 2499
rect 26789 2459 26847 2465
rect 28261 2499 28319 2505
rect 28261 2465 28273 2499
rect 28307 2465 28319 2499
rect 28261 2459 28319 2465
rect 29825 2499 29883 2505
rect 29825 2465 29837 2499
rect 29871 2496 29883 2499
rect 30282 2496 30288 2508
rect 29871 2468 30288 2496
rect 29871 2465 29883 2468
rect 29825 2459 29883 2465
rect 30282 2456 30288 2468
rect 30340 2456 30346 2508
rect 32214 2456 32220 2508
rect 32272 2456 32278 2508
rect 33413 2499 33471 2505
rect 33413 2465 33425 2499
rect 33459 2496 33471 2499
rect 36464 2496 36492 2604
rect 41598 2592 41604 2604
rect 41656 2592 41662 2644
rect 41693 2635 41751 2641
rect 41693 2601 41705 2635
rect 41739 2632 41751 2635
rect 43530 2632 43536 2644
rect 41739 2604 43536 2632
rect 41739 2601 41751 2604
rect 41693 2595 41751 2601
rect 43530 2592 43536 2604
rect 43588 2592 43594 2644
rect 44726 2592 44732 2644
rect 44784 2632 44790 2644
rect 44821 2635 44879 2641
rect 44821 2632 44833 2635
rect 44784 2604 44833 2632
rect 44784 2592 44790 2604
rect 44821 2601 44833 2604
rect 44867 2601 44879 2635
rect 44821 2595 44879 2601
rect 45830 2592 45836 2644
rect 45888 2632 45894 2644
rect 46842 2632 46848 2644
rect 45888 2604 46848 2632
rect 45888 2592 45894 2604
rect 46842 2592 46848 2604
rect 46900 2592 46906 2644
rect 49970 2592 49976 2644
rect 50028 2592 50034 2644
rect 70857 2635 70915 2641
rect 70857 2601 70869 2635
rect 70903 2632 70915 2635
rect 72234 2632 72240 2644
rect 70903 2604 72240 2632
rect 70903 2601 70915 2604
rect 70857 2595 70915 2601
rect 72234 2592 72240 2604
rect 72292 2592 72298 2644
rect 74077 2635 74135 2641
rect 74077 2601 74089 2635
rect 74123 2632 74135 2635
rect 74626 2632 74632 2644
rect 74123 2604 74632 2632
rect 74123 2601 74135 2604
rect 74077 2595 74135 2601
rect 74626 2592 74632 2604
rect 74684 2592 74690 2644
rect 76650 2592 76656 2644
rect 76708 2632 76714 2644
rect 76837 2635 76895 2641
rect 76837 2632 76849 2635
rect 76708 2604 76849 2632
rect 76708 2592 76714 2604
rect 76837 2601 76849 2604
rect 76883 2601 76895 2635
rect 76837 2595 76895 2601
rect 36541 2567 36599 2573
rect 36541 2533 36553 2567
rect 36587 2564 36599 2567
rect 40957 2567 41015 2573
rect 36587 2536 40172 2564
rect 36587 2533 36599 2536
rect 36541 2527 36599 2533
rect 33459 2468 36492 2496
rect 37553 2499 37611 2505
rect 33459 2465 33471 2468
rect 33413 2459 33471 2465
rect 37553 2465 37565 2499
rect 37599 2496 37611 2499
rect 39850 2496 39856 2508
rect 37599 2468 39856 2496
rect 37599 2465 37611 2468
rect 37553 2459 37611 2465
rect 39850 2456 39856 2468
rect 39908 2456 39914 2508
rect 39945 2499 40003 2505
rect 39945 2465 39957 2499
rect 39991 2496 40003 2499
rect 40034 2496 40040 2508
rect 39991 2468 40040 2496
rect 39991 2465 40003 2468
rect 39945 2459 40003 2465
rect 40034 2456 40040 2468
rect 40092 2456 40098 2508
rect 26329 2431 26387 2437
rect 26329 2428 26341 2431
rect 25516 2400 26341 2428
rect 26329 2397 26341 2400
rect 26375 2397 26387 2431
rect 26329 2391 26387 2397
rect 27890 2388 27896 2440
rect 27948 2388 27954 2440
rect 30098 2428 30104 2440
rect 28000 2400 30104 2428
rect 26970 2360 26976 2372
rect 24504 2332 26976 2360
rect 23753 2323 23811 2329
rect 26970 2320 26976 2332
rect 27028 2320 27034 2372
rect 11848 2264 13124 2292
rect 11848 2252 11854 2264
rect 15194 2252 15200 2304
rect 15252 2252 15258 2304
rect 15562 2252 15568 2304
rect 15620 2252 15626 2304
rect 16390 2252 16396 2304
rect 16448 2292 16454 2304
rect 17957 2295 18015 2301
rect 17957 2292 17969 2295
rect 16448 2264 17969 2292
rect 16448 2252 16454 2264
rect 17957 2261 17969 2264
rect 18003 2261 18015 2295
rect 17957 2255 18015 2261
rect 18046 2252 18052 2304
rect 18104 2252 18110 2304
rect 20346 2252 20352 2304
rect 20404 2252 20410 2304
rect 20622 2252 20628 2304
rect 20680 2252 20686 2304
rect 22094 2252 22100 2304
rect 22152 2252 22158 2304
rect 22189 2295 22247 2301
rect 22189 2261 22201 2295
rect 22235 2292 22247 2295
rect 22830 2292 22836 2304
rect 22235 2264 22836 2292
rect 22235 2261 22247 2264
rect 22189 2255 22247 2261
rect 22830 2252 22836 2264
rect 22888 2252 22894 2304
rect 23385 2295 23443 2301
rect 23385 2261 23397 2295
rect 23431 2292 23443 2295
rect 23842 2292 23848 2304
rect 23431 2264 23848 2292
rect 23431 2261 23443 2264
rect 23385 2255 23443 2261
rect 23842 2252 23848 2264
rect 23900 2252 23906 2304
rect 25133 2295 25191 2301
rect 25133 2261 25145 2295
rect 25179 2292 25191 2295
rect 28000 2292 28028 2400
rect 30098 2388 30104 2400
rect 30156 2388 30162 2440
rect 30193 2431 30251 2437
rect 30193 2397 30205 2431
rect 30239 2428 30251 2431
rect 30374 2428 30380 2440
rect 30239 2400 30380 2428
rect 30239 2397 30251 2400
rect 30193 2391 30251 2397
rect 30374 2388 30380 2400
rect 30432 2388 30438 2440
rect 30837 2431 30895 2437
rect 30837 2397 30849 2431
rect 30883 2428 30895 2431
rect 32766 2428 32772 2440
rect 30883 2400 32772 2428
rect 30883 2397 30895 2400
rect 30837 2391 30895 2397
rect 32766 2388 32772 2400
rect 32824 2388 32830 2440
rect 32861 2431 32919 2437
rect 32861 2397 32873 2431
rect 32907 2428 32919 2431
rect 33318 2428 33324 2440
rect 32907 2400 33324 2428
rect 32907 2397 32919 2400
rect 32861 2391 32919 2397
rect 33318 2388 33324 2400
rect 33376 2388 33382 2440
rect 35250 2388 35256 2440
rect 35308 2388 35314 2440
rect 35618 2388 35624 2440
rect 35676 2388 35682 2440
rect 35986 2388 35992 2440
rect 36044 2388 36050 2440
rect 37921 2431 37979 2437
rect 37921 2397 37933 2431
rect 37967 2397 37979 2431
rect 37921 2391 37979 2397
rect 28810 2320 28816 2372
rect 28868 2320 28874 2372
rect 34146 2320 34152 2372
rect 34204 2360 34210 2372
rect 34241 2363 34299 2369
rect 34241 2360 34253 2363
rect 34204 2332 34253 2360
rect 34204 2320 34210 2332
rect 34241 2329 34253 2332
rect 34287 2329 34299 2363
rect 37936 2360 37964 2391
rect 38010 2388 38016 2440
rect 38068 2428 38074 2440
rect 38289 2431 38347 2437
rect 38289 2428 38301 2431
rect 38068 2400 38301 2428
rect 38068 2388 38074 2400
rect 38289 2397 38301 2400
rect 38335 2397 38347 2431
rect 38289 2391 38347 2397
rect 38838 2388 38844 2440
rect 38896 2388 38902 2440
rect 38930 2388 38936 2440
rect 38988 2388 38994 2440
rect 39669 2431 39727 2437
rect 39669 2397 39681 2431
rect 39715 2397 39727 2431
rect 40144 2428 40172 2536
rect 40957 2533 40969 2567
rect 41003 2564 41015 2567
rect 41966 2564 41972 2576
rect 41003 2536 41972 2564
rect 41003 2533 41015 2536
rect 40957 2527 41015 2533
rect 41966 2524 41972 2536
rect 42024 2524 42030 2576
rect 44634 2524 44640 2576
rect 44692 2564 44698 2576
rect 48133 2567 48191 2573
rect 48133 2564 48145 2567
rect 44692 2536 48145 2564
rect 44692 2524 44698 2536
rect 48133 2533 48145 2536
rect 48179 2533 48191 2567
rect 48133 2527 48191 2533
rect 49602 2524 49608 2576
rect 49660 2564 49666 2576
rect 50709 2567 50767 2573
rect 50709 2564 50721 2567
rect 49660 2536 50721 2564
rect 49660 2524 49666 2536
rect 50709 2533 50721 2536
rect 50755 2533 50767 2567
rect 50709 2527 50767 2533
rect 40589 2499 40647 2505
rect 40589 2465 40601 2499
rect 40635 2496 40647 2499
rect 40635 2468 41000 2496
rect 40635 2465 40647 2468
rect 40589 2459 40647 2465
rect 40773 2431 40831 2437
rect 40773 2428 40785 2431
rect 40144 2400 40785 2428
rect 39669 2391 39727 2397
rect 40773 2397 40785 2400
rect 40819 2397 40831 2431
rect 40972 2428 41000 2468
rect 41138 2456 41144 2508
rect 41196 2456 41202 2508
rect 41386 2468 41828 2496
rect 41386 2428 41414 2468
rect 41800 2437 41828 2468
rect 41874 2456 41880 2508
rect 41932 2496 41938 2508
rect 43809 2499 43867 2505
rect 43809 2496 43821 2499
rect 41932 2468 43821 2496
rect 41932 2456 41938 2468
rect 43809 2465 43821 2468
rect 43855 2465 43867 2499
rect 43809 2459 43867 2465
rect 44266 2456 44272 2508
rect 44324 2496 44330 2508
rect 45373 2499 45431 2505
rect 45373 2496 45385 2499
rect 44324 2468 45385 2496
rect 44324 2456 44330 2468
rect 45373 2465 45385 2468
rect 45419 2465 45431 2499
rect 45373 2459 45431 2465
rect 46385 2499 46443 2505
rect 46385 2465 46397 2499
rect 46431 2465 46443 2499
rect 46385 2459 46443 2465
rect 40972 2400 41414 2428
rect 41785 2431 41843 2437
rect 40773 2391 40831 2397
rect 41785 2397 41797 2431
rect 41831 2397 41843 2431
rect 41785 2391 41843 2397
rect 42981 2431 43039 2437
rect 42981 2397 42993 2431
rect 43027 2428 43039 2431
rect 43349 2431 43407 2437
rect 43349 2428 43361 2431
rect 43027 2400 43361 2428
rect 43027 2397 43039 2400
rect 42981 2391 43039 2397
rect 43349 2397 43361 2400
rect 43395 2397 43407 2431
rect 43349 2391 43407 2397
rect 38746 2360 38752 2372
rect 37936 2332 38752 2360
rect 34241 2323 34299 2329
rect 38746 2320 38752 2332
rect 38804 2320 38810 2372
rect 39684 2360 39712 2391
rect 44818 2388 44824 2440
rect 44876 2428 44882 2440
rect 45189 2431 45247 2437
rect 45189 2428 45201 2431
rect 44876 2400 45201 2428
rect 44876 2388 44882 2400
rect 45189 2397 45201 2400
rect 45235 2397 45247 2431
rect 45189 2391 45247 2397
rect 45281 2431 45339 2437
rect 45281 2397 45293 2431
rect 45327 2428 45339 2431
rect 45830 2428 45836 2440
rect 45327 2400 45836 2428
rect 45327 2397 45339 2400
rect 45281 2391 45339 2397
rect 45830 2388 45836 2400
rect 45888 2388 45894 2440
rect 45922 2388 45928 2440
rect 45980 2388 45986 2440
rect 42702 2360 42708 2372
rect 39684 2332 42708 2360
rect 42702 2320 42708 2332
rect 42760 2320 42766 2372
rect 43806 2320 43812 2372
rect 43864 2360 43870 2372
rect 46400 2360 46428 2459
rect 47026 2456 47032 2508
rect 47084 2496 47090 2508
rect 47949 2499 48007 2505
rect 47949 2496 47961 2499
rect 47084 2468 47961 2496
rect 47084 2456 47090 2468
rect 47949 2465 47961 2468
rect 47995 2465 48007 2499
rect 47949 2459 48007 2465
rect 49421 2499 49479 2505
rect 49421 2465 49433 2499
rect 49467 2496 49479 2499
rect 49786 2496 49792 2508
rect 49467 2468 49792 2496
rect 49467 2465 49479 2468
rect 49421 2459 49479 2465
rect 49786 2456 49792 2468
rect 49844 2456 49850 2508
rect 52086 2456 52092 2508
rect 52144 2456 52150 2508
rect 54018 2456 54024 2508
rect 54076 2456 54082 2508
rect 58161 2499 58219 2505
rect 58161 2465 58173 2499
rect 58207 2496 58219 2499
rect 59265 2499 59323 2505
rect 58207 2468 58848 2496
rect 58207 2465 58219 2468
rect 58161 2459 58219 2465
rect 48314 2388 48320 2440
rect 48372 2388 48378 2440
rect 49878 2388 49884 2440
rect 49936 2388 49942 2440
rect 50522 2388 50528 2440
rect 50580 2388 50586 2440
rect 53006 2388 53012 2440
rect 53064 2388 53070 2440
rect 55033 2431 55091 2437
rect 55033 2397 55045 2431
rect 55079 2428 55091 2431
rect 55306 2428 55312 2440
rect 55079 2400 55312 2428
rect 55079 2397 55091 2400
rect 55033 2391 55091 2397
rect 55306 2388 55312 2400
rect 55364 2388 55370 2440
rect 55398 2388 55404 2440
rect 55456 2428 55462 2440
rect 55493 2431 55551 2437
rect 55493 2428 55505 2431
rect 55456 2400 55505 2428
rect 55456 2388 55462 2400
rect 55493 2397 55505 2400
rect 55539 2397 55551 2431
rect 55493 2391 55551 2397
rect 58618 2388 58624 2440
rect 58676 2388 58682 2440
rect 58820 2437 58848 2468
rect 59265 2465 59277 2499
rect 59311 2465 59323 2499
rect 59265 2459 59323 2465
rect 58805 2431 58863 2437
rect 58805 2397 58817 2431
rect 58851 2397 58863 2431
rect 58805 2391 58863 2397
rect 43864 2332 46428 2360
rect 43864 2320 43870 2332
rect 57330 2320 57336 2372
rect 57388 2360 57394 2372
rect 59280 2360 59308 2459
rect 61746 2456 61752 2508
rect 61804 2456 61810 2508
rect 65518 2456 65524 2508
rect 65576 2456 65582 2508
rect 67634 2456 67640 2508
rect 67692 2456 67698 2508
rect 69474 2456 69480 2508
rect 69532 2456 69538 2508
rect 70302 2456 70308 2508
rect 70360 2496 70366 2508
rect 70360 2468 70716 2496
rect 70360 2456 70366 2468
rect 62758 2388 62764 2440
rect 62816 2388 62822 2440
rect 63126 2388 63132 2440
rect 63184 2428 63190 2440
rect 63221 2431 63279 2437
rect 63221 2428 63233 2431
rect 63184 2400 63233 2428
rect 63184 2388 63190 2400
rect 63221 2397 63233 2400
rect 63267 2397 63279 2431
rect 63221 2391 63279 2397
rect 66254 2388 66260 2440
rect 66312 2388 66318 2440
rect 68278 2388 68284 2440
rect 68336 2388 68342 2440
rect 70486 2388 70492 2440
rect 70544 2388 70550 2440
rect 70688 2437 70716 2468
rect 72602 2456 72608 2508
rect 72660 2456 72666 2508
rect 72786 2456 72792 2508
rect 72844 2496 72850 2508
rect 73157 2499 73215 2505
rect 73157 2496 73169 2499
rect 72844 2468 73169 2496
rect 72844 2456 72850 2468
rect 73157 2465 73169 2468
rect 73203 2465 73215 2499
rect 73157 2459 73215 2465
rect 73525 2499 73583 2505
rect 73525 2465 73537 2499
rect 73571 2496 73583 2499
rect 75454 2496 75460 2508
rect 73571 2468 75460 2496
rect 73571 2465 73583 2468
rect 73525 2459 73583 2465
rect 75454 2456 75460 2468
rect 75512 2456 75518 2508
rect 75733 2499 75791 2505
rect 75733 2465 75745 2499
rect 75779 2496 75791 2499
rect 77389 2499 77447 2505
rect 77389 2496 77401 2499
rect 75779 2468 77401 2496
rect 75779 2465 75791 2468
rect 75733 2459 75791 2465
rect 77389 2465 77401 2468
rect 77435 2465 77447 2499
rect 77389 2459 77447 2465
rect 70673 2431 70731 2437
rect 70673 2397 70685 2431
rect 70719 2397 70731 2431
rect 70673 2391 70731 2397
rect 73062 2388 73068 2440
rect 73120 2388 73126 2440
rect 76190 2388 76196 2440
rect 76248 2388 76254 2440
rect 57388 2332 59308 2360
rect 57388 2320 57394 2332
rect 25179 2264 28028 2292
rect 25179 2261 25191 2264
rect 25133 2255 25191 2261
rect 28074 2252 28080 2304
rect 28132 2252 28138 2304
rect 31386 2252 31392 2304
rect 31444 2252 31450 2304
rect 34974 2252 34980 2304
rect 35032 2292 35038 2304
rect 38289 2295 38347 2301
rect 38289 2292 38301 2295
rect 35032 2264 38301 2292
rect 35032 2252 35038 2264
rect 38289 2261 38301 2264
rect 38335 2261 38347 2295
rect 38289 2255 38347 2261
rect 47394 2252 47400 2304
rect 47452 2252 47458 2304
rect 2024 2202 77924 2224
rect 2024 2150 5794 2202
rect 5846 2150 5858 2202
rect 5910 2150 5922 2202
rect 5974 2150 5986 2202
rect 6038 2150 6050 2202
rect 6102 2150 36514 2202
rect 36566 2150 36578 2202
rect 36630 2150 36642 2202
rect 36694 2150 36706 2202
rect 36758 2150 36770 2202
rect 36822 2150 67234 2202
rect 67286 2150 67298 2202
rect 67350 2150 67362 2202
rect 67414 2150 67426 2202
rect 67478 2150 67490 2202
rect 67542 2150 77924 2202
rect 2024 2128 77924 2150
rect 6270 2048 6276 2100
rect 6328 2088 6334 2100
rect 11606 2088 11612 2100
rect 6328 2060 11612 2088
rect 6328 2048 6334 2060
rect 11606 2048 11612 2060
rect 11664 2048 11670 2100
rect 12986 2048 12992 2100
rect 13044 2088 13050 2100
rect 13044 2060 16620 2088
rect 13044 2048 13050 2060
rect 9122 1980 9128 2032
rect 9180 2020 9186 2032
rect 16390 2020 16396 2032
rect 9180 1992 16396 2020
rect 9180 1980 9186 1992
rect 16390 1980 16396 1992
rect 16448 1980 16454 2032
rect 10594 1912 10600 1964
rect 10652 1952 10658 1964
rect 13354 1952 13360 1964
rect 10652 1924 13360 1952
rect 10652 1912 10658 1924
rect 13354 1912 13360 1924
rect 13412 1912 13418 1964
rect 16592 1952 16620 2060
rect 20622 2048 20628 2100
rect 20680 2088 20686 2100
rect 27522 2088 27528 2100
rect 20680 2060 27528 2088
rect 20680 2048 20686 2060
rect 27522 2048 27528 2060
rect 27580 2048 27586 2100
rect 35986 2048 35992 2100
rect 36044 2088 36050 2100
rect 47394 2088 47400 2100
rect 36044 2060 47400 2088
rect 36044 2048 36050 2060
rect 47394 2048 47400 2060
rect 47452 2048 47458 2100
rect 22094 1980 22100 2032
rect 22152 2020 22158 2032
rect 22152 1992 30604 2020
rect 22152 1980 22158 1992
rect 23566 1952 23572 1964
rect 16592 1924 23572 1952
rect 23566 1912 23572 1924
rect 23624 1912 23630 1964
rect 23842 1912 23848 1964
rect 23900 1952 23906 1964
rect 30466 1952 30472 1964
rect 23900 1924 30472 1952
rect 23900 1912 23906 1924
rect 30466 1912 30472 1924
rect 30524 1912 30530 1964
rect 5718 1844 5724 1896
rect 5776 1884 5782 1896
rect 11698 1884 11704 1896
rect 5776 1856 11704 1884
rect 5776 1844 5782 1856
rect 11698 1844 11704 1856
rect 11756 1844 11762 1896
rect 16298 1844 16304 1896
rect 16356 1884 16362 1896
rect 16356 1856 26924 1884
rect 16356 1844 16362 1856
rect 8294 1776 8300 1828
rect 8352 1816 8358 1828
rect 18046 1816 18052 1828
rect 8352 1788 18052 1816
rect 8352 1776 8358 1788
rect 18046 1776 18052 1788
rect 18104 1776 18110 1828
rect 20162 1776 20168 1828
rect 20220 1816 20226 1828
rect 26326 1816 26332 1828
rect 20220 1788 26332 1816
rect 20220 1776 20226 1788
rect 26326 1776 26332 1788
rect 26384 1776 26390 1828
rect 8938 1708 8944 1760
rect 8996 1748 9002 1760
rect 18138 1748 18144 1760
rect 8996 1720 18144 1748
rect 8996 1708 9002 1720
rect 18138 1708 18144 1720
rect 18196 1708 18202 1760
rect 8570 1640 8576 1692
rect 8628 1680 8634 1692
rect 8628 1652 12434 1680
rect 8628 1640 8634 1652
rect 12406 1612 12434 1652
rect 13354 1640 13360 1692
rect 13412 1680 13418 1692
rect 25682 1680 25688 1692
rect 13412 1652 25688 1680
rect 13412 1640 13418 1652
rect 25682 1640 25688 1652
rect 25740 1640 25746 1692
rect 15194 1612 15200 1624
rect 12406 1584 15200 1612
rect 15194 1572 15200 1584
rect 15252 1572 15258 1624
rect 20346 1572 20352 1624
rect 20404 1612 20410 1624
rect 25774 1612 25780 1624
rect 20404 1584 25780 1612
rect 20404 1572 20410 1584
rect 25774 1572 25780 1584
rect 25832 1572 25838 1624
rect 26896 1612 26924 1856
rect 30576 1680 30604 1992
rect 31570 1980 31576 2032
rect 31628 2020 31634 2032
rect 38930 2020 38936 2032
rect 31628 1992 38936 2020
rect 31628 1980 31634 1992
rect 38930 1980 38936 1992
rect 38988 1980 38994 2032
rect 44450 1980 44456 2032
rect 44508 2020 44514 2032
rect 50522 2020 50528 2032
rect 44508 1992 50528 2020
rect 44508 1980 44514 1992
rect 50522 1980 50528 1992
rect 50580 1980 50586 2032
rect 35618 1912 35624 1964
rect 35676 1952 35682 1964
rect 40678 1952 40684 1964
rect 35676 1924 40684 1952
rect 35676 1912 35682 1924
rect 40678 1912 40684 1924
rect 40736 1912 40742 1964
rect 35802 1844 35808 1896
rect 35860 1884 35866 1896
rect 40494 1884 40500 1896
rect 35860 1856 40500 1884
rect 35860 1844 35866 1856
rect 40494 1844 40500 1856
rect 40552 1844 40558 1896
rect 32766 1776 32772 1828
rect 32824 1816 32830 1828
rect 39206 1816 39212 1828
rect 32824 1788 39212 1816
rect 32824 1776 32830 1788
rect 39206 1776 39212 1788
rect 39264 1776 39270 1828
rect 31386 1708 31392 1760
rect 31444 1748 31450 1760
rect 41230 1748 41236 1760
rect 31444 1720 41236 1748
rect 31444 1708 31450 1720
rect 41230 1708 41236 1720
rect 41288 1708 41294 1760
rect 36906 1680 36912 1692
rect 30576 1652 36912 1680
rect 36906 1640 36912 1652
rect 36964 1640 36970 1692
rect 35710 1612 35716 1624
rect 26896 1584 35716 1612
rect 35710 1572 35716 1584
rect 35768 1572 35774 1624
rect 14918 1300 14924 1352
rect 14976 1340 14982 1352
rect 16114 1340 16120 1352
rect 14976 1312 16120 1340
rect 14976 1300 14982 1312
rect 16114 1300 16120 1312
rect 16172 1300 16178 1352
rect 42518 1300 42524 1352
rect 42576 1340 42582 1352
rect 47118 1340 47124 1352
rect 42576 1312 47124 1340
rect 42576 1300 42582 1312
rect 47118 1300 47124 1312
rect 47176 1300 47182 1352
rect 40586 1096 40592 1148
rect 40644 1136 40650 1148
rect 45186 1136 45192 1148
rect 40644 1108 45192 1136
rect 40644 1096 40650 1108
rect 45186 1096 45192 1108
rect 45244 1096 45250 1148
rect 7650 280 7656 332
rect 7708 320 7714 332
rect 18598 320 18604 332
rect 7708 292 18604 320
rect 7708 280 7714 292
rect 18598 280 18604 292
rect 18656 280 18662 332
rect 21726 280 21732 332
rect 21784 320 21790 332
rect 31478 320 31484 332
rect 21784 292 31484 320
rect 21784 280 21790 292
rect 31478 280 31484 292
rect 31536 280 31542 332
rect 10134 212 10140 264
rect 10192 252 10198 264
rect 21174 252 21180 264
rect 10192 224 21180 252
rect 10192 212 10198 224
rect 21174 212 21180 224
rect 21232 212 21238 264
rect 21634 212 21640 264
rect 21692 252 21698 264
rect 32766 252 32772 264
rect 21692 224 32772 252
rect 21692 212 21698 224
rect 32766 212 32772 224
rect 32824 212 32830 264
rect 8386 144 8392 196
rect 8444 184 8450 196
rect 23106 184 23112 196
rect 8444 156 23112 184
rect 8444 144 8450 156
rect 23106 144 23112 156
rect 23164 144 23170 196
rect 9122 76 9128 128
rect 9180 116 9186 128
rect 23474 116 23480 128
rect 9180 88 23480 116
rect 9180 76 9186 88
rect 23474 76 23480 88
rect 23532 76 23538 128
<< via1 >>
rect 5134 37510 5186 37562
rect 5198 37510 5250 37562
rect 5262 37510 5314 37562
rect 5326 37510 5378 37562
rect 5390 37510 5442 37562
rect 35854 37510 35906 37562
rect 35918 37510 35970 37562
rect 35982 37510 36034 37562
rect 36046 37510 36098 37562
rect 36110 37510 36162 37562
rect 66574 37510 66626 37562
rect 66638 37510 66690 37562
rect 66702 37510 66754 37562
rect 66766 37510 66818 37562
rect 66830 37510 66882 37562
rect 2228 37272 2280 37324
rect 13268 37272 13320 37324
rect 33508 37272 33560 37324
rect 39028 37272 39080 37324
rect 3516 37247 3568 37256
rect 3516 37213 3525 37247
rect 3525 37213 3559 37247
rect 3559 37213 3568 37247
rect 3516 37204 3568 37213
rect 5908 37247 5960 37256
rect 5908 37213 5917 37247
rect 5917 37213 5951 37247
rect 5951 37213 5960 37247
rect 5908 37204 5960 37213
rect 7012 37247 7064 37256
rect 7012 37213 7021 37247
rect 7021 37213 7055 37247
rect 7055 37213 7064 37247
rect 7012 37204 7064 37213
rect 7748 37204 7800 37256
rect 7932 37204 7984 37256
rect 11428 37204 11480 37256
rect 11888 37204 11940 37256
rect 14556 37247 14608 37256
rect 14556 37213 14565 37247
rect 14565 37213 14599 37247
rect 14599 37213 14608 37247
rect 14556 37204 14608 37213
rect 15108 37204 15160 37256
rect 18696 37247 18748 37256
rect 18696 37213 18705 37247
rect 18705 37213 18739 37247
rect 18739 37213 18748 37247
rect 18696 37204 18748 37213
rect 18788 37204 18840 37256
rect 20628 37204 20680 37256
rect 21916 37247 21968 37256
rect 21916 37213 21925 37247
rect 21925 37213 21959 37247
rect 21959 37213 21968 37247
rect 21916 37204 21968 37213
rect 22468 37204 22520 37256
rect 26056 37204 26108 37256
rect 27988 37204 28040 37256
rect 29276 37247 29328 37256
rect 29276 37213 29285 37247
rect 29285 37213 29319 37247
rect 29319 37213 29328 37247
rect 29276 37204 29328 37213
rect 31668 37204 31720 37256
rect 32772 37247 32824 37256
rect 32772 37213 32781 37247
rect 32781 37213 32815 37247
rect 32815 37213 32824 37247
rect 32772 37204 32824 37213
rect 33784 37247 33836 37256
rect 33784 37213 33793 37247
rect 33793 37213 33827 37247
rect 33827 37213 33836 37247
rect 33784 37204 33836 37213
rect 37004 37204 37056 37256
rect 37188 37204 37240 37256
rect 39120 37247 39172 37256
rect 39120 37213 39129 37247
rect 39129 37213 39163 37247
rect 39163 37213 39172 37247
rect 39120 37204 39172 37213
rect 40868 37204 40920 37256
rect 41052 37204 41104 37256
rect 43352 37247 43404 37256
rect 43352 37213 43361 37247
rect 43361 37213 43395 37247
rect 43395 37213 43404 37247
rect 43352 37204 43404 37213
rect 46480 37247 46532 37256
rect 46480 37213 46489 37247
rect 46489 37213 46523 37247
rect 46523 37213 46532 37247
rect 46480 37204 46532 37213
rect 48228 37204 48280 37256
rect 51908 37204 51960 37256
rect 52092 37204 52144 37256
rect 53840 37247 53892 37256
rect 53840 37213 53849 37247
rect 53849 37213 53883 37247
rect 53883 37213 53892 37247
rect 53840 37204 53892 37213
rect 55588 37204 55640 37256
rect 58808 37247 58860 37256
rect 58808 37213 58817 37247
rect 58817 37213 58851 37247
rect 58851 37213 58860 37247
rect 58808 37204 58860 37213
rect 15016 37136 15068 37188
rect 22560 37136 22612 37188
rect 26148 37136 26200 37188
rect 42708 37136 42760 37188
rect 46388 37136 46440 37188
rect 48136 37136 48188 37188
rect 53748 37136 53800 37188
rect 55680 37136 55732 37188
rect 57428 37136 57480 37188
rect 5794 36966 5846 37018
rect 5858 36966 5910 37018
rect 5922 36966 5974 37018
rect 5986 36966 6038 37018
rect 6050 36966 6102 37018
rect 36514 36966 36566 37018
rect 36578 36966 36630 37018
rect 36642 36966 36694 37018
rect 36706 36966 36758 37018
rect 36770 36966 36822 37018
rect 67234 36966 67286 37018
rect 67298 36966 67350 37018
rect 67362 36966 67414 37018
rect 67426 36966 67478 37018
rect 67490 36966 67542 37018
rect 7748 36907 7800 36916
rect 7748 36873 7757 36907
rect 7757 36873 7791 36907
rect 7791 36873 7800 36907
rect 7748 36864 7800 36873
rect 11888 36907 11940 36916
rect 11888 36873 11897 36907
rect 11897 36873 11931 36907
rect 11931 36873 11940 36907
rect 11888 36864 11940 36873
rect 15108 36907 15160 36916
rect 15108 36873 15117 36907
rect 15117 36873 15151 36907
rect 15151 36873 15160 36907
rect 15108 36864 15160 36873
rect 18696 36864 18748 36916
rect 22468 36907 22520 36916
rect 22468 36873 22477 36907
rect 22477 36873 22511 36907
rect 22511 36873 22520 36907
rect 22468 36864 22520 36873
rect 26056 36864 26108 36916
rect 4068 36796 4120 36848
rect 9588 36796 9640 36848
rect 16948 36796 17000 36848
rect 24308 36796 24360 36848
rect 10876 36771 10928 36780
rect 10876 36737 10885 36771
rect 10885 36737 10919 36771
rect 10919 36737 10928 36771
rect 10876 36728 10928 36737
rect 11796 36771 11848 36780
rect 11796 36737 11805 36771
rect 11805 36737 11839 36771
rect 11839 36737 11848 36771
rect 11796 36728 11848 36737
rect 18972 36771 19024 36780
rect 18972 36737 18981 36771
rect 18981 36737 19015 36771
rect 19015 36737 19024 36771
rect 18972 36728 19024 36737
rect 25780 36771 25832 36780
rect 25780 36737 25789 36771
rect 25789 36737 25823 36771
rect 25823 36737 25832 36771
rect 25780 36728 25832 36737
rect 29828 36796 29880 36848
rect 33784 36907 33836 36916
rect 33784 36873 33793 36907
rect 33793 36873 33827 36907
rect 33827 36873 33836 36907
rect 33784 36864 33836 36873
rect 37004 36907 37056 36916
rect 37004 36873 37013 36907
rect 37013 36873 37047 36907
rect 37047 36873 37056 36907
rect 37004 36864 37056 36873
rect 40868 36907 40920 36916
rect 40868 36873 40877 36907
rect 40877 36873 40911 36907
rect 40911 36873 40920 36907
rect 40868 36864 40920 36873
rect 48228 36907 48280 36916
rect 48228 36873 48237 36907
rect 48237 36873 48271 36907
rect 48271 36873 48280 36907
rect 48228 36864 48280 36873
rect 51908 36907 51960 36916
rect 51908 36873 51917 36907
rect 51917 36873 51951 36907
rect 51951 36873 51960 36907
rect 51908 36864 51960 36873
rect 55588 36907 55640 36916
rect 55588 36873 55597 36907
rect 55597 36873 55631 36907
rect 55631 36873 55640 36907
rect 55588 36864 55640 36873
rect 11796 36592 11848 36644
rect 35440 36771 35492 36780
rect 35440 36737 35449 36771
rect 35449 36737 35483 36771
rect 35483 36737 35492 36771
rect 35440 36728 35492 36737
rect 35348 36660 35400 36712
rect 44732 36660 44784 36712
rect 50160 36771 50212 36780
rect 50160 36737 50169 36771
rect 50169 36737 50203 36771
rect 50203 36737 50212 36771
rect 50160 36728 50212 36737
rect 59268 36796 59320 36848
rect 50068 36660 50120 36712
rect 5134 36422 5186 36474
rect 5198 36422 5250 36474
rect 5262 36422 5314 36474
rect 5326 36422 5378 36474
rect 5390 36422 5442 36474
rect 35854 36422 35906 36474
rect 35918 36422 35970 36474
rect 35982 36422 36034 36474
rect 36046 36422 36098 36474
rect 36110 36422 36162 36474
rect 66574 36422 66626 36474
rect 66638 36422 66690 36474
rect 66702 36422 66754 36474
rect 66766 36422 66818 36474
rect 66830 36422 66882 36474
rect 5794 35878 5846 35930
rect 5858 35878 5910 35930
rect 5922 35878 5974 35930
rect 5986 35878 6038 35930
rect 6050 35878 6102 35930
rect 36514 35878 36566 35930
rect 36578 35878 36630 35930
rect 36642 35878 36694 35930
rect 36706 35878 36758 35930
rect 36770 35878 36822 35930
rect 67234 35878 67286 35930
rect 67298 35878 67350 35930
rect 67362 35878 67414 35930
rect 67426 35878 67478 35930
rect 67490 35878 67542 35930
rect 5134 35334 5186 35386
rect 5198 35334 5250 35386
rect 5262 35334 5314 35386
rect 5326 35334 5378 35386
rect 5390 35334 5442 35386
rect 35854 35334 35906 35386
rect 35918 35334 35970 35386
rect 35982 35334 36034 35386
rect 36046 35334 36098 35386
rect 36110 35334 36162 35386
rect 66574 35334 66626 35386
rect 66638 35334 66690 35386
rect 66702 35334 66754 35386
rect 66766 35334 66818 35386
rect 66830 35334 66882 35386
rect 5794 34790 5846 34842
rect 5858 34790 5910 34842
rect 5922 34790 5974 34842
rect 5986 34790 6038 34842
rect 6050 34790 6102 34842
rect 36514 34790 36566 34842
rect 36578 34790 36630 34842
rect 36642 34790 36694 34842
rect 36706 34790 36758 34842
rect 36770 34790 36822 34842
rect 67234 34790 67286 34842
rect 67298 34790 67350 34842
rect 67362 34790 67414 34842
rect 67426 34790 67478 34842
rect 67490 34790 67542 34842
rect 5134 34246 5186 34298
rect 5198 34246 5250 34298
rect 5262 34246 5314 34298
rect 5326 34246 5378 34298
rect 5390 34246 5442 34298
rect 35854 34246 35906 34298
rect 35918 34246 35970 34298
rect 35982 34246 36034 34298
rect 36046 34246 36098 34298
rect 36110 34246 36162 34298
rect 66574 34246 66626 34298
rect 66638 34246 66690 34298
rect 66702 34246 66754 34298
rect 66766 34246 66818 34298
rect 66830 34246 66882 34298
rect 5794 33702 5846 33754
rect 5858 33702 5910 33754
rect 5922 33702 5974 33754
rect 5986 33702 6038 33754
rect 6050 33702 6102 33754
rect 36514 33702 36566 33754
rect 36578 33702 36630 33754
rect 36642 33702 36694 33754
rect 36706 33702 36758 33754
rect 36770 33702 36822 33754
rect 67234 33702 67286 33754
rect 67298 33702 67350 33754
rect 67362 33702 67414 33754
rect 67426 33702 67478 33754
rect 67490 33702 67542 33754
rect 5134 33158 5186 33210
rect 5198 33158 5250 33210
rect 5262 33158 5314 33210
rect 5326 33158 5378 33210
rect 5390 33158 5442 33210
rect 35854 33158 35906 33210
rect 35918 33158 35970 33210
rect 35982 33158 36034 33210
rect 36046 33158 36098 33210
rect 36110 33158 36162 33210
rect 66574 33158 66626 33210
rect 66638 33158 66690 33210
rect 66702 33158 66754 33210
rect 66766 33158 66818 33210
rect 66830 33158 66882 33210
rect 25780 33056 25832 33108
rect 27344 33056 27396 33108
rect 5794 32614 5846 32666
rect 5858 32614 5910 32666
rect 5922 32614 5974 32666
rect 5986 32614 6038 32666
rect 6050 32614 6102 32666
rect 36514 32614 36566 32666
rect 36578 32614 36630 32666
rect 36642 32614 36694 32666
rect 36706 32614 36758 32666
rect 36770 32614 36822 32666
rect 67234 32614 67286 32666
rect 67298 32614 67350 32666
rect 67362 32614 67414 32666
rect 67426 32614 67478 32666
rect 67490 32614 67542 32666
rect 26332 32376 26384 32428
rect 43352 32376 43404 32428
rect 5134 32070 5186 32122
rect 5198 32070 5250 32122
rect 5262 32070 5314 32122
rect 5326 32070 5378 32122
rect 5390 32070 5442 32122
rect 35854 32070 35906 32122
rect 35918 32070 35970 32122
rect 35982 32070 36034 32122
rect 36046 32070 36098 32122
rect 36110 32070 36162 32122
rect 66574 32070 66626 32122
rect 66638 32070 66690 32122
rect 66702 32070 66754 32122
rect 66766 32070 66818 32122
rect 66830 32070 66882 32122
rect 5794 31526 5846 31578
rect 5858 31526 5910 31578
rect 5922 31526 5974 31578
rect 5986 31526 6038 31578
rect 6050 31526 6102 31578
rect 36514 31526 36566 31578
rect 36578 31526 36630 31578
rect 36642 31526 36694 31578
rect 36706 31526 36758 31578
rect 36770 31526 36822 31578
rect 67234 31526 67286 31578
rect 67298 31526 67350 31578
rect 67362 31526 67414 31578
rect 67426 31526 67478 31578
rect 67490 31526 67542 31578
rect 5134 30982 5186 31034
rect 5198 30982 5250 31034
rect 5262 30982 5314 31034
rect 5326 30982 5378 31034
rect 5390 30982 5442 31034
rect 35854 30982 35906 31034
rect 35918 30982 35970 31034
rect 35982 30982 36034 31034
rect 36046 30982 36098 31034
rect 36110 30982 36162 31034
rect 66574 30982 66626 31034
rect 66638 30982 66690 31034
rect 66702 30982 66754 31034
rect 66766 30982 66818 31034
rect 66830 30982 66882 31034
rect 5794 30438 5846 30490
rect 5858 30438 5910 30490
rect 5922 30438 5974 30490
rect 5986 30438 6038 30490
rect 6050 30438 6102 30490
rect 36514 30438 36566 30490
rect 36578 30438 36630 30490
rect 36642 30438 36694 30490
rect 36706 30438 36758 30490
rect 36770 30438 36822 30490
rect 67234 30438 67286 30490
rect 67298 30438 67350 30490
rect 67362 30438 67414 30490
rect 67426 30438 67478 30490
rect 67490 30438 67542 30490
rect 5134 29894 5186 29946
rect 5198 29894 5250 29946
rect 5262 29894 5314 29946
rect 5326 29894 5378 29946
rect 5390 29894 5442 29946
rect 35854 29894 35906 29946
rect 35918 29894 35970 29946
rect 35982 29894 36034 29946
rect 36046 29894 36098 29946
rect 36110 29894 36162 29946
rect 66574 29894 66626 29946
rect 66638 29894 66690 29946
rect 66702 29894 66754 29946
rect 66766 29894 66818 29946
rect 66830 29894 66882 29946
rect 26056 29588 26108 29640
rect 50160 29588 50212 29640
rect 5794 29350 5846 29402
rect 5858 29350 5910 29402
rect 5922 29350 5974 29402
rect 5986 29350 6038 29402
rect 6050 29350 6102 29402
rect 36514 29350 36566 29402
rect 36578 29350 36630 29402
rect 36642 29350 36694 29402
rect 36706 29350 36758 29402
rect 36770 29350 36822 29402
rect 67234 29350 67286 29402
rect 67298 29350 67350 29402
rect 67362 29350 67414 29402
rect 67426 29350 67478 29402
rect 67490 29350 67542 29402
rect 5134 28806 5186 28858
rect 5198 28806 5250 28858
rect 5262 28806 5314 28858
rect 5326 28806 5378 28858
rect 5390 28806 5442 28858
rect 35854 28806 35906 28858
rect 35918 28806 35970 28858
rect 35982 28806 36034 28858
rect 36046 28806 36098 28858
rect 36110 28806 36162 28858
rect 66574 28806 66626 28858
rect 66638 28806 66690 28858
rect 66702 28806 66754 28858
rect 66766 28806 66818 28858
rect 66830 28806 66882 28858
rect 5794 28262 5846 28314
rect 5858 28262 5910 28314
rect 5922 28262 5974 28314
rect 5986 28262 6038 28314
rect 6050 28262 6102 28314
rect 36514 28262 36566 28314
rect 36578 28262 36630 28314
rect 36642 28262 36694 28314
rect 36706 28262 36758 28314
rect 36770 28262 36822 28314
rect 67234 28262 67286 28314
rect 67298 28262 67350 28314
rect 67362 28262 67414 28314
rect 67426 28262 67478 28314
rect 67490 28262 67542 28314
rect 5134 27718 5186 27770
rect 5198 27718 5250 27770
rect 5262 27718 5314 27770
rect 5326 27718 5378 27770
rect 5390 27718 5442 27770
rect 35854 27718 35906 27770
rect 35918 27718 35970 27770
rect 35982 27718 36034 27770
rect 36046 27718 36098 27770
rect 36110 27718 36162 27770
rect 66574 27718 66626 27770
rect 66638 27718 66690 27770
rect 66702 27718 66754 27770
rect 66766 27718 66818 27770
rect 66830 27718 66882 27770
rect 5794 27174 5846 27226
rect 5858 27174 5910 27226
rect 5922 27174 5974 27226
rect 5986 27174 6038 27226
rect 6050 27174 6102 27226
rect 36514 27174 36566 27226
rect 36578 27174 36630 27226
rect 36642 27174 36694 27226
rect 36706 27174 36758 27226
rect 36770 27174 36822 27226
rect 67234 27174 67286 27226
rect 67298 27174 67350 27226
rect 67362 27174 67414 27226
rect 67426 27174 67478 27226
rect 67490 27174 67542 27226
rect 25688 26868 25740 26920
rect 53840 26868 53892 26920
rect 5134 26630 5186 26682
rect 5198 26630 5250 26682
rect 5262 26630 5314 26682
rect 5326 26630 5378 26682
rect 5390 26630 5442 26682
rect 35854 26630 35906 26682
rect 35918 26630 35970 26682
rect 35982 26630 36034 26682
rect 36046 26630 36098 26682
rect 36110 26630 36162 26682
rect 66574 26630 66626 26682
rect 66638 26630 66690 26682
rect 66702 26630 66754 26682
rect 66766 26630 66818 26682
rect 66830 26630 66882 26682
rect 5794 26086 5846 26138
rect 5858 26086 5910 26138
rect 5922 26086 5974 26138
rect 5986 26086 6038 26138
rect 6050 26086 6102 26138
rect 36514 26086 36566 26138
rect 36578 26086 36630 26138
rect 36642 26086 36694 26138
rect 36706 26086 36758 26138
rect 36770 26086 36822 26138
rect 67234 26086 67286 26138
rect 67298 26086 67350 26138
rect 67362 26086 67414 26138
rect 67426 26086 67478 26138
rect 67490 26086 67542 26138
rect 5134 25542 5186 25594
rect 5198 25542 5250 25594
rect 5262 25542 5314 25594
rect 5326 25542 5378 25594
rect 5390 25542 5442 25594
rect 35854 25542 35906 25594
rect 35918 25542 35970 25594
rect 35982 25542 36034 25594
rect 36046 25542 36098 25594
rect 36110 25542 36162 25594
rect 66574 25542 66626 25594
rect 66638 25542 66690 25594
rect 66702 25542 66754 25594
rect 66766 25542 66818 25594
rect 66830 25542 66882 25594
rect 5794 24998 5846 25050
rect 5858 24998 5910 25050
rect 5922 24998 5974 25050
rect 5986 24998 6038 25050
rect 6050 24998 6102 25050
rect 36514 24998 36566 25050
rect 36578 24998 36630 25050
rect 36642 24998 36694 25050
rect 36706 24998 36758 25050
rect 36770 24998 36822 25050
rect 67234 24998 67286 25050
rect 67298 24998 67350 25050
rect 67362 24998 67414 25050
rect 67426 24998 67478 25050
rect 67490 24998 67542 25050
rect 5134 24454 5186 24506
rect 5198 24454 5250 24506
rect 5262 24454 5314 24506
rect 5326 24454 5378 24506
rect 5390 24454 5442 24506
rect 35854 24454 35906 24506
rect 35918 24454 35970 24506
rect 35982 24454 36034 24506
rect 36046 24454 36098 24506
rect 36110 24454 36162 24506
rect 66574 24454 66626 24506
rect 66638 24454 66690 24506
rect 66702 24454 66754 24506
rect 66766 24454 66818 24506
rect 66830 24454 66882 24506
rect 25504 24080 25556 24132
rect 46480 24080 46532 24132
rect 5794 23910 5846 23962
rect 5858 23910 5910 23962
rect 5922 23910 5974 23962
rect 5986 23910 6038 23962
rect 6050 23910 6102 23962
rect 36514 23910 36566 23962
rect 36578 23910 36630 23962
rect 36642 23910 36694 23962
rect 36706 23910 36758 23962
rect 36770 23910 36822 23962
rect 67234 23910 67286 23962
rect 67298 23910 67350 23962
rect 67362 23910 67414 23962
rect 67426 23910 67478 23962
rect 67490 23910 67542 23962
rect 5134 23366 5186 23418
rect 5198 23366 5250 23418
rect 5262 23366 5314 23418
rect 5326 23366 5378 23418
rect 5390 23366 5442 23418
rect 35854 23366 35906 23418
rect 35918 23366 35970 23418
rect 35982 23366 36034 23418
rect 36046 23366 36098 23418
rect 36110 23366 36162 23418
rect 66574 23366 66626 23418
rect 66638 23366 66690 23418
rect 66702 23366 66754 23418
rect 66766 23366 66818 23418
rect 66830 23366 66882 23418
rect 5794 22822 5846 22874
rect 5858 22822 5910 22874
rect 5922 22822 5974 22874
rect 5986 22822 6038 22874
rect 6050 22822 6102 22874
rect 36514 22822 36566 22874
rect 36578 22822 36630 22874
rect 36642 22822 36694 22874
rect 36706 22822 36758 22874
rect 36770 22822 36822 22874
rect 67234 22822 67286 22874
rect 67298 22822 67350 22874
rect 67362 22822 67414 22874
rect 67426 22822 67478 22874
rect 67490 22822 67542 22874
rect 5134 22278 5186 22330
rect 5198 22278 5250 22330
rect 5262 22278 5314 22330
rect 5326 22278 5378 22330
rect 5390 22278 5442 22330
rect 35854 22278 35906 22330
rect 35918 22278 35970 22330
rect 35982 22278 36034 22330
rect 36046 22278 36098 22330
rect 36110 22278 36162 22330
rect 66574 22278 66626 22330
rect 66638 22278 66690 22330
rect 66702 22278 66754 22330
rect 66766 22278 66818 22330
rect 66830 22278 66882 22330
rect 5794 21734 5846 21786
rect 5858 21734 5910 21786
rect 5922 21734 5974 21786
rect 5986 21734 6038 21786
rect 6050 21734 6102 21786
rect 36514 21734 36566 21786
rect 36578 21734 36630 21786
rect 36642 21734 36694 21786
rect 36706 21734 36758 21786
rect 36770 21734 36822 21786
rect 67234 21734 67286 21786
rect 67298 21734 67350 21786
rect 67362 21734 67414 21786
rect 67426 21734 67478 21786
rect 67490 21734 67542 21786
rect 5134 21190 5186 21242
rect 5198 21190 5250 21242
rect 5262 21190 5314 21242
rect 5326 21190 5378 21242
rect 5390 21190 5442 21242
rect 35854 21190 35906 21242
rect 35918 21190 35970 21242
rect 35982 21190 36034 21242
rect 36046 21190 36098 21242
rect 36110 21190 36162 21242
rect 66574 21190 66626 21242
rect 66638 21190 66690 21242
rect 66702 21190 66754 21242
rect 66766 21190 66818 21242
rect 66830 21190 66882 21242
rect 5794 20646 5846 20698
rect 5858 20646 5910 20698
rect 5922 20646 5974 20698
rect 5986 20646 6038 20698
rect 6050 20646 6102 20698
rect 36514 20646 36566 20698
rect 36578 20646 36630 20698
rect 36642 20646 36694 20698
rect 36706 20646 36758 20698
rect 36770 20646 36822 20698
rect 67234 20646 67286 20698
rect 67298 20646 67350 20698
rect 67362 20646 67414 20698
rect 67426 20646 67478 20698
rect 67490 20646 67542 20698
rect 5134 20102 5186 20154
rect 5198 20102 5250 20154
rect 5262 20102 5314 20154
rect 5326 20102 5378 20154
rect 5390 20102 5442 20154
rect 35854 20102 35906 20154
rect 35918 20102 35970 20154
rect 35982 20102 36034 20154
rect 36046 20102 36098 20154
rect 36110 20102 36162 20154
rect 66574 20102 66626 20154
rect 66638 20102 66690 20154
rect 66702 20102 66754 20154
rect 66766 20102 66818 20154
rect 66830 20102 66882 20154
rect 5794 19558 5846 19610
rect 5858 19558 5910 19610
rect 5922 19558 5974 19610
rect 5986 19558 6038 19610
rect 6050 19558 6102 19610
rect 36514 19558 36566 19610
rect 36578 19558 36630 19610
rect 36642 19558 36694 19610
rect 36706 19558 36758 19610
rect 36770 19558 36822 19610
rect 67234 19558 67286 19610
rect 67298 19558 67350 19610
rect 67362 19558 67414 19610
rect 67426 19558 67478 19610
rect 67490 19558 67542 19610
rect 5134 19014 5186 19066
rect 5198 19014 5250 19066
rect 5262 19014 5314 19066
rect 5326 19014 5378 19066
rect 5390 19014 5442 19066
rect 35854 19014 35906 19066
rect 35918 19014 35970 19066
rect 35982 19014 36034 19066
rect 36046 19014 36098 19066
rect 36110 19014 36162 19066
rect 66574 19014 66626 19066
rect 66638 19014 66690 19066
rect 66702 19014 66754 19066
rect 66766 19014 66818 19066
rect 66830 19014 66882 19066
rect 5794 18470 5846 18522
rect 5858 18470 5910 18522
rect 5922 18470 5974 18522
rect 5986 18470 6038 18522
rect 6050 18470 6102 18522
rect 36514 18470 36566 18522
rect 36578 18470 36630 18522
rect 36642 18470 36694 18522
rect 36706 18470 36758 18522
rect 36770 18470 36822 18522
rect 67234 18470 67286 18522
rect 67298 18470 67350 18522
rect 67362 18470 67414 18522
rect 67426 18470 67478 18522
rect 67490 18470 67542 18522
rect 5134 17926 5186 17978
rect 5198 17926 5250 17978
rect 5262 17926 5314 17978
rect 5326 17926 5378 17978
rect 5390 17926 5442 17978
rect 35854 17926 35906 17978
rect 35918 17926 35970 17978
rect 35982 17926 36034 17978
rect 36046 17926 36098 17978
rect 36110 17926 36162 17978
rect 66574 17926 66626 17978
rect 66638 17926 66690 17978
rect 66702 17926 66754 17978
rect 66766 17926 66818 17978
rect 66830 17926 66882 17978
rect 29276 17824 29328 17876
rect 31116 17824 31168 17876
rect 31668 17824 31720 17876
rect 35440 17824 35492 17876
rect 5794 17382 5846 17434
rect 5858 17382 5910 17434
rect 5922 17382 5974 17434
rect 5986 17382 6038 17434
rect 6050 17382 6102 17434
rect 36514 17382 36566 17434
rect 36578 17382 36630 17434
rect 36642 17382 36694 17434
rect 36706 17382 36758 17434
rect 36770 17382 36822 17434
rect 67234 17382 67286 17434
rect 67298 17382 67350 17434
rect 67362 17382 67414 17434
rect 67426 17382 67478 17434
rect 67490 17382 67542 17434
rect 5134 16838 5186 16890
rect 5198 16838 5250 16890
rect 5262 16838 5314 16890
rect 5326 16838 5378 16890
rect 5390 16838 5442 16890
rect 35854 16838 35906 16890
rect 35918 16838 35970 16890
rect 35982 16838 36034 16890
rect 36046 16838 36098 16890
rect 36110 16838 36162 16890
rect 66574 16838 66626 16890
rect 66638 16838 66690 16890
rect 66702 16838 66754 16890
rect 66766 16838 66818 16890
rect 66830 16838 66882 16890
rect 5794 16294 5846 16346
rect 5858 16294 5910 16346
rect 5922 16294 5974 16346
rect 5986 16294 6038 16346
rect 6050 16294 6102 16346
rect 36514 16294 36566 16346
rect 36578 16294 36630 16346
rect 36642 16294 36694 16346
rect 36706 16294 36758 16346
rect 36770 16294 36822 16346
rect 67234 16294 67286 16346
rect 67298 16294 67350 16346
rect 67362 16294 67414 16346
rect 67426 16294 67478 16346
rect 67490 16294 67542 16346
rect 5134 15750 5186 15802
rect 5198 15750 5250 15802
rect 5262 15750 5314 15802
rect 5326 15750 5378 15802
rect 5390 15750 5442 15802
rect 35854 15750 35906 15802
rect 35918 15750 35970 15802
rect 35982 15750 36034 15802
rect 36046 15750 36098 15802
rect 36110 15750 36162 15802
rect 66574 15750 66626 15802
rect 66638 15750 66690 15802
rect 66702 15750 66754 15802
rect 66766 15750 66818 15802
rect 66830 15750 66882 15802
rect 5794 15206 5846 15258
rect 5858 15206 5910 15258
rect 5922 15206 5974 15258
rect 5986 15206 6038 15258
rect 6050 15206 6102 15258
rect 36514 15206 36566 15258
rect 36578 15206 36630 15258
rect 36642 15206 36694 15258
rect 36706 15206 36758 15258
rect 36770 15206 36822 15258
rect 67234 15206 67286 15258
rect 67298 15206 67350 15258
rect 67362 15206 67414 15258
rect 67426 15206 67478 15258
rect 67490 15206 67542 15258
rect 5134 14662 5186 14714
rect 5198 14662 5250 14714
rect 5262 14662 5314 14714
rect 5326 14662 5378 14714
rect 5390 14662 5442 14714
rect 35854 14662 35906 14714
rect 35918 14662 35970 14714
rect 35982 14662 36034 14714
rect 36046 14662 36098 14714
rect 36110 14662 36162 14714
rect 66574 14662 66626 14714
rect 66638 14662 66690 14714
rect 66702 14662 66754 14714
rect 66766 14662 66818 14714
rect 66830 14662 66882 14714
rect 25964 14424 26016 14476
rect 58808 14424 58860 14476
rect 5794 14118 5846 14170
rect 5858 14118 5910 14170
rect 5922 14118 5974 14170
rect 5986 14118 6038 14170
rect 6050 14118 6102 14170
rect 36514 14118 36566 14170
rect 36578 14118 36630 14170
rect 36642 14118 36694 14170
rect 36706 14118 36758 14170
rect 36770 14118 36822 14170
rect 67234 14118 67286 14170
rect 67298 14118 67350 14170
rect 67362 14118 67414 14170
rect 67426 14118 67478 14170
rect 67490 14118 67542 14170
rect 5134 13574 5186 13626
rect 5198 13574 5250 13626
rect 5262 13574 5314 13626
rect 5326 13574 5378 13626
rect 5390 13574 5442 13626
rect 35854 13574 35906 13626
rect 35918 13574 35970 13626
rect 35982 13574 36034 13626
rect 36046 13574 36098 13626
rect 36110 13574 36162 13626
rect 66574 13574 66626 13626
rect 66638 13574 66690 13626
rect 66702 13574 66754 13626
rect 66766 13574 66818 13626
rect 66830 13574 66882 13626
rect 5794 13030 5846 13082
rect 5858 13030 5910 13082
rect 5922 13030 5974 13082
rect 5986 13030 6038 13082
rect 6050 13030 6102 13082
rect 36514 13030 36566 13082
rect 36578 13030 36630 13082
rect 36642 13030 36694 13082
rect 36706 13030 36758 13082
rect 36770 13030 36822 13082
rect 67234 13030 67286 13082
rect 67298 13030 67350 13082
rect 67362 13030 67414 13082
rect 67426 13030 67478 13082
rect 67490 13030 67542 13082
rect 14188 12656 14240 12708
rect 27896 12656 27948 12708
rect 17592 12588 17644 12640
rect 38016 12588 38068 12640
rect 5134 12486 5186 12538
rect 5198 12486 5250 12538
rect 5262 12486 5314 12538
rect 5326 12486 5378 12538
rect 5390 12486 5442 12538
rect 35854 12486 35906 12538
rect 35918 12486 35970 12538
rect 35982 12486 36034 12538
rect 36046 12486 36098 12538
rect 36110 12486 36162 12538
rect 66574 12486 66626 12538
rect 66638 12486 66690 12538
rect 66702 12486 66754 12538
rect 66766 12486 66818 12538
rect 66830 12486 66882 12538
rect 25688 12044 25740 12096
rect 30840 12044 30892 12096
rect 5794 11942 5846 11994
rect 5858 11942 5910 11994
rect 5922 11942 5974 11994
rect 5986 11942 6038 11994
rect 6050 11942 6102 11994
rect 36514 11942 36566 11994
rect 36578 11942 36630 11994
rect 36642 11942 36694 11994
rect 36706 11942 36758 11994
rect 36770 11942 36822 11994
rect 67234 11942 67286 11994
rect 67298 11942 67350 11994
rect 67362 11942 67414 11994
rect 67426 11942 67478 11994
rect 67490 11942 67542 11994
rect 23112 11840 23164 11892
rect 25320 11840 25372 11892
rect 22192 11772 22244 11824
rect 27068 11772 27120 11824
rect 28080 11772 28132 11824
rect 24308 11704 24360 11756
rect 24768 11704 24820 11756
rect 26240 11704 26292 11756
rect 36360 11840 36412 11892
rect 30288 11772 30340 11824
rect 19432 11636 19484 11688
rect 23940 11636 23992 11688
rect 27252 11636 27304 11688
rect 21916 11568 21968 11620
rect 24860 11568 24912 11620
rect 25964 11568 26016 11620
rect 12992 11500 13044 11552
rect 29644 11747 29696 11756
rect 29644 11713 29653 11747
rect 29653 11713 29687 11747
rect 29687 11713 29696 11747
rect 29644 11704 29696 11713
rect 28908 11636 28960 11688
rect 29000 11568 29052 11620
rect 38844 11568 38896 11620
rect 29276 11543 29328 11552
rect 29276 11509 29285 11543
rect 29285 11509 29319 11543
rect 29319 11509 29328 11543
rect 29276 11500 29328 11509
rect 5134 11398 5186 11450
rect 5198 11398 5250 11450
rect 5262 11398 5314 11450
rect 5326 11398 5378 11450
rect 5390 11398 5442 11450
rect 35854 11398 35906 11450
rect 35918 11398 35970 11450
rect 35982 11398 36034 11450
rect 36046 11398 36098 11450
rect 36110 11398 36162 11450
rect 66574 11398 66626 11450
rect 66638 11398 66690 11450
rect 66702 11398 66754 11450
rect 66766 11398 66818 11450
rect 66830 11398 66882 11450
rect 20352 11296 20404 11348
rect 22100 11271 22152 11280
rect 22100 11237 22109 11271
rect 22109 11237 22143 11271
rect 22143 11237 22152 11271
rect 22100 11228 22152 11237
rect 16580 11160 16632 11212
rect 23388 11228 23440 11280
rect 23480 11271 23532 11280
rect 23480 11237 23489 11271
rect 23489 11237 23523 11271
rect 23523 11237 23532 11271
rect 23480 11228 23532 11237
rect 24676 11296 24728 11348
rect 20812 11092 20864 11144
rect 21916 11135 21968 11144
rect 21916 11101 21925 11135
rect 21925 11101 21959 11135
rect 21959 11101 21968 11135
rect 21916 11092 21968 11101
rect 24492 11160 24544 11212
rect 22468 11135 22520 11144
rect 22468 11101 22477 11135
rect 22477 11101 22511 11135
rect 22511 11101 22520 11135
rect 22468 11092 22520 11101
rect 22560 11092 22612 11144
rect 23940 11135 23992 11144
rect 23940 11101 23949 11135
rect 23949 11101 23983 11135
rect 23983 11101 23992 11135
rect 23940 11092 23992 11101
rect 24860 11160 24912 11212
rect 26976 11296 27028 11348
rect 27436 11296 27488 11348
rect 29000 11296 29052 11348
rect 27988 11271 28040 11280
rect 27988 11237 27997 11271
rect 27997 11237 28031 11271
rect 28031 11237 28040 11271
rect 27988 11228 28040 11237
rect 30380 11228 30432 11280
rect 28540 11203 28592 11212
rect 28540 11169 28549 11203
rect 28549 11169 28583 11203
rect 28583 11169 28592 11203
rect 28540 11160 28592 11169
rect 28724 11160 28776 11212
rect 20260 11024 20312 11076
rect 22192 11067 22244 11076
rect 22192 11033 22201 11067
rect 22201 11033 22235 11067
rect 22235 11033 22244 11067
rect 22192 11024 22244 11033
rect 24216 11024 24268 11076
rect 24676 11135 24728 11144
rect 24676 11101 24685 11135
rect 24685 11101 24719 11135
rect 24719 11101 24728 11135
rect 24676 11092 24728 11101
rect 24768 11135 24820 11144
rect 24768 11101 24777 11135
rect 24777 11101 24811 11135
rect 24811 11101 24820 11135
rect 24768 11092 24820 11101
rect 24952 11135 25004 11144
rect 24952 11101 24961 11135
rect 24961 11101 24995 11135
rect 24995 11101 25004 11135
rect 24952 11092 25004 11101
rect 25320 11092 25372 11144
rect 25688 11135 25740 11144
rect 25688 11101 25697 11135
rect 25697 11101 25731 11135
rect 25731 11101 25740 11135
rect 25688 11092 25740 11101
rect 25780 11092 25832 11144
rect 26240 11135 26292 11144
rect 26240 11101 26249 11135
rect 26249 11101 26283 11135
rect 26283 11101 26292 11135
rect 26240 11092 26292 11101
rect 26332 11135 26384 11144
rect 26332 11101 26341 11135
rect 26341 11101 26375 11135
rect 26375 11101 26384 11135
rect 26332 11092 26384 11101
rect 24860 11067 24912 11076
rect 24860 11033 24869 11067
rect 24869 11033 24903 11067
rect 24903 11033 24912 11067
rect 24860 11024 24912 11033
rect 26700 11092 26752 11144
rect 27068 11135 27120 11144
rect 27068 11101 27077 11135
rect 27077 11101 27111 11135
rect 27111 11101 27120 11135
rect 27068 11092 27120 11101
rect 27252 11135 27304 11144
rect 27252 11101 27261 11135
rect 27261 11101 27295 11135
rect 27295 11101 27304 11135
rect 27252 11092 27304 11101
rect 27344 11135 27396 11144
rect 27344 11101 27353 11135
rect 27353 11101 27387 11135
rect 27387 11101 27396 11135
rect 27344 11092 27396 11101
rect 28172 11135 28224 11144
rect 28172 11101 28181 11135
rect 28181 11101 28215 11135
rect 28215 11101 28224 11135
rect 28172 11092 28224 11101
rect 28264 11092 28316 11144
rect 29828 11135 29880 11144
rect 29828 11101 29837 11135
rect 29837 11101 29871 11135
rect 29871 11101 29880 11135
rect 29828 11092 29880 11101
rect 18236 10956 18288 11008
rect 24584 10956 24636 11008
rect 24676 10956 24728 11008
rect 24768 10956 24820 11008
rect 29184 11024 29236 11076
rect 32128 11024 32180 11076
rect 27160 10956 27212 11008
rect 29644 10956 29696 11008
rect 5794 10854 5846 10906
rect 5858 10854 5910 10906
rect 5922 10854 5974 10906
rect 5986 10854 6038 10906
rect 6050 10854 6102 10906
rect 36514 10854 36566 10906
rect 36578 10854 36630 10906
rect 36642 10854 36694 10906
rect 36706 10854 36758 10906
rect 36770 10854 36822 10906
rect 67234 10854 67286 10906
rect 67298 10854 67350 10906
rect 67362 10854 67414 10906
rect 67426 10854 67478 10906
rect 67490 10854 67542 10906
rect 20076 10752 20128 10804
rect 20720 10752 20772 10804
rect 17500 10684 17552 10736
rect 21640 10684 21692 10736
rect 22744 10752 22796 10804
rect 23020 10752 23072 10804
rect 27804 10752 27856 10804
rect 27896 10795 27948 10804
rect 27896 10761 27905 10795
rect 27905 10761 27939 10795
rect 27939 10761 27948 10795
rect 27896 10752 27948 10761
rect 28172 10752 28224 10804
rect 29644 10752 29696 10804
rect 19248 10616 19300 10668
rect 20720 10659 20772 10668
rect 20720 10625 20729 10659
rect 20729 10625 20763 10659
rect 20763 10625 20772 10659
rect 20720 10616 20772 10625
rect 21272 10659 21324 10668
rect 21272 10625 21281 10659
rect 21281 10625 21315 10659
rect 21315 10625 21324 10659
rect 21272 10616 21324 10625
rect 16672 10548 16724 10600
rect 22284 10616 22336 10668
rect 22836 10684 22888 10736
rect 23296 10684 23348 10736
rect 23388 10727 23440 10736
rect 23388 10693 23397 10727
rect 23397 10693 23431 10727
rect 23431 10693 23440 10727
rect 23388 10684 23440 10693
rect 27988 10684 28040 10736
rect 22744 10616 22796 10668
rect 27804 10616 27856 10668
rect 10508 10480 10560 10532
rect 24124 10591 24176 10600
rect 24124 10557 24133 10591
rect 24133 10557 24167 10591
rect 24167 10557 24176 10591
rect 24124 10548 24176 10557
rect 24584 10548 24636 10600
rect 25136 10548 25188 10600
rect 25412 10548 25464 10600
rect 26056 10548 26108 10600
rect 26240 10591 26292 10600
rect 26240 10557 26249 10591
rect 26249 10557 26283 10591
rect 26283 10557 26292 10591
rect 26240 10548 26292 10557
rect 26608 10548 26660 10600
rect 26884 10548 26936 10600
rect 28816 10659 28868 10668
rect 28816 10625 28825 10659
rect 28825 10625 28859 10659
rect 28859 10625 28868 10659
rect 28816 10616 28868 10625
rect 30288 10616 30340 10668
rect 31300 10752 31352 10804
rect 31208 10727 31260 10736
rect 31208 10693 31217 10727
rect 31217 10693 31251 10727
rect 31251 10693 31260 10727
rect 31208 10684 31260 10693
rect 34244 10684 34296 10736
rect 33876 10616 33928 10668
rect 34888 10659 34940 10668
rect 34888 10625 34897 10659
rect 34897 10625 34931 10659
rect 34931 10625 34940 10659
rect 34888 10616 34940 10625
rect 35164 10659 35216 10668
rect 35164 10625 35173 10659
rect 35173 10625 35207 10659
rect 35207 10625 35216 10659
rect 35164 10616 35216 10625
rect 29000 10548 29052 10600
rect 29736 10548 29788 10600
rect 31484 10548 31536 10600
rect 33140 10548 33192 10600
rect 33324 10591 33376 10600
rect 33324 10557 33333 10591
rect 33333 10557 33367 10591
rect 33367 10557 33376 10591
rect 33324 10548 33376 10557
rect 14740 10412 14792 10464
rect 21364 10455 21416 10464
rect 21364 10421 21373 10455
rect 21373 10421 21407 10455
rect 21407 10421 21416 10455
rect 21364 10412 21416 10421
rect 21548 10455 21600 10464
rect 21548 10421 21557 10455
rect 21557 10421 21591 10455
rect 21591 10421 21600 10455
rect 21548 10412 21600 10421
rect 22652 10412 22704 10464
rect 22744 10455 22796 10464
rect 22744 10421 22753 10455
rect 22753 10421 22787 10455
rect 22787 10421 22796 10455
rect 22744 10412 22796 10421
rect 23112 10455 23164 10464
rect 23112 10421 23121 10455
rect 23121 10421 23155 10455
rect 23155 10421 23164 10455
rect 23112 10412 23164 10421
rect 23204 10412 23256 10464
rect 23848 10412 23900 10464
rect 24584 10412 24636 10464
rect 24676 10412 24728 10464
rect 25412 10412 25464 10464
rect 25964 10455 26016 10464
rect 25964 10421 25973 10455
rect 25973 10421 26007 10455
rect 26007 10421 26016 10455
rect 25964 10412 26016 10421
rect 26056 10455 26108 10464
rect 26056 10421 26065 10455
rect 26065 10421 26099 10455
rect 26099 10421 26108 10455
rect 26056 10412 26108 10421
rect 26608 10412 26660 10464
rect 27528 10455 27580 10464
rect 27528 10421 27537 10455
rect 27537 10421 27571 10455
rect 27571 10421 27580 10455
rect 27528 10412 27580 10421
rect 28632 10455 28684 10464
rect 28632 10421 28641 10455
rect 28641 10421 28675 10455
rect 28675 10421 28684 10455
rect 28632 10412 28684 10421
rect 28816 10412 28868 10464
rect 31668 10480 31720 10532
rect 33600 10548 33652 10600
rect 30196 10455 30248 10464
rect 30196 10421 30205 10455
rect 30205 10421 30239 10455
rect 30239 10421 30248 10455
rect 30196 10412 30248 10421
rect 32312 10412 32364 10464
rect 32496 10412 32548 10464
rect 34796 10412 34848 10464
rect 35440 10455 35492 10464
rect 35440 10421 35449 10455
rect 35449 10421 35483 10455
rect 35483 10421 35492 10455
rect 35440 10412 35492 10421
rect 5134 10310 5186 10362
rect 5198 10310 5250 10362
rect 5262 10310 5314 10362
rect 5326 10310 5378 10362
rect 5390 10310 5442 10362
rect 35854 10310 35906 10362
rect 35918 10310 35970 10362
rect 35982 10310 36034 10362
rect 36046 10310 36098 10362
rect 36110 10310 36162 10362
rect 66574 10310 66626 10362
rect 66638 10310 66690 10362
rect 66702 10310 66754 10362
rect 66766 10310 66818 10362
rect 66830 10310 66882 10362
rect 19892 10208 19944 10260
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 16856 10140 16908 10192
rect 21456 10208 21508 10260
rect 23204 10208 23256 10260
rect 23296 10208 23348 10260
rect 24676 10208 24728 10260
rect 27160 10208 27212 10260
rect 27436 10208 27488 10260
rect 28540 10251 28592 10260
rect 28540 10217 28549 10251
rect 28549 10217 28583 10251
rect 28583 10217 28592 10251
rect 28540 10208 28592 10217
rect 30288 10208 30340 10260
rect 34336 10208 34388 10260
rect 20812 10072 20864 10124
rect 19432 10004 19484 10056
rect 19708 10047 19760 10056
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 13728 9936 13780 9988
rect 20904 10047 20956 10056
rect 20904 10013 20913 10047
rect 20913 10013 20947 10047
rect 20947 10013 20956 10047
rect 20904 10004 20956 10013
rect 20536 9911 20588 9920
rect 20536 9877 20545 9911
rect 20545 9877 20579 9911
rect 20579 9877 20588 9911
rect 20536 9868 20588 9877
rect 21088 9936 21140 9988
rect 21456 10072 21508 10124
rect 21824 10004 21876 10056
rect 22652 10115 22704 10124
rect 22652 10081 22661 10115
rect 22661 10081 22695 10115
rect 22695 10081 22704 10115
rect 22652 10072 22704 10081
rect 22744 10004 22796 10056
rect 22928 10004 22980 10056
rect 23848 10072 23900 10124
rect 37188 10140 37240 10192
rect 31208 10115 31260 10124
rect 31208 10081 31217 10115
rect 31217 10081 31251 10115
rect 31251 10081 31260 10115
rect 31208 10072 31260 10081
rect 23480 10047 23532 10056
rect 23480 10013 23489 10047
rect 23489 10013 23523 10047
rect 23523 10013 23532 10047
rect 23480 10004 23532 10013
rect 24124 10047 24176 10056
rect 24124 10013 24133 10047
rect 24133 10013 24167 10047
rect 24167 10013 24176 10047
rect 24124 10004 24176 10013
rect 25136 10004 25188 10056
rect 25504 10047 25556 10056
rect 25504 10013 25513 10047
rect 25513 10013 25547 10047
rect 25547 10013 25556 10047
rect 25504 10004 25556 10013
rect 25596 10004 25648 10056
rect 22008 9936 22060 9988
rect 23296 9936 23348 9988
rect 26056 10004 26108 10056
rect 26608 10004 26660 10056
rect 27344 10004 27396 10056
rect 27804 10047 27856 10056
rect 27804 10013 27813 10047
rect 27813 10013 27847 10047
rect 27847 10013 27856 10047
rect 27804 10004 27856 10013
rect 29460 10004 29512 10056
rect 25872 9979 25924 9988
rect 25872 9945 25881 9979
rect 25881 9945 25915 9979
rect 25915 9945 25924 9979
rect 25872 9936 25924 9945
rect 29552 9936 29604 9988
rect 32956 10072 33008 10124
rect 34796 10115 34848 10124
rect 34796 10081 34805 10115
rect 34805 10081 34839 10115
rect 34839 10081 34848 10115
rect 34796 10072 34848 10081
rect 31852 10047 31904 10056
rect 31852 10013 31861 10047
rect 31861 10013 31895 10047
rect 31895 10013 31904 10047
rect 31852 10004 31904 10013
rect 32588 10004 32640 10056
rect 32864 10004 32916 10056
rect 35624 10047 35676 10056
rect 35624 10013 35633 10047
rect 35633 10013 35667 10047
rect 35667 10013 35676 10047
rect 35624 10004 35676 10013
rect 36912 10004 36964 10056
rect 32404 9936 32456 9988
rect 21364 9911 21416 9920
rect 21364 9877 21373 9911
rect 21373 9877 21407 9911
rect 21407 9877 21416 9911
rect 21364 9868 21416 9877
rect 22100 9911 22152 9920
rect 22100 9877 22109 9911
rect 22109 9877 22143 9911
rect 22143 9877 22152 9911
rect 22100 9868 22152 9877
rect 22376 9868 22428 9920
rect 23112 9868 23164 9920
rect 23480 9868 23532 9920
rect 25044 9868 25096 9920
rect 25228 9868 25280 9920
rect 25412 9868 25464 9920
rect 26056 9868 26108 9920
rect 26148 9911 26200 9920
rect 26148 9877 26157 9911
rect 26157 9877 26191 9911
rect 26191 9877 26200 9911
rect 26148 9868 26200 9877
rect 28632 9911 28684 9920
rect 28632 9877 28641 9911
rect 28641 9877 28675 9911
rect 28675 9877 28684 9911
rect 28632 9868 28684 9877
rect 29000 9911 29052 9920
rect 29000 9877 29009 9911
rect 29009 9877 29043 9911
rect 29043 9877 29052 9911
rect 29000 9868 29052 9877
rect 30012 9868 30064 9920
rect 30472 9911 30524 9920
rect 30472 9877 30481 9911
rect 30481 9877 30515 9911
rect 30515 9877 30524 9911
rect 30472 9868 30524 9877
rect 32680 9868 32732 9920
rect 33416 9868 33468 9920
rect 36268 9911 36320 9920
rect 36268 9877 36277 9911
rect 36277 9877 36311 9911
rect 36311 9877 36320 9911
rect 36268 9868 36320 9877
rect 38752 9868 38804 9920
rect 5794 9766 5846 9818
rect 5858 9766 5910 9818
rect 5922 9766 5974 9818
rect 5986 9766 6038 9818
rect 6050 9766 6102 9818
rect 36514 9766 36566 9818
rect 36578 9766 36630 9818
rect 36642 9766 36694 9818
rect 36706 9766 36758 9818
rect 36770 9766 36822 9818
rect 67234 9766 67286 9818
rect 67298 9766 67350 9818
rect 67362 9766 67414 9818
rect 67426 9766 67478 9818
rect 67490 9766 67542 9818
rect 15568 9596 15620 9648
rect 18880 9596 18932 9648
rect 19340 9596 19392 9648
rect 18696 9571 18748 9580
rect 18696 9537 18705 9571
rect 18705 9537 18739 9571
rect 18739 9537 18748 9571
rect 18696 9528 18748 9537
rect 19156 9571 19208 9580
rect 19156 9537 19165 9571
rect 19165 9537 19199 9571
rect 19199 9537 19208 9571
rect 19156 9528 19208 9537
rect 19432 9571 19484 9614
rect 19432 9562 19435 9571
rect 19435 9562 19469 9571
rect 19469 9562 19484 9571
rect 19616 9562 19668 9614
rect 23572 9664 23624 9716
rect 24124 9707 24176 9716
rect 24124 9673 24133 9707
rect 24133 9673 24167 9707
rect 24167 9673 24176 9707
rect 24124 9664 24176 9673
rect 22560 9639 22612 9648
rect 22560 9605 22569 9639
rect 22569 9605 22603 9639
rect 22603 9605 22612 9639
rect 22560 9596 22612 9605
rect 19064 9460 19116 9512
rect 19984 9528 20036 9580
rect 21824 9460 21876 9512
rect 22008 9571 22060 9580
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 24492 9596 24544 9648
rect 24676 9596 24728 9648
rect 27804 9664 27856 9716
rect 33324 9664 33376 9716
rect 26516 9596 26568 9648
rect 26884 9596 26936 9648
rect 27712 9596 27764 9648
rect 22836 9571 22888 9580
rect 22836 9537 22845 9571
rect 22845 9537 22879 9571
rect 22879 9537 22888 9571
rect 22836 9528 22888 9537
rect 23020 9571 23072 9580
rect 23020 9537 23029 9571
rect 23029 9537 23063 9571
rect 23063 9537 23072 9571
rect 23020 9528 23072 9537
rect 25964 9571 26016 9580
rect 25964 9537 25973 9571
rect 25973 9537 26007 9571
rect 26007 9537 26016 9571
rect 25964 9528 26016 9537
rect 28540 9596 28592 9648
rect 30656 9596 30708 9648
rect 31576 9596 31628 9648
rect 32864 9639 32916 9648
rect 32864 9605 32873 9639
rect 32873 9605 32907 9639
rect 32907 9605 32916 9639
rect 32864 9596 32916 9605
rect 23296 9460 23348 9512
rect 13820 9324 13872 9376
rect 20996 9324 21048 9376
rect 21732 9392 21784 9444
rect 23112 9392 23164 9444
rect 25228 9460 25280 9512
rect 25504 9460 25556 9512
rect 27160 9503 27212 9512
rect 27160 9469 27169 9503
rect 27169 9469 27203 9503
rect 27203 9469 27212 9503
rect 27160 9460 27212 9469
rect 33048 9571 33100 9580
rect 33048 9537 33057 9571
rect 33057 9537 33091 9571
rect 33091 9537 33100 9571
rect 33048 9528 33100 9537
rect 33232 9528 33284 9580
rect 33508 9528 33560 9580
rect 36268 9528 36320 9580
rect 38752 9571 38804 9580
rect 38752 9537 38761 9571
rect 38761 9537 38795 9571
rect 38795 9537 38804 9571
rect 38752 9528 38804 9537
rect 24216 9435 24268 9444
rect 24216 9401 24225 9435
rect 24225 9401 24259 9435
rect 24259 9401 24268 9435
rect 24216 9392 24268 9401
rect 24676 9435 24728 9444
rect 24676 9401 24685 9435
rect 24685 9401 24719 9435
rect 24719 9401 24728 9435
rect 24676 9392 24728 9401
rect 23204 9367 23256 9376
rect 23204 9333 23213 9367
rect 23213 9333 23247 9367
rect 23247 9333 23256 9367
rect 23204 9324 23256 9333
rect 23296 9367 23348 9376
rect 23296 9333 23305 9367
rect 23305 9333 23339 9367
rect 23339 9333 23348 9367
rect 23296 9324 23348 9333
rect 23572 9324 23624 9376
rect 23848 9324 23900 9376
rect 25320 9324 25372 9376
rect 28448 9392 28500 9444
rect 28632 9460 28684 9512
rect 29644 9460 29696 9512
rect 30932 9460 30984 9512
rect 31300 9503 31352 9512
rect 31300 9469 31309 9503
rect 31309 9469 31343 9503
rect 31343 9469 31352 9503
rect 31300 9460 31352 9469
rect 31576 9460 31628 9512
rect 32036 9503 32088 9512
rect 32036 9469 32045 9503
rect 32045 9469 32079 9503
rect 32079 9469 32088 9503
rect 32036 9460 32088 9469
rect 32220 9503 32272 9512
rect 32220 9469 32229 9503
rect 32229 9469 32263 9503
rect 32263 9469 32272 9503
rect 32220 9460 32272 9469
rect 29000 9392 29052 9444
rect 29092 9392 29144 9444
rect 28356 9324 28408 9376
rect 29184 9324 29236 9376
rect 30748 9367 30800 9376
rect 30748 9333 30757 9367
rect 30757 9333 30791 9367
rect 30791 9333 30800 9367
rect 30748 9324 30800 9333
rect 31392 9324 31444 9376
rect 34980 9503 35032 9512
rect 34980 9469 34989 9503
rect 34989 9469 35023 9503
rect 35023 9469 35032 9503
rect 34980 9460 35032 9469
rect 36360 9460 36412 9512
rect 37924 9460 37976 9512
rect 32772 9324 32824 9376
rect 35072 9392 35124 9444
rect 35348 9392 35400 9444
rect 37096 9392 37148 9444
rect 34152 9324 34204 9376
rect 35256 9367 35308 9376
rect 35256 9333 35265 9367
rect 35265 9333 35299 9367
rect 35299 9333 35308 9367
rect 35256 9324 35308 9333
rect 37004 9324 37056 9376
rect 38200 9367 38252 9376
rect 38200 9333 38209 9367
rect 38209 9333 38243 9367
rect 38243 9333 38252 9367
rect 38200 9324 38252 9333
rect 5134 9222 5186 9274
rect 5198 9222 5250 9274
rect 5262 9222 5314 9274
rect 5326 9222 5378 9274
rect 5390 9222 5442 9274
rect 35854 9222 35906 9274
rect 35918 9222 35970 9274
rect 35982 9222 36034 9274
rect 36046 9222 36098 9274
rect 36110 9222 36162 9274
rect 66574 9222 66626 9274
rect 66638 9222 66690 9274
rect 66702 9222 66754 9274
rect 66766 9222 66818 9274
rect 66830 9222 66882 9274
rect 11796 9163 11848 9172
rect 11796 9129 11805 9163
rect 11805 9129 11839 9163
rect 11839 9129 11848 9163
rect 11796 9120 11848 9129
rect 15936 9120 15988 9172
rect 17592 9163 17644 9172
rect 17592 9129 17601 9163
rect 17601 9129 17635 9163
rect 17635 9129 17644 9163
rect 17592 9120 17644 9129
rect 17684 9120 17736 9172
rect 18972 9052 19024 9104
rect 10876 8984 10928 9036
rect 17776 8984 17828 9036
rect 9956 8916 10008 8968
rect 17960 8916 18012 8968
rect 18052 8891 18104 8900
rect 18052 8857 18061 8891
rect 18061 8857 18095 8891
rect 18095 8857 18104 8891
rect 18052 8848 18104 8857
rect 18144 8848 18196 8900
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 19616 8848 19668 8900
rect 20260 8916 20312 8968
rect 23204 9120 23256 9172
rect 21916 9052 21968 9104
rect 23296 9052 23348 9104
rect 22100 8984 22152 9036
rect 22928 8984 22980 9036
rect 23572 9027 23624 9036
rect 23572 8993 23581 9027
rect 23581 8993 23615 9027
rect 23615 8993 23624 9027
rect 23572 8984 23624 8993
rect 18420 8780 18472 8832
rect 18604 8823 18656 8832
rect 18604 8789 18613 8823
rect 18613 8789 18647 8823
rect 18647 8789 18656 8823
rect 18604 8780 18656 8789
rect 19524 8780 19576 8832
rect 20168 8780 20220 8832
rect 20260 8823 20312 8832
rect 20260 8789 20269 8823
rect 20269 8789 20303 8823
rect 20303 8789 20312 8823
rect 20260 8780 20312 8789
rect 20444 8891 20496 8900
rect 20444 8857 20453 8891
rect 20453 8857 20487 8891
rect 20487 8857 20496 8891
rect 20444 8848 20496 8857
rect 20812 8848 20864 8900
rect 21548 8848 21600 8900
rect 24308 8959 24360 8968
rect 24308 8925 24317 8959
rect 24317 8925 24351 8959
rect 24351 8925 24360 8959
rect 24308 8916 24360 8925
rect 24492 8959 24544 8968
rect 24492 8925 24501 8959
rect 24501 8925 24535 8959
rect 24535 8925 24544 8959
rect 24492 8916 24544 8925
rect 25136 8916 25188 8968
rect 25688 9120 25740 9172
rect 32864 9120 32916 9172
rect 33140 9120 33192 9172
rect 33508 9120 33560 9172
rect 35624 9120 35676 9172
rect 25964 9052 26016 9104
rect 27528 8984 27580 9036
rect 28448 8984 28500 9036
rect 29276 8984 29328 9036
rect 27712 8959 27764 8968
rect 27712 8925 27721 8959
rect 27721 8925 27755 8959
rect 27755 8925 27764 8959
rect 27712 8916 27764 8925
rect 30472 8984 30524 9036
rect 29644 8959 29696 8968
rect 29644 8925 29653 8959
rect 29653 8925 29687 8959
rect 29687 8925 29696 8959
rect 29644 8916 29696 8925
rect 31944 9052 31996 9104
rect 36084 9052 36136 9104
rect 36452 9052 36504 9104
rect 34060 8984 34112 9036
rect 31852 8916 31904 8968
rect 32404 8959 32456 8968
rect 32404 8925 32413 8959
rect 32413 8925 32447 8959
rect 32447 8925 32456 8959
rect 32404 8916 32456 8925
rect 33140 8959 33192 8968
rect 33140 8925 33149 8959
rect 33149 8925 33183 8959
rect 33183 8925 33192 8959
rect 33140 8916 33192 8925
rect 34520 8916 34572 8968
rect 35072 8916 35124 8968
rect 35440 8984 35492 9036
rect 38292 8984 38344 9036
rect 27436 8848 27488 8900
rect 29000 8848 29052 8900
rect 30472 8848 30524 8900
rect 31116 8848 31168 8900
rect 31668 8891 31720 8900
rect 31668 8857 31677 8891
rect 31677 8857 31711 8891
rect 31711 8857 31720 8891
rect 31668 8848 31720 8857
rect 20720 8780 20772 8832
rect 21456 8780 21508 8832
rect 23480 8780 23532 8832
rect 25044 8780 25096 8832
rect 25228 8780 25280 8832
rect 27252 8780 27304 8832
rect 28448 8823 28500 8832
rect 28448 8789 28457 8823
rect 28457 8789 28491 8823
rect 28491 8789 28500 8823
rect 28448 8780 28500 8789
rect 29368 8780 29420 8832
rect 31760 8823 31812 8832
rect 31760 8789 31769 8823
rect 31769 8789 31803 8823
rect 31803 8789 31812 8823
rect 31760 8780 31812 8789
rect 31944 8780 31996 8832
rect 32404 8780 32456 8832
rect 33324 8823 33376 8832
rect 33324 8789 33333 8823
rect 33333 8789 33367 8823
rect 33367 8789 33376 8823
rect 33324 8780 33376 8789
rect 33508 8848 33560 8900
rect 36268 8848 36320 8900
rect 33876 8780 33928 8832
rect 34520 8780 34572 8832
rect 35072 8780 35124 8832
rect 35716 8780 35768 8832
rect 37464 8916 37516 8968
rect 37372 8891 37424 8900
rect 37372 8857 37381 8891
rect 37381 8857 37415 8891
rect 37415 8857 37424 8891
rect 37372 8848 37424 8857
rect 38660 8823 38712 8832
rect 38660 8789 38669 8823
rect 38669 8789 38703 8823
rect 38703 8789 38712 8823
rect 38660 8780 38712 8789
rect 5794 8678 5846 8730
rect 5858 8678 5910 8730
rect 5922 8678 5974 8730
rect 5986 8678 6038 8730
rect 6050 8678 6102 8730
rect 36514 8678 36566 8730
rect 36578 8678 36630 8730
rect 36642 8678 36694 8730
rect 36706 8678 36758 8730
rect 36770 8678 36822 8730
rect 67234 8678 67286 8730
rect 67298 8678 67350 8730
rect 67362 8678 67414 8730
rect 67426 8678 67478 8730
rect 67490 8678 67542 8730
rect 15108 8576 15160 8628
rect 18144 8576 18196 8628
rect 19248 8619 19300 8628
rect 19248 8585 19257 8619
rect 19257 8585 19291 8619
rect 19291 8585 19300 8619
rect 19248 8576 19300 8585
rect 19432 8576 19484 8628
rect 13912 8508 13964 8560
rect 19892 8508 19944 8560
rect 8208 8440 8260 8492
rect 16120 8440 16172 8492
rect 23296 8576 23348 8628
rect 12900 8372 12952 8424
rect 3976 8304 4028 8356
rect 17132 8372 17184 8424
rect 16396 8304 16448 8356
rect 18144 8372 18196 8424
rect 18880 8372 18932 8424
rect 19340 8372 19392 8424
rect 17316 8347 17368 8356
rect 17316 8313 17325 8347
rect 17325 8313 17359 8347
rect 17359 8313 17368 8347
rect 17316 8304 17368 8313
rect 19248 8304 19300 8356
rect 19432 8347 19484 8356
rect 19432 8313 19441 8347
rect 19441 8313 19475 8347
rect 19475 8313 19484 8347
rect 19432 8304 19484 8313
rect 21916 8508 21968 8560
rect 22008 8508 22060 8560
rect 23664 8508 23716 8560
rect 21640 8440 21692 8492
rect 22100 8440 22152 8492
rect 22376 8440 22428 8492
rect 25780 8576 25832 8628
rect 29644 8576 29696 8628
rect 30196 8576 30248 8628
rect 25872 8508 25924 8560
rect 26884 8508 26936 8560
rect 27804 8440 27856 8492
rect 20444 8415 20496 8424
rect 20444 8381 20453 8415
rect 20453 8381 20487 8415
rect 20487 8381 20496 8415
rect 20444 8372 20496 8381
rect 20812 8372 20864 8424
rect 21916 8415 21968 8424
rect 21916 8381 21925 8415
rect 21925 8381 21959 8415
rect 21959 8381 21968 8415
rect 21916 8372 21968 8381
rect 23388 8372 23440 8424
rect 24032 8415 24084 8424
rect 24032 8381 24041 8415
rect 24041 8381 24075 8415
rect 24075 8381 24084 8415
rect 24032 8372 24084 8381
rect 24308 8415 24360 8424
rect 24308 8381 24317 8415
rect 24317 8381 24351 8415
rect 24351 8381 24360 8415
rect 24308 8372 24360 8381
rect 24676 8372 24728 8424
rect 25688 8372 25740 8424
rect 26056 8415 26108 8424
rect 26056 8381 26065 8415
rect 26065 8381 26099 8415
rect 26099 8381 26108 8415
rect 26056 8372 26108 8381
rect 26424 8372 26476 8424
rect 26976 8415 27028 8424
rect 26976 8381 26985 8415
rect 26985 8381 27019 8415
rect 27019 8381 27028 8415
rect 26976 8372 27028 8381
rect 21088 8347 21140 8356
rect 21088 8313 21097 8347
rect 21097 8313 21131 8347
rect 21131 8313 21140 8347
rect 21088 8304 21140 8313
rect 21180 8347 21232 8356
rect 21180 8313 21189 8347
rect 21189 8313 21223 8347
rect 21223 8313 21232 8347
rect 21180 8304 21232 8313
rect 19800 8236 19852 8288
rect 22376 8236 22428 8288
rect 23756 8304 23808 8356
rect 23940 8236 23992 8288
rect 25596 8304 25648 8356
rect 28172 8415 28224 8424
rect 28172 8381 28181 8415
rect 28181 8381 28215 8415
rect 28215 8381 28224 8415
rect 28172 8372 28224 8381
rect 27252 8304 27304 8356
rect 27896 8347 27948 8356
rect 27896 8313 27905 8347
rect 27905 8313 27939 8347
rect 27939 8313 27948 8347
rect 27896 8304 27948 8313
rect 28080 8304 28132 8356
rect 29644 8415 29696 8424
rect 29644 8381 29653 8415
rect 29653 8381 29687 8415
rect 29687 8381 29696 8415
rect 29644 8372 29696 8381
rect 29920 8415 29972 8424
rect 29920 8381 29929 8415
rect 29929 8381 29963 8415
rect 29963 8381 29972 8415
rect 29920 8372 29972 8381
rect 30656 8372 30708 8424
rect 31944 8440 31996 8492
rect 32220 8415 32272 8424
rect 32220 8381 32229 8415
rect 32229 8381 32263 8415
rect 32263 8381 32272 8415
rect 32220 8372 32272 8381
rect 32404 8576 32456 8628
rect 33140 8508 33192 8560
rect 33048 8483 33100 8492
rect 33048 8449 33057 8483
rect 33057 8449 33091 8483
rect 33091 8449 33100 8483
rect 33048 8440 33100 8449
rect 32404 8372 32456 8424
rect 33508 8483 33560 8492
rect 33508 8449 33517 8483
rect 33517 8449 33551 8483
rect 33551 8449 33560 8483
rect 33508 8440 33560 8449
rect 34152 8508 34204 8560
rect 34796 8508 34848 8560
rect 35072 8551 35124 8560
rect 35072 8517 35081 8551
rect 35081 8517 35115 8551
rect 35115 8517 35124 8551
rect 35072 8508 35124 8517
rect 33784 8483 33836 8492
rect 33784 8449 33793 8483
rect 33793 8449 33827 8483
rect 33827 8449 33836 8483
rect 33784 8440 33836 8449
rect 33876 8440 33928 8492
rect 34428 8440 34480 8492
rect 36084 8440 36136 8492
rect 36728 8440 36780 8492
rect 26700 8236 26752 8288
rect 31116 8304 31168 8356
rect 34612 8415 34664 8424
rect 34612 8381 34621 8415
rect 34621 8381 34655 8415
rect 34655 8381 34664 8415
rect 34612 8372 34664 8381
rect 33876 8304 33928 8356
rect 34152 8304 34204 8356
rect 35072 8372 35124 8424
rect 35716 8372 35768 8424
rect 35808 8372 35860 8424
rect 37188 8372 37240 8424
rect 39304 8415 39356 8424
rect 39304 8381 39313 8415
rect 39313 8381 39347 8415
rect 39347 8381 39356 8415
rect 39304 8372 39356 8381
rect 37648 8304 37700 8356
rect 41420 8304 41472 8356
rect 31208 8236 31260 8288
rect 31668 8236 31720 8288
rect 33324 8236 33376 8288
rect 37556 8279 37608 8288
rect 37556 8245 37565 8279
rect 37565 8245 37599 8279
rect 37599 8245 37608 8279
rect 37556 8236 37608 8245
rect 5134 8134 5186 8186
rect 5198 8134 5250 8186
rect 5262 8134 5314 8186
rect 5326 8134 5378 8186
rect 5390 8134 5442 8186
rect 35854 8134 35906 8186
rect 35918 8134 35970 8186
rect 35982 8134 36034 8186
rect 36046 8134 36098 8186
rect 36110 8134 36162 8186
rect 66574 8134 66626 8186
rect 66638 8134 66690 8186
rect 66702 8134 66754 8186
rect 66766 8134 66818 8186
rect 66830 8134 66882 8186
rect 17960 8032 18012 8084
rect 19156 8032 19208 8084
rect 19800 8032 19852 8084
rect 21916 8032 21968 8084
rect 22192 8032 22244 8084
rect 22468 8032 22520 8084
rect 26516 8032 26568 8084
rect 27528 8032 27580 8084
rect 11152 7896 11204 7948
rect 18328 7896 18380 7948
rect 19432 7896 19484 7948
rect 6920 7828 6972 7880
rect 15384 7871 15436 7880
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 17408 7828 17460 7880
rect 18788 7871 18840 7880
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 23572 7964 23624 8016
rect 23940 7964 23992 8016
rect 24216 7964 24268 8016
rect 24768 7964 24820 8016
rect 25504 7964 25556 8016
rect 28264 7964 28316 8016
rect 29552 8007 29604 8016
rect 29552 7973 29561 8007
rect 29561 7973 29595 8007
rect 29595 7973 29604 8007
rect 29552 7964 29604 7973
rect 21640 7896 21692 7948
rect 21732 7939 21784 7948
rect 21732 7905 21741 7939
rect 21741 7905 21775 7939
rect 21775 7905 21784 7939
rect 21732 7896 21784 7905
rect 24032 7896 24084 7948
rect 24124 7939 24176 7948
rect 24124 7905 24133 7939
rect 24133 7905 24167 7939
rect 24167 7905 24176 7939
rect 24124 7896 24176 7905
rect 18604 7760 18656 7812
rect 23940 7828 23992 7880
rect 25872 7896 25924 7948
rect 26700 7896 26752 7948
rect 25044 7871 25096 7880
rect 25044 7837 25053 7871
rect 25053 7837 25087 7871
rect 25087 7837 25096 7871
rect 25044 7828 25096 7837
rect 26056 7828 26108 7880
rect 27528 7828 27580 7880
rect 27620 7871 27672 7880
rect 27620 7837 27629 7871
rect 27629 7837 27663 7871
rect 27663 7837 27672 7871
rect 27620 7828 27672 7837
rect 27804 7871 27856 7880
rect 27804 7837 27813 7871
rect 27813 7837 27847 7871
rect 27847 7837 27856 7871
rect 27804 7828 27856 7837
rect 28816 7939 28868 7948
rect 28816 7905 28825 7939
rect 28825 7905 28859 7939
rect 28859 7905 28868 7939
rect 28816 7896 28868 7905
rect 29092 7896 29144 7948
rect 29920 8032 29972 8084
rect 30380 8032 30432 8084
rect 30196 7964 30248 8016
rect 34888 8032 34940 8084
rect 37556 8032 37608 8084
rect 30840 7964 30892 8016
rect 22376 7803 22428 7812
rect 22376 7769 22385 7803
rect 22385 7769 22419 7803
rect 22419 7769 22428 7803
rect 22376 7760 22428 7769
rect 23664 7760 23716 7812
rect 10232 7692 10284 7744
rect 14832 7692 14884 7744
rect 18236 7735 18288 7744
rect 18236 7701 18245 7735
rect 18245 7701 18279 7735
rect 18279 7701 18288 7735
rect 18236 7692 18288 7701
rect 19800 7735 19852 7744
rect 19800 7701 19809 7735
rect 19809 7701 19843 7735
rect 19843 7701 19852 7735
rect 19800 7692 19852 7701
rect 21824 7692 21876 7744
rect 25688 7760 25740 7812
rect 28540 7828 28592 7880
rect 30656 7871 30708 7880
rect 30656 7837 30665 7871
rect 30665 7837 30699 7871
rect 30699 7837 30708 7871
rect 30656 7828 30708 7837
rect 31208 7828 31260 7880
rect 31392 7828 31444 7880
rect 31760 7871 31812 7880
rect 31760 7837 31769 7871
rect 31769 7837 31803 7871
rect 31803 7837 31812 7871
rect 31760 7828 31812 7837
rect 29552 7760 29604 7812
rect 29920 7760 29972 7812
rect 33508 7896 33560 7948
rect 33876 7939 33928 7948
rect 33876 7905 33885 7939
rect 33885 7905 33919 7939
rect 33919 7905 33928 7939
rect 33876 7896 33928 7905
rect 34152 7939 34204 7948
rect 34152 7905 34161 7939
rect 34161 7905 34195 7939
rect 34195 7905 34204 7939
rect 34152 7896 34204 7905
rect 24768 7692 24820 7744
rect 27160 7692 27212 7744
rect 27988 7692 28040 7744
rect 29092 7692 29144 7744
rect 30196 7692 30248 7744
rect 30288 7692 30340 7744
rect 30840 7692 30892 7744
rect 31392 7692 31444 7744
rect 32404 7760 32456 7812
rect 32312 7692 32364 7744
rect 34336 7828 34388 7880
rect 34796 7871 34848 7880
rect 34796 7837 34805 7871
rect 34805 7837 34839 7871
rect 34839 7837 34848 7871
rect 34796 7828 34848 7837
rect 34888 7828 34940 7880
rect 34428 7760 34480 7812
rect 40408 7896 40460 7948
rect 38200 7828 38252 7880
rect 35992 7803 36044 7812
rect 35992 7769 36001 7803
rect 36001 7769 36035 7803
rect 36035 7769 36044 7803
rect 35992 7760 36044 7769
rect 34336 7735 34388 7744
rect 34336 7701 34345 7735
rect 34345 7701 34379 7735
rect 34379 7701 34388 7735
rect 34336 7692 34388 7701
rect 35624 7692 35676 7744
rect 36728 7692 36780 7744
rect 38384 7760 38436 7812
rect 41604 7828 41656 7880
rect 40868 7760 40920 7812
rect 37464 7692 37516 7744
rect 39212 7692 39264 7744
rect 40132 7735 40184 7744
rect 40132 7701 40141 7735
rect 40141 7701 40175 7735
rect 40175 7701 40184 7735
rect 40132 7692 40184 7701
rect 40500 7735 40552 7744
rect 40500 7701 40509 7735
rect 40509 7701 40543 7735
rect 40543 7701 40552 7735
rect 40500 7692 40552 7701
rect 5794 7590 5846 7642
rect 5858 7590 5910 7642
rect 5922 7590 5974 7642
rect 5986 7590 6038 7642
rect 6050 7590 6102 7642
rect 36514 7590 36566 7642
rect 36578 7590 36630 7642
rect 36642 7590 36694 7642
rect 36706 7590 36758 7642
rect 36770 7590 36822 7642
rect 67234 7590 67286 7642
rect 67298 7590 67350 7642
rect 67362 7590 67414 7642
rect 67426 7590 67478 7642
rect 67490 7590 67542 7642
rect 10784 7488 10836 7540
rect 11060 7352 11112 7404
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 14464 7352 14516 7404
rect 16304 7488 16356 7540
rect 22284 7488 22336 7540
rect 23388 7531 23440 7540
rect 23388 7497 23397 7531
rect 23397 7497 23431 7531
rect 23431 7497 23440 7531
rect 23388 7488 23440 7497
rect 16488 7420 16540 7472
rect 15476 7352 15528 7404
rect 19708 7420 19760 7472
rect 20720 7352 20772 7404
rect 21824 7420 21876 7472
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 15200 7216 15252 7268
rect 12348 7148 12400 7200
rect 14556 7191 14608 7200
rect 14556 7157 14565 7191
rect 14565 7157 14599 7191
rect 14599 7157 14608 7191
rect 14556 7148 14608 7157
rect 15016 7148 15068 7200
rect 15476 7148 15528 7200
rect 15844 7148 15896 7200
rect 16028 7191 16080 7200
rect 16028 7157 16037 7191
rect 16037 7157 16071 7191
rect 16071 7157 16080 7191
rect 16028 7148 16080 7157
rect 16212 7148 16264 7200
rect 19432 7284 19484 7336
rect 20628 7284 20680 7336
rect 21456 7395 21508 7404
rect 21456 7361 21465 7395
rect 21465 7361 21499 7395
rect 21499 7361 21508 7395
rect 21456 7352 21508 7361
rect 21548 7395 21600 7404
rect 21548 7361 21557 7395
rect 21557 7361 21591 7395
rect 21591 7361 21600 7395
rect 21548 7352 21600 7361
rect 21640 7395 21692 7404
rect 21640 7361 21654 7395
rect 21654 7361 21688 7395
rect 21688 7361 21692 7395
rect 21640 7352 21692 7361
rect 21732 7284 21784 7336
rect 22008 7327 22060 7336
rect 22008 7293 22017 7327
rect 22017 7293 22051 7327
rect 22051 7293 22060 7327
rect 22008 7284 22060 7293
rect 22560 7284 22612 7336
rect 23020 7420 23072 7472
rect 27620 7488 27672 7540
rect 29828 7488 29880 7540
rect 30196 7488 30248 7540
rect 31668 7488 31720 7540
rect 32220 7531 32272 7540
rect 32220 7497 32229 7531
rect 32229 7497 32263 7531
rect 32263 7497 32272 7531
rect 32220 7488 32272 7497
rect 32864 7488 32916 7540
rect 33048 7488 33100 7540
rect 34612 7488 34664 7540
rect 36268 7488 36320 7540
rect 24492 7420 24544 7472
rect 26792 7420 26844 7472
rect 26424 7352 26476 7404
rect 26976 7352 27028 7404
rect 27436 7463 27488 7472
rect 27436 7429 27445 7463
rect 27445 7429 27479 7463
rect 27479 7429 27488 7463
rect 27436 7420 27488 7429
rect 27528 7463 27580 7472
rect 27528 7429 27537 7463
rect 27537 7429 27571 7463
rect 27571 7429 27580 7463
rect 27528 7420 27580 7429
rect 29644 7420 29696 7472
rect 28172 7352 28224 7404
rect 28724 7352 28776 7404
rect 30288 7420 30340 7472
rect 31392 7420 31444 7472
rect 31116 7352 31168 7404
rect 31668 7352 31720 7404
rect 32312 7352 32364 7404
rect 32496 7395 32548 7404
rect 32496 7361 32505 7395
rect 32505 7361 32539 7395
rect 32539 7361 32548 7395
rect 32496 7352 32548 7361
rect 33140 7420 33192 7472
rect 33232 7352 33284 7404
rect 33508 7352 33560 7404
rect 34060 7395 34112 7404
rect 34060 7361 34069 7395
rect 34069 7361 34103 7395
rect 34103 7361 34112 7395
rect 34060 7352 34112 7361
rect 35716 7352 35768 7404
rect 37464 7395 37516 7404
rect 37464 7361 37473 7395
rect 37473 7361 37507 7395
rect 37507 7361 37516 7395
rect 37464 7352 37516 7361
rect 38568 7352 38620 7404
rect 41420 7395 41472 7404
rect 41420 7361 41429 7395
rect 41429 7361 41463 7395
rect 41463 7361 41472 7395
rect 41420 7352 41472 7361
rect 23664 7327 23716 7336
rect 23664 7293 23673 7327
rect 23673 7293 23707 7327
rect 23707 7293 23716 7327
rect 23664 7284 23716 7293
rect 23940 7284 23992 7336
rect 24400 7284 24452 7336
rect 24952 7327 25004 7336
rect 24952 7293 24961 7327
rect 24961 7293 24995 7327
rect 24995 7293 25004 7327
rect 24952 7284 25004 7293
rect 25044 7327 25096 7336
rect 25044 7293 25053 7327
rect 25053 7293 25087 7327
rect 25087 7293 25096 7327
rect 25044 7284 25096 7293
rect 23204 7216 23256 7268
rect 18788 7148 18840 7200
rect 20720 7148 20772 7200
rect 21824 7191 21876 7200
rect 21824 7157 21833 7191
rect 21833 7157 21867 7191
rect 21867 7157 21876 7191
rect 21824 7148 21876 7157
rect 22008 7148 22060 7200
rect 22192 7148 22244 7200
rect 22560 7191 22612 7200
rect 22560 7157 22569 7191
rect 22569 7157 22603 7191
rect 22603 7157 22612 7191
rect 22560 7148 22612 7157
rect 22836 7148 22888 7200
rect 24768 7216 24820 7268
rect 27160 7259 27212 7268
rect 27160 7225 27169 7259
rect 27169 7225 27203 7259
rect 27203 7225 27212 7259
rect 27160 7216 27212 7225
rect 23480 7191 23532 7200
rect 23480 7157 23489 7191
rect 23489 7157 23523 7191
rect 23523 7157 23532 7191
rect 23480 7148 23532 7157
rect 23664 7148 23716 7200
rect 25872 7148 25924 7200
rect 28540 7216 28592 7268
rect 27804 7148 27856 7200
rect 30196 7148 30248 7200
rect 32220 7216 32272 7268
rect 32404 7148 32456 7200
rect 32864 7327 32916 7336
rect 32864 7293 32873 7327
rect 32873 7293 32907 7327
rect 32907 7293 32916 7327
rect 32864 7284 32916 7293
rect 34336 7327 34388 7336
rect 34336 7293 34345 7327
rect 34345 7293 34379 7327
rect 34379 7293 34388 7327
rect 34336 7284 34388 7293
rect 34428 7284 34480 7336
rect 35532 7216 35584 7268
rect 37464 7216 37516 7268
rect 34244 7191 34296 7200
rect 34244 7157 34253 7191
rect 34253 7157 34287 7191
rect 34287 7157 34296 7191
rect 34244 7148 34296 7157
rect 35716 7148 35768 7200
rect 37280 7148 37332 7200
rect 40684 7148 40736 7200
rect 5134 7046 5186 7098
rect 5198 7046 5250 7098
rect 5262 7046 5314 7098
rect 5326 7046 5378 7098
rect 5390 7046 5442 7098
rect 35854 7046 35906 7098
rect 35918 7046 35970 7098
rect 35982 7046 36034 7098
rect 36046 7046 36098 7098
rect 36110 7046 36162 7098
rect 66574 7046 66626 7098
rect 66638 7046 66690 7098
rect 66702 7046 66754 7098
rect 66766 7046 66818 7098
rect 66830 7046 66882 7098
rect 4528 6876 4580 6928
rect 14280 6944 14332 6996
rect 15844 6944 15896 6996
rect 18788 6944 18840 6996
rect 10968 6876 11020 6928
rect 4344 6808 4396 6860
rect 14648 6876 14700 6928
rect 16488 6876 16540 6928
rect 19892 6944 19944 6996
rect 10600 6783 10652 6792
rect 10600 6749 10609 6783
rect 10609 6749 10643 6783
rect 10643 6749 10652 6783
rect 10600 6740 10652 6749
rect 10692 6740 10744 6792
rect 11612 6740 11664 6792
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 12440 6783 12492 6792
rect 12440 6749 12449 6783
rect 12449 6749 12483 6783
rect 12483 6749 12492 6783
rect 12440 6740 12492 6749
rect 11336 6672 11388 6724
rect 8392 6604 8444 6656
rect 12532 6604 12584 6656
rect 14924 6740 14976 6792
rect 16304 6808 16356 6860
rect 15476 6672 15528 6724
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 17776 6851 17828 6860
rect 17776 6817 17785 6851
rect 17785 6817 17819 6851
rect 17819 6817 17828 6851
rect 17776 6808 17828 6817
rect 18052 6808 18104 6860
rect 20536 6944 20588 6996
rect 22744 6944 22796 6996
rect 23388 6944 23440 6996
rect 21824 6876 21876 6928
rect 16488 6783 16540 6792
rect 16488 6749 16497 6783
rect 16497 6749 16531 6783
rect 16531 6749 16540 6783
rect 16488 6740 16540 6749
rect 17868 6740 17920 6792
rect 19064 6740 19116 6792
rect 19340 6740 19392 6792
rect 19616 6740 19668 6792
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 22192 6783 22244 6792
rect 22192 6749 22201 6783
rect 22201 6749 22235 6783
rect 22235 6749 22244 6783
rect 22192 6740 22244 6749
rect 14280 6647 14332 6656
rect 14280 6613 14289 6647
rect 14289 6613 14323 6647
rect 14323 6613 14332 6647
rect 14280 6604 14332 6613
rect 14372 6604 14424 6656
rect 17224 6604 17276 6656
rect 20536 6672 20588 6724
rect 22100 6672 22152 6724
rect 22376 6808 22428 6860
rect 22652 6919 22704 6928
rect 22652 6885 22661 6919
rect 22661 6885 22695 6919
rect 22695 6885 22704 6919
rect 22652 6876 22704 6885
rect 22928 6808 22980 6860
rect 23296 6808 23348 6860
rect 23480 6851 23532 6860
rect 23480 6817 23489 6851
rect 23489 6817 23523 6851
rect 23523 6817 23532 6851
rect 23480 6808 23532 6817
rect 24492 6944 24544 6996
rect 25872 6987 25924 6996
rect 25872 6953 25881 6987
rect 25881 6953 25915 6987
rect 25915 6953 25924 6987
rect 25872 6944 25924 6953
rect 27436 6944 27488 6996
rect 30564 6944 30616 6996
rect 31024 6987 31076 6996
rect 31024 6953 31033 6987
rect 31033 6953 31067 6987
rect 31067 6953 31076 6987
rect 31024 6944 31076 6953
rect 32864 6944 32916 6996
rect 35164 6944 35216 6996
rect 36360 6944 36412 6996
rect 24032 6876 24084 6928
rect 25044 6876 25096 6928
rect 24124 6808 24176 6860
rect 24492 6808 24544 6860
rect 28172 6876 28224 6928
rect 26976 6808 27028 6860
rect 28448 6808 28500 6860
rect 28632 6808 28684 6860
rect 29920 6808 29972 6860
rect 30104 6808 30156 6860
rect 22560 6740 22612 6792
rect 23572 6740 23624 6792
rect 23756 6740 23808 6792
rect 23940 6740 23992 6792
rect 18144 6604 18196 6656
rect 18512 6647 18564 6656
rect 18512 6613 18521 6647
rect 18521 6613 18555 6647
rect 18555 6613 18564 6647
rect 18512 6604 18564 6613
rect 19340 6647 19392 6656
rect 19340 6613 19349 6647
rect 19349 6613 19383 6647
rect 19383 6613 19392 6647
rect 19340 6604 19392 6613
rect 23112 6604 23164 6656
rect 23940 6604 23992 6656
rect 25504 6783 25556 6792
rect 25504 6749 25513 6783
rect 25513 6749 25547 6783
rect 25547 6749 25556 6783
rect 25504 6740 25556 6749
rect 25872 6740 25924 6792
rect 26056 6783 26108 6792
rect 26056 6749 26065 6783
rect 26065 6749 26099 6783
rect 26099 6749 26108 6783
rect 26056 6740 26108 6749
rect 28264 6740 28316 6792
rect 28540 6740 28592 6792
rect 30656 6851 30708 6860
rect 30656 6817 30665 6851
rect 30665 6817 30699 6851
rect 30699 6817 30708 6851
rect 30656 6808 30708 6817
rect 31392 6876 31444 6928
rect 31760 6876 31812 6928
rect 31668 6808 31720 6860
rect 31116 6783 31168 6792
rect 31116 6749 31125 6783
rect 31125 6749 31159 6783
rect 31159 6749 31168 6783
rect 31116 6740 31168 6749
rect 33232 6808 33284 6860
rect 34612 6876 34664 6928
rect 35256 6876 35308 6928
rect 35440 6919 35492 6928
rect 35440 6885 35449 6919
rect 35449 6885 35483 6919
rect 35483 6885 35492 6919
rect 35440 6876 35492 6885
rect 34428 6808 34480 6860
rect 34704 6808 34756 6860
rect 31852 6783 31904 6792
rect 31852 6749 31861 6783
rect 31861 6749 31895 6783
rect 31895 6749 31904 6783
rect 31852 6740 31904 6749
rect 31944 6740 31996 6792
rect 26332 6672 26384 6724
rect 30472 6672 30524 6724
rect 33140 6783 33192 6792
rect 33140 6749 33149 6783
rect 33149 6749 33183 6783
rect 33183 6749 33192 6783
rect 33140 6740 33192 6749
rect 33508 6740 33560 6792
rect 34888 6783 34940 6792
rect 34888 6749 34897 6783
rect 34897 6749 34931 6783
rect 34931 6749 34940 6783
rect 34888 6740 34940 6749
rect 38200 6808 38252 6860
rect 39396 6851 39448 6860
rect 39396 6817 39405 6851
rect 39405 6817 39439 6851
rect 39439 6817 39448 6851
rect 39396 6808 39448 6817
rect 40224 6808 40276 6860
rect 35164 6783 35216 6792
rect 35164 6749 35173 6783
rect 35173 6749 35207 6783
rect 35207 6749 35216 6783
rect 35164 6740 35216 6749
rect 35808 6783 35860 6792
rect 35808 6749 35817 6783
rect 35817 6749 35851 6783
rect 35851 6749 35860 6783
rect 35808 6740 35860 6749
rect 34244 6672 34296 6724
rect 34428 6672 34480 6724
rect 34612 6672 34664 6724
rect 28264 6604 28316 6656
rect 29000 6604 29052 6656
rect 29920 6604 29972 6656
rect 31208 6604 31260 6656
rect 31944 6604 31996 6656
rect 33508 6604 33560 6656
rect 34060 6604 34112 6656
rect 35164 6604 35216 6656
rect 35992 6672 36044 6724
rect 35900 6604 35952 6656
rect 36360 6672 36412 6724
rect 38384 6672 38436 6724
rect 44088 6740 44140 6792
rect 39580 6672 39632 6724
rect 43352 6672 43404 6724
rect 39120 6604 39172 6656
rect 40592 6647 40644 6656
rect 40592 6613 40601 6647
rect 40601 6613 40635 6647
rect 40635 6613 40644 6647
rect 40592 6604 40644 6613
rect 41420 6647 41472 6656
rect 41420 6613 41429 6647
rect 41429 6613 41463 6647
rect 41463 6613 41472 6647
rect 41420 6604 41472 6613
rect 41512 6647 41564 6656
rect 41512 6613 41521 6647
rect 41521 6613 41555 6647
rect 41555 6613 41564 6647
rect 41512 6604 41564 6613
rect 41788 6604 41840 6656
rect 5794 6502 5846 6554
rect 5858 6502 5910 6554
rect 5922 6502 5974 6554
rect 5986 6502 6038 6554
rect 6050 6502 6102 6554
rect 36514 6502 36566 6554
rect 36578 6502 36630 6554
rect 36642 6502 36694 6554
rect 36706 6502 36758 6554
rect 36770 6502 36822 6554
rect 67234 6502 67286 6554
rect 67298 6502 67350 6554
rect 67362 6502 67414 6554
rect 67426 6502 67478 6554
rect 67490 6502 67542 6554
rect 7012 6400 7064 6452
rect 10692 6400 10744 6452
rect 11612 6400 11664 6452
rect 13360 6400 13412 6452
rect 15660 6400 15712 6452
rect 16120 6400 16172 6452
rect 16672 6443 16724 6452
rect 16672 6409 16681 6443
rect 16681 6409 16715 6443
rect 16715 6409 16724 6443
rect 16672 6400 16724 6409
rect 18420 6443 18472 6452
rect 18420 6409 18429 6443
rect 18429 6409 18463 6443
rect 18463 6409 18472 6443
rect 18420 6400 18472 6409
rect 10600 6332 10652 6384
rect 13636 6332 13688 6384
rect 8116 6264 8168 6316
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 20812 6400 20864 6452
rect 21088 6400 21140 6452
rect 14556 6307 14608 6316
rect 14556 6273 14565 6307
rect 14565 6273 14599 6307
rect 14599 6273 14608 6307
rect 14556 6264 14608 6273
rect 16396 6264 16448 6316
rect 19340 6264 19392 6316
rect 19432 6264 19484 6316
rect 21640 6332 21692 6384
rect 8944 6196 8996 6248
rect 12256 6196 12308 6248
rect 15200 6196 15252 6248
rect 16580 6196 16632 6248
rect 3792 6128 3844 6180
rect 11796 6128 11848 6180
rect 11888 6128 11940 6180
rect 18144 6196 18196 6248
rect 18604 6196 18656 6248
rect 17592 6128 17644 6180
rect 19156 6239 19208 6248
rect 19156 6205 19165 6239
rect 19165 6205 19199 6239
rect 19199 6205 19208 6239
rect 19156 6196 19208 6205
rect 19800 6239 19852 6248
rect 19800 6205 19809 6239
rect 19809 6205 19843 6239
rect 19843 6205 19852 6239
rect 24400 6400 24452 6452
rect 24676 6400 24728 6452
rect 25780 6400 25832 6452
rect 26056 6400 26108 6452
rect 27252 6443 27304 6452
rect 27252 6409 27261 6443
rect 27261 6409 27295 6443
rect 27295 6409 27304 6443
rect 27252 6400 27304 6409
rect 27896 6400 27948 6452
rect 28908 6400 28960 6452
rect 30288 6443 30340 6452
rect 30288 6409 30297 6443
rect 30297 6409 30331 6443
rect 30331 6409 30340 6443
rect 30288 6400 30340 6409
rect 30380 6400 30432 6452
rect 19800 6196 19852 6205
rect 20260 6196 20312 6248
rect 22008 6239 22060 6248
rect 22008 6205 22017 6239
rect 22017 6205 22051 6239
rect 22051 6205 22060 6239
rect 22008 6196 22060 6205
rect 22652 6332 22704 6384
rect 22192 6196 22244 6248
rect 22560 6196 22612 6248
rect 22652 6196 22704 6248
rect 7932 6060 7984 6112
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 9864 6060 9916 6112
rect 12716 6103 12768 6112
rect 12716 6069 12725 6103
rect 12725 6069 12759 6103
rect 12759 6069 12768 6103
rect 12716 6060 12768 6069
rect 14648 6060 14700 6112
rect 18696 6060 18748 6112
rect 20260 6060 20312 6112
rect 23756 6264 23808 6316
rect 23296 6196 23348 6248
rect 23480 6196 23532 6248
rect 28172 6332 28224 6384
rect 24124 6264 24176 6316
rect 25412 6264 25464 6316
rect 25688 6264 25740 6316
rect 26516 6307 26568 6316
rect 26516 6273 26525 6307
rect 26525 6273 26559 6307
rect 26559 6273 26568 6307
rect 26516 6264 26568 6273
rect 24400 6239 24452 6248
rect 24400 6205 24409 6239
rect 24409 6205 24443 6239
rect 24443 6205 24452 6239
rect 24400 6196 24452 6205
rect 25780 6239 25832 6248
rect 25780 6205 25789 6239
rect 25789 6205 25823 6239
rect 25823 6205 25832 6239
rect 25780 6196 25832 6205
rect 25872 6196 25924 6248
rect 27528 6239 27580 6248
rect 27528 6205 27537 6239
rect 27537 6205 27571 6239
rect 27571 6205 27580 6239
rect 27528 6196 27580 6205
rect 28264 6307 28316 6316
rect 28264 6273 28273 6307
rect 28273 6273 28307 6307
rect 28307 6273 28316 6307
rect 28264 6264 28316 6273
rect 31484 6332 31536 6384
rect 31852 6375 31904 6384
rect 31852 6341 31861 6375
rect 31861 6341 31895 6375
rect 31895 6341 31904 6375
rect 31852 6332 31904 6341
rect 32128 6332 32180 6384
rect 30104 6264 30156 6316
rect 30472 6307 30524 6316
rect 30472 6273 30481 6307
rect 30481 6273 30515 6307
rect 30515 6273 30524 6307
rect 30472 6264 30524 6273
rect 31944 6264 31996 6316
rect 32220 6264 32272 6316
rect 34152 6400 34204 6452
rect 34244 6400 34296 6452
rect 35992 6400 36044 6452
rect 36360 6400 36412 6452
rect 38614 6400 38666 6452
rect 40592 6400 40644 6452
rect 40868 6400 40920 6452
rect 33232 6332 33284 6384
rect 33784 6332 33836 6384
rect 34612 6332 34664 6384
rect 35440 6264 35492 6316
rect 38384 6332 38436 6384
rect 38936 6332 38988 6384
rect 36176 6307 36228 6316
rect 36176 6273 36185 6307
rect 36185 6273 36219 6307
rect 36219 6273 36228 6307
rect 36176 6264 36228 6273
rect 36268 6307 36320 6316
rect 36268 6273 36277 6307
rect 36277 6273 36311 6307
rect 36311 6273 36320 6307
rect 36268 6264 36320 6273
rect 37832 6264 37884 6316
rect 38200 6307 38252 6316
rect 38200 6273 38209 6307
rect 38209 6273 38243 6307
rect 38243 6273 38252 6307
rect 38200 6264 38252 6273
rect 28816 6196 28868 6248
rect 29828 6196 29880 6248
rect 25504 6128 25556 6180
rect 30472 6128 30524 6180
rect 32220 6128 32272 6180
rect 35716 6239 35768 6248
rect 35716 6205 35725 6239
rect 35725 6205 35759 6239
rect 35759 6205 35768 6239
rect 35716 6196 35768 6205
rect 37280 6239 37332 6248
rect 37280 6205 37289 6239
rect 37289 6205 37323 6239
rect 37323 6205 37332 6239
rect 37280 6196 37332 6205
rect 21088 6060 21140 6112
rect 21272 6103 21324 6112
rect 21272 6069 21281 6103
rect 21281 6069 21315 6103
rect 21315 6069 21324 6103
rect 21272 6060 21324 6069
rect 21364 6103 21416 6112
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 21364 6060 21416 6069
rect 21456 6060 21508 6112
rect 21640 6060 21692 6112
rect 22008 6060 22060 6112
rect 22192 6060 22244 6112
rect 22284 6060 22336 6112
rect 22560 6103 22612 6112
rect 22560 6069 22569 6103
rect 22569 6069 22603 6103
rect 22603 6069 22612 6103
rect 22560 6060 22612 6069
rect 25044 6060 25096 6112
rect 25320 6060 25372 6112
rect 27436 6060 27488 6112
rect 30840 6060 30892 6112
rect 33876 6060 33928 6112
rect 35440 6060 35492 6112
rect 36912 6060 36964 6112
rect 37556 6128 37608 6180
rect 38568 6196 38620 6248
rect 40500 6332 40552 6384
rect 42524 6332 42576 6384
rect 41420 6264 41472 6316
rect 40224 6239 40276 6248
rect 40224 6205 40233 6239
rect 40233 6205 40267 6239
rect 40267 6205 40276 6239
rect 40224 6196 40276 6205
rect 41328 6196 41380 6248
rect 43076 6264 43128 6316
rect 41972 6239 42024 6248
rect 41972 6205 41981 6239
rect 41981 6205 42015 6239
rect 42015 6205 42024 6239
rect 41972 6196 42024 6205
rect 39856 6060 39908 6112
rect 41144 6103 41196 6112
rect 41144 6069 41153 6103
rect 41153 6069 41187 6103
rect 41187 6069 41196 6103
rect 41144 6060 41196 6069
rect 42616 6103 42668 6112
rect 42616 6069 42625 6103
rect 42625 6069 42659 6103
rect 42659 6069 42668 6103
rect 42616 6060 42668 6069
rect 42800 6060 42852 6112
rect 5134 5958 5186 6010
rect 5198 5958 5250 6010
rect 5262 5958 5314 6010
rect 5326 5958 5378 6010
rect 5390 5958 5442 6010
rect 35854 5958 35906 6010
rect 35918 5958 35970 6010
rect 35982 5958 36034 6010
rect 36046 5958 36098 6010
rect 36110 5958 36162 6010
rect 66574 5958 66626 6010
rect 66638 5958 66690 6010
rect 66702 5958 66754 6010
rect 66766 5958 66818 6010
rect 66830 5958 66882 6010
rect 3608 5856 3660 5908
rect 9772 5856 9824 5908
rect 10140 5899 10192 5908
rect 10140 5865 10149 5899
rect 10149 5865 10183 5899
rect 10183 5865 10192 5899
rect 10140 5856 10192 5865
rect 11152 5899 11204 5908
rect 11152 5865 11161 5899
rect 11161 5865 11195 5899
rect 11195 5865 11204 5899
rect 11152 5856 11204 5865
rect 7564 5788 7616 5840
rect 9864 5788 9916 5840
rect 7840 5720 7892 5772
rect 12440 5856 12492 5908
rect 14464 5856 14516 5908
rect 15108 5856 15160 5908
rect 15568 5788 15620 5840
rect 8300 5652 8352 5704
rect 8024 5584 8076 5636
rect 10324 5652 10376 5704
rect 10692 5652 10744 5704
rect 11336 5652 11388 5704
rect 11428 5695 11480 5704
rect 11428 5661 11437 5695
rect 11437 5661 11471 5695
rect 11471 5661 11480 5695
rect 11428 5652 11480 5661
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 16028 5720 16080 5772
rect 16304 5763 16356 5772
rect 16304 5729 16313 5763
rect 16313 5729 16347 5763
rect 16347 5729 16356 5763
rect 16304 5720 16356 5729
rect 12440 5584 12492 5636
rect 4712 5516 4764 5568
rect 9772 5516 9824 5568
rect 12072 5516 12124 5568
rect 13820 5652 13872 5704
rect 14096 5652 14148 5704
rect 14740 5584 14792 5636
rect 13268 5516 13320 5568
rect 15292 5627 15344 5636
rect 15292 5593 15301 5627
rect 15301 5593 15335 5627
rect 15335 5593 15344 5627
rect 15292 5584 15344 5593
rect 18420 5856 18472 5908
rect 18604 5856 18656 5908
rect 19432 5856 19484 5908
rect 19524 5856 19576 5908
rect 21180 5856 21232 5908
rect 16488 5788 16540 5840
rect 22928 5856 22980 5908
rect 21732 5788 21784 5840
rect 24768 5856 24820 5908
rect 27528 5856 27580 5908
rect 19156 5720 19208 5772
rect 19340 5763 19392 5772
rect 19340 5729 19349 5763
rect 19349 5729 19383 5763
rect 19383 5729 19392 5763
rect 19340 5720 19392 5729
rect 17684 5652 17736 5704
rect 16580 5584 16632 5636
rect 18696 5652 18748 5704
rect 20444 5720 20496 5772
rect 21824 5720 21876 5772
rect 22468 5720 22520 5772
rect 23020 5720 23072 5772
rect 23480 5788 23532 5840
rect 23756 5788 23808 5840
rect 23848 5788 23900 5840
rect 24308 5788 24360 5840
rect 26976 5788 27028 5840
rect 23572 5720 23624 5772
rect 33784 5856 33836 5908
rect 35256 5856 35308 5908
rect 35716 5856 35768 5908
rect 35992 5856 36044 5908
rect 36452 5856 36504 5908
rect 37556 5856 37608 5908
rect 38660 5856 38712 5908
rect 39580 5856 39632 5908
rect 41604 5856 41656 5908
rect 20720 5652 20772 5704
rect 20904 5695 20956 5704
rect 20904 5661 20913 5695
rect 20913 5661 20947 5695
rect 20947 5661 20956 5695
rect 20904 5652 20956 5661
rect 22652 5652 22704 5704
rect 15200 5516 15252 5568
rect 16304 5516 16356 5568
rect 16396 5559 16448 5568
rect 16396 5525 16405 5559
rect 16405 5525 16439 5559
rect 16439 5525 16448 5559
rect 16396 5516 16448 5525
rect 17868 5516 17920 5568
rect 17960 5516 18012 5568
rect 21272 5584 21324 5636
rect 23756 5652 23808 5704
rect 23848 5695 23900 5704
rect 23848 5661 23857 5695
rect 23857 5661 23891 5695
rect 23891 5661 23900 5695
rect 23848 5652 23900 5661
rect 24492 5695 24544 5704
rect 24492 5661 24501 5695
rect 24501 5661 24535 5695
rect 24535 5661 24544 5695
rect 24492 5652 24544 5661
rect 25504 5695 25556 5704
rect 25504 5661 25513 5695
rect 25513 5661 25547 5695
rect 25547 5661 25556 5695
rect 25504 5652 25556 5661
rect 25964 5652 26016 5704
rect 30104 5652 30156 5704
rect 30840 5720 30892 5772
rect 19432 5516 19484 5568
rect 20352 5516 20404 5568
rect 21364 5516 21416 5568
rect 23480 5584 23532 5636
rect 26976 5584 27028 5636
rect 22192 5559 22244 5568
rect 22192 5525 22201 5559
rect 22201 5525 22235 5559
rect 22235 5525 22244 5559
rect 22192 5516 22244 5525
rect 22284 5516 22336 5568
rect 22468 5516 22520 5568
rect 22560 5516 22612 5568
rect 25412 5516 25464 5568
rect 26056 5559 26108 5568
rect 26056 5525 26065 5559
rect 26065 5525 26099 5559
rect 26099 5525 26108 5559
rect 26056 5516 26108 5525
rect 27252 5516 27304 5568
rect 27896 5516 27948 5568
rect 29184 5516 29236 5568
rect 30196 5516 30248 5568
rect 30656 5516 30708 5568
rect 31208 5720 31260 5772
rect 33508 5788 33560 5840
rect 34152 5788 34204 5840
rect 31484 5695 31536 5704
rect 31484 5661 31493 5695
rect 31493 5661 31527 5695
rect 31527 5661 31536 5695
rect 31484 5652 31536 5661
rect 31668 5652 31720 5704
rect 31944 5695 31996 5704
rect 31944 5661 31953 5695
rect 31953 5661 31987 5695
rect 31987 5661 31996 5695
rect 31944 5652 31996 5661
rect 32220 5584 32272 5636
rect 33692 5652 33744 5704
rect 34336 5720 34388 5772
rect 36268 5788 36320 5840
rect 35532 5652 35584 5704
rect 34336 5627 34388 5636
rect 34336 5593 34345 5627
rect 34345 5593 34379 5627
rect 34379 5593 34388 5627
rect 34336 5584 34388 5593
rect 33692 5516 33744 5568
rect 33968 5516 34020 5568
rect 34704 5516 34756 5568
rect 34980 5516 35032 5568
rect 35992 5695 36044 5704
rect 35992 5661 36001 5695
rect 36001 5661 36035 5695
rect 36035 5661 36044 5695
rect 35992 5652 36044 5661
rect 36176 5695 36228 5704
rect 36176 5661 36185 5695
rect 36185 5661 36219 5695
rect 36219 5661 36228 5695
rect 36176 5652 36228 5661
rect 37280 5720 37332 5772
rect 39120 5763 39172 5772
rect 39120 5729 39129 5763
rect 39129 5729 39163 5763
rect 39163 5729 39172 5763
rect 39120 5720 39172 5729
rect 37832 5652 37884 5704
rect 38568 5652 38620 5704
rect 39396 5652 39448 5704
rect 41420 5788 41472 5840
rect 41144 5720 41196 5772
rect 42616 5720 42668 5772
rect 41788 5652 41840 5704
rect 42064 5695 42116 5704
rect 42064 5661 42073 5695
rect 42073 5661 42107 5695
rect 42107 5661 42116 5695
rect 42064 5652 42116 5661
rect 42984 5652 43036 5704
rect 43168 5652 43220 5704
rect 45928 5652 45980 5704
rect 48780 5652 48832 5704
rect 36268 5584 36320 5636
rect 40868 5584 40920 5636
rect 49792 5584 49844 5636
rect 37832 5516 37884 5568
rect 38200 5559 38252 5568
rect 38200 5525 38209 5559
rect 38209 5525 38243 5559
rect 38243 5525 38252 5559
rect 38200 5516 38252 5525
rect 39028 5516 39080 5568
rect 40500 5516 40552 5568
rect 41696 5516 41748 5568
rect 44272 5559 44324 5568
rect 44272 5525 44281 5559
rect 44281 5525 44315 5559
rect 44315 5525 44324 5559
rect 44272 5516 44324 5525
rect 46940 5516 46992 5568
rect 5794 5414 5846 5466
rect 5858 5414 5910 5466
rect 5922 5414 5974 5466
rect 5986 5414 6038 5466
rect 6050 5414 6102 5466
rect 36514 5414 36566 5466
rect 36578 5414 36630 5466
rect 36642 5414 36694 5466
rect 36706 5414 36758 5466
rect 36770 5414 36822 5466
rect 67234 5414 67286 5466
rect 67298 5414 67350 5466
rect 67362 5414 67414 5466
rect 67426 5414 67478 5466
rect 67490 5414 67542 5466
rect 10692 5312 10744 5364
rect 10784 5355 10836 5364
rect 10784 5321 10793 5355
rect 10793 5321 10827 5355
rect 10827 5321 10836 5355
rect 10784 5312 10836 5321
rect 11888 5312 11940 5364
rect 15016 5312 15068 5364
rect 15200 5355 15252 5364
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 15936 5355 15988 5364
rect 15936 5321 15945 5355
rect 15945 5321 15979 5355
rect 15979 5321 15988 5355
rect 15936 5312 15988 5321
rect 18144 5355 18196 5364
rect 18144 5321 18153 5355
rect 18153 5321 18187 5355
rect 18187 5321 18196 5355
rect 18144 5312 18196 5321
rect 18972 5312 19024 5364
rect 19156 5312 19208 5364
rect 12532 5244 12584 5296
rect 12992 5287 13044 5296
rect 12992 5253 13001 5287
rect 13001 5253 13035 5287
rect 13035 5253 13044 5287
rect 12992 5244 13044 5253
rect 16212 5244 16264 5296
rect 18512 5244 18564 5296
rect 20536 5312 20588 5364
rect 21548 5312 21600 5364
rect 9864 5176 9916 5228
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 10416 5176 10468 5228
rect 11612 5219 11664 5228
rect 11612 5185 11621 5219
rect 11621 5185 11655 5219
rect 11655 5185 11664 5219
rect 11612 5176 11664 5185
rect 12348 5176 12400 5228
rect 15016 5176 15068 5228
rect 16856 5176 16908 5228
rect 17592 5219 17644 5228
rect 17592 5185 17601 5219
rect 17601 5185 17635 5219
rect 17635 5185 17644 5219
rect 17592 5176 17644 5185
rect 17684 5176 17736 5228
rect 18144 5176 18196 5228
rect 20352 5176 20404 5228
rect 13176 5151 13228 5160
rect 13176 5117 13185 5151
rect 13185 5117 13219 5151
rect 13219 5117 13228 5151
rect 13176 5108 13228 5117
rect 13820 5151 13872 5160
rect 13820 5117 13829 5151
rect 13829 5117 13863 5151
rect 13863 5117 13872 5151
rect 13820 5108 13872 5117
rect 13912 5108 13964 5160
rect 15292 5151 15344 5160
rect 15292 5117 15301 5151
rect 15301 5117 15335 5151
rect 15335 5117 15344 5151
rect 15292 5108 15344 5117
rect 15752 5108 15804 5160
rect 16304 5108 16356 5160
rect 16764 5151 16816 5160
rect 16764 5117 16773 5151
rect 16773 5117 16807 5151
rect 16807 5117 16816 5151
rect 16764 5108 16816 5117
rect 18236 5151 18288 5160
rect 18236 5117 18245 5151
rect 18245 5117 18279 5151
rect 18279 5117 18288 5151
rect 18236 5108 18288 5117
rect 18512 5108 18564 5160
rect 20996 5244 21048 5296
rect 21732 5355 21784 5364
rect 21732 5321 21741 5355
rect 21741 5321 21775 5355
rect 21775 5321 21784 5355
rect 21732 5312 21784 5321
rect 21824 5312 21876 5364
rect 23664 5312 23716 5364
rect 24032 5355 24084 5364
rect 24032 5321 24041 5355
rect 24041 5321 24075 5355
rect 24075 5321 24084 5355
rect 24032 5312 24084 5321
rect 24860 5312 24912 5364
rect 28816 5312 28868 5364
rect 20812 5176 20864 5228
rect 21456 5176 21508 5228
rect 22284 5244 22336 5296
rect 23572 5244 23624 5296
rect 23848 5244 23900 5296
rect 28172 5287 28224 5296
rect 28172 5253 28181 5287
rect 28181 5253 28215 5287
rect 28215 5253 28224 5287
rect 28172 5244 28224 5253
rect 9956 4972 10008 5024
rect 10416 5040 10468 5092
rect 12440 4972 12492 5024
rect 14556 4972 14608 5024
rect 17592 4972 17644 5024
rect 18512 4972 18564 5024
rect 20444 5040 20496 5092
rect 21732 5108 21784 5160
rect 21824 5040 21876 5092
rect 23112 5108 23164 5160
rect 25412 5108 25464 5160
rect 25688 5219 25740 5228
rect 25688 5185 25697 5219
rect 25697 5185 25731 5219
rect 25731 5185 25740 5219
rect 25688 5176 25740 5185
rect 28724 5176 28776 5228
rect 31852 5312 31904 5364
rect 26884 5108 26936 5160
rect 26976 5108 27028 5160
rect 23020 4972 23072 5024
rect 24124 5040 24176 5092
rect 24308 5040 24360 5092
rect 29000 5108 29052 5160
rect 27528 5040 27580 5092
rect 29276 5176 29328 5228
rect 30380 5176 30432 5228
rect 32404 5312 32456 5364
rect 33140 5312 33192 5364
rect 33692 5312 33744 5364
rect 33508 5244 33560 5296
rect 32312 5176 32364 5228
rect 29552 5151 29604 5160
rect 29552 5117 29561 5151
rect 29561 5117 29595 5151
rect 29595 5117 29604 5151
rect 29552 5108 29604 5117
rect 29368 5040 29420 5092
rect 32956 5108 33008 5160
rect 33876 5151 33928 5160
rect 33876 5117 33885 5151
rect 33885 5117 33919 5151
rect 33919 5117 33928 5151
rect 33876 5108 33928 5117
rect 34060 5219 34112 5228
rect 34060 5185 34069 5219
rect 34069 5185 34103 5219
rect 34103 5185 34112 5219
rect 34060 5176 34112 5185
rect 36820 5312 36872 5364
rect 39764 5312 39816 5364
rect 39856 5312 39908 5364
rect 41604 5312 41656 5364
rect 42064 5312 42116 5364
rect 42524 5312 42576 5364
rect 34612 5176 34664 5228
rect 36544 5244 36596 5296
rect 37740 5244 37792 5296
rect 40132 5244 40184 5296
rect 42156 5244 42208 5296
rect 35164 5176 35216 5228
rect 36084 5176 36136 5228
rect 37556 5176 37608 5228
rect 35440 5108 35492 5160
rect 36452 5108 36504 5160
rect 40500 5219 40552 5228
rect 40500 5185 40509 5219
rect 40509 5185 40543 5219
rect 40543 5185 40552 5219
rect 40500 5176 40552 5185
rect 43076 5176 43128 5228
rect 43536 5176 43588 5228
rect 44272 5176 44324 5228
rect 46940 5219 46992 5228
rect 46940 5185 46949 5219
rect 46949 5185 46983 5219
rect 46983 5185 46992 5219
rect 46940 5176 46992 5185
rect 23756 4972 23808 5024
rect 25412 5015 25464 5024
rect 25412 4981 25421 5015
rect 25421 4981 25455 5015
rect 25455 4981 25464 5015
rect 25412 4972 25464 4981
rect 30196 4972 30248 5024
rect 30564 4972 30616 5024
rect 34244 5040 34296 5092
rect 34888 5040 34940 5092
rect 36544 5040 36596 5092
rect 37740 5040 37792 5092
rect 38660 5108 38712 5160
rect 39028 5151 39080 5160
rect 39028 5117 39037 5151
rect 39037 5117 39071 5151
rect 39071 5117 39080 5151
rect 39028 5108 39080 5117
rect 41604 5108 41656 5160
rect 42064 5108 42116 5160
rect 44640 5108 44692 5160
rect 44732 5151 44784 5160
rect 44732 5117 44741 5151
rect 44741 5117 44775 5151
rect 44775 5117 44784 5151
rect 44732 5108 44784 5117
rect 76932 5108 76984 5160
rect 31852 4972 31904 5024
rect 33232 4972 33284 5024
rect 35164 4972 35216 5024
rect 37924 4972 37976 5024
rect 42892 5040 42944 5092
rect 39948 4972 40000 5024
rect 43076 5015 43128 5024
rect 43076 4981 43085 5015
rect 43085 4981 43119 5015
rect 43119 4981 43128 5015
rect 43076 4972 43128 4981
rect 45836 4972 45888 5024
rect 46296 5015 46348 5024
rect 46296 4981 46305 5015
rect 46305 4981 46339 5015
rect 46339 4981 46348 5015
rect 46296 4972 46348 4981
rect 76656 4972 76708 5024
rect 5134 4870 5186 4922
rect 5198 4870 5250 4922
rect 5262 4870 5314 4922
rect 5326 4870 5378 4922
rect 5390 4870 5442 4922
rect 35854 4870 35906 4922
rect 35918 4870 35970 4922
rect 35982 4870 36034 4922
rect 36046 4870 36098 4922
rect 36110 4870 36162 4922
rect 66574 4870 66626 4922
rect 66638 4870 66690 4922
rect 66702 4870 66754 4922
rect 66766 4870 66818 4922
rect 66830 4870 66882 4922
rect 8944 4811 8996 4820
rect 8944 4777 8953 4811
rect 8953 4777 8987 4811
rect 8987 4777 8996 4811
rect 8944 4768 8996 4777
rect 11060 4768 11112 4820
rect 11980 4768 12032 4820
rect 12624 4811 12676 4820
rect 12624 4777 12633 4811
rect 12633 4777 12667 4811
rect 12667 4777 12676 4811
rect 12624 4768 12676 4777
rect 13544 4768 13596 4820
rect 16580 4768 16632 4820
rect 17040 4811 17092 4820
rect 17040 4777 17049 4811
rect 17049 4777 17083 4811
rect 17083 4777 17092 4811
rect 17040 4768 17092 4777
rect 9772 4632 9824 4684
rect 9956 4632 10008 4684
rect 11244 4632 11296 4684
rect 11612 4632 11664 4684
rect 7380 4607 7432 4616
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 10692 4564 10744 4616
rect 9956 4496 10008 4548
rect 10048 4539 10100 4548
rect 10048 4505 10057 4539
rect 10057 4505 10091 4539
rect 10091 4505 10100 4539
rect 10048 4496 10100 4505
rect 11060 4496 11112 4548
rect 12440 4700 12492 4752
rect 13176 4700 13228 4752
rect 14188 4700 14240 4752
rect 12164 4632 12216 4684
rect 14372 4632 14424 4684
rect 14464 4632 14516 4684
rect 17684 4700 17736 4752
rect 18512 4743 18564 4752
rect 18512 4709 18521 4743
rect 18521 4709 18555 4743
rect 18555 4709 18564 4743
rect 18512 4700 18564 4709
rect 19248 4743 19300 4752
rect 19248 4709 19257 4743
rect 19257 4709 19291 4743
rect 19291 4709 19300 4743
rect 19248 4700 19300 4709
rect 19616 4700 19668 4752
rect 20444 4700 20496 4752
rect 22100 4768 22152 4820
rect 22744 4768 22796 4820
rect 22928 4811 22980 4820
rect 22928 4777 22937 4811
rect 22937 4777 22971 4811
rect 22971 4777 22980 4811
rect 22928 4768 22980 4777
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 13544 4564 13596 4616
rect 15108 4607 15160 4616
rect 15108 4573 15117 4607
rect 15117 4573 15151 4607
rect 15151 4573 15160 4607
rect 15108 4564 15160 4573
rect 15660 4564 15712 4616
rect 15844 4564 15896 4616
rect 18604 4564 18656 4616
rect 18696 4607 18748 4616
rect 18696 4573 18705 4607
rect 18705 4573 18739 4607
rect 18739 4573 18748 4607
rect 18696 4564 18748 4573
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 19616 4564 19668 4616
rect 19984 4564 20036 4616
rect 21180 4564 21232 4616
rect 23020 4632 23072 4684
rect 22100 4564 22152 4616
rect 22284 4607 22336 4616
rect 22284 4573 22293 4607
rect 22293 4573 22327 4607
rect 22327 4573 22336 4607
rect 22284 4564 22336 4573
rect 14280 4496 14332 4548
rect 6828 4471 6880 4480
rect 6828 4437 6837 4471
rect 6837 4437 6871 4471
rect 6871 4437 6880 4471
rect 6828 4428 6880 4437
rect 9404 4428 9456 4480
rect 11152 4471 11204 4480
rect 11152 4437 11161 4471
rect 11161 4437 11195 4471
rect 11195 4437 11204 4471
rect 11152 4428 11204 4437
rect 11428 4428 11480 4480
rect 12808 4428 12860 4480
rect 20260 4496 20312 4548
rect 24124 4632 24176 4684
rect 24400 4700 24452 4752
rect 25412 4700 25464 4752
rect 26608 4700 26660 4752
rect 29828 4768 29880 4820
rect 31300 4768 31352 4820
rect 31576 4768 31628 4820
rect 32772 4768 32824 4820
rect 33784 4768 33836 4820
rect 36084 4768 36136 4820
rect 36268 4768 36320 4820
rect 36452 4768 36504 4820
rect 37464 4768 37516 4820
rect 37924 4768 37976 4820
rect 47032 4768 47084 4820
rect 76932 4811 76984 4820
rect 76932 4777 76941 4811
rect 76941 4777 76975 4811
rect 76975 4777 76984 4811
rect 76932 4768 76984 4777
rect 28264 4632 28316 4684
rect 28356 4675 28408 4684
rect 28356 4641 28365 4675
rect 28365 4641 28399 4675
rect 28399 4641 28408 4675
rect 28356 4632 28408 4641
rect 24768 4564 24820 4616
rect 25228 4564 25280 4616
rect 26516 4607 26568 4616
rect 26516 4573 26525 4607
rect 26525 4573 26559 4607
rect 26559 4573 26568 4607
rect 26516 4564 26568 4573
rect 27528 4564 27580 4616
rect 27620 4564 27672 4616
rect 28908 4675 28960 4684
rect 28908 4641 28917 4675
rect 28917 4641 28951 4675
rect 28951 4641 28960 4675
rect 28908 4632 28960 4641
rect 29092 4632 29144 4684
rect 29276 4632 29328 4684
rect 30472 4564 30524 4616
rect 30840 4632 30892 4684
rect 16120 4428 16172 4480
rect 16304 4471 16356 4480
rect 16304 4437 16313 4471
rect 16313 4437 16347 4471
rect 16347 4437 16356 4471
rect 16304 4428 16356 4437
rect 16672 4428 16724 4480
rect 19524 4428 19576 4480
rect 19984 4471 20036 4480
rect 19984 4437 19993 4471
rect 19993 4437 20027 4471
rect 20027 4437 20036 4471
rect 19984 4428 20036 4437
rect 22100 4471 22152 4480
rect 22100 4437 22109 4471
rect 22109 4437 22143 4471
rect 22143 4437 22152 4471
rect 22100 4428 22152 4437
rect 23664 4428 23716 4480
rect 25412 4428 25464 4480
rect 28816 4496 28868 4548
rect 27068 4428 27120 4480
rect 28080 4428 28132 4480
rect 28448 4428 28500 4480
rect 30288 4471 30340 4480
rect 30288 4437 30297 4471
rect 30297 4437 30331 4471
rect 30331 4437 30340 4471
rect 30288 4428 30340 4437
rect 31208 4564 31260 4616
rect 31668 4700 31720 4752
rect 31852 4675 31904 4684
rect 31852 4641 31861 4675
rect 31861 4641 31895 4675
rect 31895 4641 31904 4675
rect 31852 4632 31904 4641
rect 32220 4632 32272 4684
rect 32956 4675 33008 4684
rect 32956 4641 32965 4675
rect 32965 4641 32999 4675
rect 32999 4641 33008 4675
rect 32956 4632 33008 4641
rect 34980 4700 35032 4752
rect 41328 4700 41380 4752
rect 34888 4675 34940 4684
rect 34888 4641 34897 4675
rect 34897 4641 34931 4675
rect 34931 4641 34940 4675
rect 34888 4632 34940 4641
rect 36912 4632 36964 4684
rect 31576 4496 31628 4548
rect 34612 4564 34664 4616
rect 36084 4496 36136 4548
rect 37740 4607 37792 4616
rect 37740 4573 37749 4607
rect 37749 4573 37783 4607
rect 37783 4573 37792 4607
rect 37740 4564 37792 4573
rect 37832 4607 37884 4616
rect 37832 4573 37841 4607
rect 37841 4573 37875 4607
rect 37875 4573 37884 4607
rect 37832 4564 37884 4573
rect 39856 4675 39908 4684
rect 39856 4641 39865 4675
rect 39865 4641 39899 4675
rect 39899 4641 39908 4675
rect 39856 4632 39908 4641
rect 39948 4675 40000 4684
rect 39948 4641 39957 4675
rect 39957 4641 39991 4675
rect 39991 4641 40000 4675
rect 39948 4632 40000 4641
rect 43076 4700 43128 4752
rect 43352 4632 43404 4684
rect 44088 4632 44140 4684
rect 45192 4632 45244 4684
rect 47216 4632 47268 4684
rect 41788 4607 41840 4616
rect 41788 4573 41797 4607
rect 41797 4573 41831 4607
rect 41831 4573 41840 4607
rect 41788 4564 41840 4573
rect 42616 4564 42668 4616
rect 38384 4496 38436 4548
rect 32128 4428 32180 4480
rect 33784 4428 33836 4480
rect 35440 4471 35492 4480
rect 35440 4437 35449 4471
rect 35449 4437 35483 4471
rect 35483 4437 35492 4471
rect 35440 4428 35492 4437
rect 37556 4428 37608 4480
rect 39488 4496 39540 4548
rect 40040 4496 40092 4548
rect 40132 4496 40184 4548
rect 40960 4496 41012 4548
rect 43076 4564 43128 4616
rect 44180 4607 44232 4616
rect 44180 4573 44189 4607
rect 44189 4573 44223 4607
rect 44223 4573 44232 4607
rect 44180 4564 44232 4573
rect 45468 4496 45520 4548
rect 45652 4496 45704 4548
rect 48044 4607 48096 4616
rect 48044 4573 48053 4607
rect 48053 4573 48087 4607
rect 48087 4573 48096 4607
rect 48044 4564 48096 4573
rect 48872 4607 48924 4616
rect 48872 4573 48881 4607
rect 48881 4573 48915 4607
rect 48915 4573 48924 4607
rect 48872 4564 48924 4573
rect 77576 4607 77628 4616
rect 77576 4573 77585 4607
rect 77585 4573 77619 4607
rect 77619 4573 77628 4607
rect 77576 4564 77628 4573
rect 49976 4496 50028 4548
rect 42248 4428 42300 4480
rect 43260 4428 43312 4480
rect 43352 4471 43404 4480
rect 43352 4437 43361 4471
rect 43361 4437 43395 4471
rect 43395 4437 43404 4471
rect 43352 4428 43404 4437
rect 45560 4428 45612 4480
rect 48320 4428 48372 4480
rect 50528 4428 50580 4480
rect 5794 4326 5846 4378
rect 5858 4326 5910 4378
rect 5922 4326 5974 4378
rect 5986 4326 6038 4378
rect 6050 4326 6102 4378
rect 36514 4326 36566 4378
rect 36578 4326 36630 4378
rect 36642 4326 36694 4378
rect 36706 4326 36758 4378
rect 36770 4326 36822 4378
rect 67234 4326 67286 4378
rect 67298 4326 67350 4378
rect 67362 4326 67414 4378
rect 67426 4326 67478 4378
rect 67490 4326 67542 4378
rect 7380 4224 7432 4276
rect 9772 4224 9824 4276
rect 9956 4224 10008 4276
rect 11244 4224 11296 4276
rect 13452 4224 13504 4276
rect 14464 4224 14516 4276
rect 15108 4224 15160 4276
rect 16672 4224 16724 4276
rect 19892 4267 19944 4276
rect 19892 4233 19901 4267
rect 19901 4233 19935 4267
rect 19935 4233 19944 4267
rect 19892 4224 19944 4233
rect 26424 4224 26476 4276
rect 26700 4224 26752 4276
rect 28816 4224 28868 4276
rect 30656 4224 30708 4276
rect 31116 4224 31168 4276
rect 32220 4224 32272 4276
rect 32496 4224 32548 4276
rect 32956 4224 33008 4276
rect 34060 4224 34112 4276
rect 40960 4224 41012 4276
rect 41328 4224 41380 4276
rect 44180 4224 44232 4276
rect 6368 4156 6420 4208
rect 6920 4156 6972 4208
rect 10232 4156 10284 4208
rect 6000 4088 6052 4140
rect 8576 4020 8628 4072
rect 10324 4088 10376 4140
rect 16764 4156 16816 4208
rect 11152 4088 11204 4140
rect 12624 4088 12676 4140
rect 13728 4088 13780 4140
rect 14648 4088 14700 4140
rect 4896 3952 4948 4004
rect 8116 3952 8168 4004
rect 10140 4020 10192 4072
rect 10416 4020 10468 4072
rect 10876 4063 10928 4072
rect 10876 4029 10885 4063
rect 10885 4029 10919 4063
rect 10919 4029 10928 4063
rect 10876 4020 10928 4029
rect 11612 4020 11664 4072
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 11888 4020 11940 4072
rect 9956 3952 10008 4004
rect 11980 3952 12032 4004
rect 5540 3884 5592 3936
rect 13820 3952 13872 4004
rect 14648 3952 14700 4004
rect 14832 4131 14884 4140
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 15016 4131 15068 4140
rect 15016 4097 15025 4131
rect 15025 4097 15059 4131
rect 15059 4097 15068 4131
rect 15016 4088 15068 4097
rect 15108 4020 15160 4072
rect 16396 4088 16448 4140
rect 16580 4088 16632 4140
rect 17224 4131 17276 4140
rect 17224 4097 17233 4131
rect 17233 4097 17267 4131
rect 17267 4097 17276 4131
rect 17224 4088 17276 4097
rect 17592 4156 17644 4208
rect 19340 4156 19392 4208
rect 19524 4156 19576 4208
rect 18236 4020 18288 4072
rect 18144 3995 18196 4004
rect 18144 3961 18153 3995
rect 18153 3961 18187 3995
rect 18187 3961 18196 3995
rect 18144 3952 18196 3961
rect 19156 4088 19208 4140
rect 20444 4199 20496 4208
rect 20444 4165 20453 4199
rect 20453 4165 20487 4199
rect 20487 4165 20496 4199
rect 20444 4156 20496 4165
rect 20628 4199 20680 4208
rect 20628 4165 20653 4199
rect 20653 4165 20680 4199
rect 20628 4156 20680 4165
rect 21088 4156 21140 4208
rect 18788 4020 18840 4072
rect 20260 4020 20312 4072
rect 24124 4156 24176 4208
rect 25872 4156 25924 4208
rect 22836 4131 22888 4140
rect 22836 4097 22845 4131
rect 22845 4097 22879 4131
rect 22879 4097 22888 4131
rect 22836 4088 22888 4097
rect 23572 4088 23624 4140
rect 24032 4088 24084 4140
rect 26056 4088 26108 4140
rect 26424 4131 26476 4140
rect 26424 4097 26433 4131
rect 26433 4097 26467 4131
rect 26467 4097 26476 4131
rect 26424 4088 26476 4097
rect 27988 4156 28040 4208
rect 28264 4156 28316 4208
rect 21824 4020 21876 4072
rect 22652 4020 22704 4072
rect 23664 4063 23716 4072
rect 23664 4029 23673 4063
rect 23673 4029 23707 4063
rect 23707 4029 23716 4063
rect 23664 4020 23716 4029
rect 25964 4020 26016 4072
rect 27068 4020 27120 4072
rect 28448 4131 28500 4140
rect 28448 4097 28457 4131
rect 28457 4097 28491 4131
rect 28491 4097 28500 4131
rect 28448 4088 28500 4097
rect 26700 3995 26752 4004
rect 26700 3961 26709 3995
rect 26709 3961 26743 3995
rect 26743 3961 26752 3995
rect 26700 3952 26752 3961
rect 29092 4063 29144 4072
rect 29092 4029 29101 4063
rect 29101 4029 29135 4063
rect 29135 4029 29144 4063
rect 29092 4020 29144 4029
rect 29644 4020 29696 4072
rect 31116 4088 31168 4140
rect 32496 4020 32548 4072
rect 13268 3884 13320 3936
rect 14464 3884 14516 3936
rect 19432 3884 19484 3936
rect 19524 3927 19576 3936
rect 19524 3893 19533 3927
rect 19533 3893 19567 3927
rect 19567 3893 19576 3927
rect 19524 3884 19576 3893
rect 20076 3884 20128 3936
rect 20720 3884 20772 3936
rect 20904 3927 20956 3936
rect 20904 3893 20913 3927
rect 20913 3893 20947 3927
rect 20947 3893 20956 3927
rect 20904 3884 20956 3893
rect 20996 3884 21048 3936
rect 26424 3884 26476 3936
rect 27436 3927 27488 3936
rect 27436 3893 27445 3927
rect 27445 3893 27479 3927
rect 27479 3893 27488 3927
rect 27436 3884 27488 3893
rect 29184 3952 29236 4004
rect 29460 3952 29512 4004
rect 31576 3952 31628 4004
rect 31668 3952 31720 4004
rect 32680 4131 32732 4140
rect 32680 4097 32689 4131
rect 32689 4097 32723 4131
rect 32723 4097 32732 4131
rect 32680 4088 32732 4097
rect 33048 4131 33100 4140
rect 33048 4097 33057 4131
rect 33057 4097 33091 4131
rect 33091 4097 33100 4131
rect 33048 4088 33100 4097
rect 33232 4131 33284 4140
rect 33232 4097 33241 4131
rect 33241 4097 33275 4131
rect 33275 4097 33284 4131
rect 33232 4088 33284 4097
rect 34612 4156 34664 4208
rect 39948 4156 40000 4208
rect 40040 4156 40092 4208
rect 41604 4156 41656 4208
rect 42248 4156 42300 4208
rect 42616 4156 42668 4208
rect 45376 4156 45428 4208
rect 52644 4199 52696 4208
rect 52644 4165 52653 4199
rect 52653 4165 52687 4199
rect 52687 4165 52696 4199
rect 52644 4156 52696 4165
rect 33968 4063 34020 4072
rect 33968 4029 33977 4063
rect 33977 4029 34011 4063
rect 34011 4029 34020 4063
rect 33968 4020 34020 4029
rect 34520 4020 34572 4072
rect 34888 4020 34940 4072
rect 35164 4020 35216 4072
rect 35256 3952 35308 4004
rect 32772 3884 32824 3936
rect 35532 3884 35584 3936
rect 36084 4131 36136 4140
rect 36084 4097 36093 4131
rect 36093 4097 36127 4131
rect 36127 4097 36136 4131
rect 36084 4088 36136 4097
rect 36176 4131 36228 4140
rect 36176 4097 36185 4131
rect 36185 4097 36219 4131
rect 36219 4097 36228 4131
rect 36176 4088 36228 4097
rect 36820 4131 36872 4140
rect 36820 4097 36829 4131
rect 36829 4097 36863 4131
rect 36863 4097 36872 4131
rect 36820 4088 36872 4097
rect 38200 4131 38252 4140
rect 38200 4097 38209 4131
rect 38209 4097 38243 4131
rect 38243 4097 38252 4131
rect 38200 4088 38252 4097
rect 38568 4088 38620 4140
rect 38660 4131 38712 4140
rect 38660 4097 38669 4131
rect 38669 4097 38703 4131
rect 38703 4097 38712 4131
rect 38660 4088 38712 4097
rect 37280 4063 37332 4072
rect 37280 4029 37289 4063
rect 37289 4029 37323 4063
rect 37323 4029 37332 4063
rect 37280 4020 37332 4029
rect 38108 4020 38160 4072
rect 41604 4020 41656 4072
rect 41696 4063 41748 4072
rect 41696 4029 41705 4063
rect 41705 4029 41739 4063
rect 41739 4029 41748 4063
rect 41696 4020 41748 4029
rect 42800 4020 42852 4072
rect 43076 4020 43128 4072
rect 43812 4020 43864 4072
rect 44824 4063 44876 4072
rect 44824 4029 44833 4063
rect 44833 4029 44867 4063
rect 44867 4029 44876 4063
rect 44824 4020 44876 4029
rect 44916 4063 44968 4072
rect 44916 4029 44925 4063
rect 44925 4029 44959 4063
rect 44959 4029 44968 4063
rect 44916 4020 44968 4029
rect 42248 3952 42300 4004
rect 43260 3952 43312 4004
rect 36452 3884 36504 3936
rect 37188 3884 37240 3936
rect 38936 3884 38988 3936
rect 42892 3884 42944 3936
rect 43536 3884 43588 3936
rect 50528 4131 50580 4140
rect 50528 4097 50537 4131
rect 50537 4097 50571 4131
rect 50571 4097 50580 4131
rect 50528 4088 50580 4097
rect 74632 4088 74684 4140
rect 46940 4063 46992 4072
rect 46940 4029 46949 4063
rect 46949 4029 46983 4063
rect 46983 4029 46992 4063
rect 46940 4020 46992 4029
rect 47124 4063 47176 4072
rect 47124 4029 47133 4063
rect 47133 4029 47167 4063
rect 47167 4029 47176 4063
rect 47124 4020 47176 4029
rect 47216 4020 47268 4072
rect 48596 4020 48648 4072
rect 50068 4020 50120 4072
rect 65432 4020 65484 4072
rect 67916 4020 67968 4072
rect 71688 4020 71740 4072
rect 74080 4020 74132 4072
rect 76564 4020 76616 4072
rect 77024 4063 77076 4072
rect 77024 4029 77033 4063
rect 77033 4029 77067 4063
rect 77067 4029 77076 4063
rect 77024 4020 77076 4029
rect 48872 3952 48924 4004
rect 46112 3884 46164 3936
rect 46388 3927 46440 3936
rect 46388 3893 46397 3927
rect 46397 3893 46431 3927
rect 46431 3893 46440 3927
rect 46388 3884 46440 3893
rect 47492 3884 47544 3936
rect 49240 3927 49292 3936
rect 49240 3893 49249 3927
rect 49249 3893 49283 3927
rect 49283 3893 49292 3927
rect 49240 3884 49292 3893
rect 49884 3884 49936 3936
rect 51080 3884 51132 3936
rect 52368 3884 52420 3936
rect 66260 3884 66312 3936
rect 68284 3884 68336 3936
rect 72424 3884 72476 3936
rect 5134 3782 5186 3834
rect 5198 3782 5250 3834
rect 5262 3782 5314 3834
rect 5326 3782 5378 3834
rect 5390 3782 5442 3834
rect 35854 3782 35906 3834
rect 35918 3782 35970 3834
rect 35982 3782 36034 3834
rect 36046 3782 36098 3834
rect 36110 3782 36162 3834
rect 66574 3782 66626 3834
rect 66638 3782 66690 3834
rect 66702 3782 66754 3834
rect 66766 3782 66818 3834
rect 66830 3782 66882 3834
rect 5724 3680 5776 3732
rect 6000 3723 6052 3732
rect 6000 3689 6009 3723
rect 6009 3689 6043 3723
rect 6043 3689 6052 3723
rect 6000 3680 6052 3689
rect 8300 3612 8352 3664
rect 9864 3680 9916 3732
rect 11888 3723 11940 3732
rect 11888 3689 11897 3723
rect 11897 3689 11931 3723
rect 11931 3689 11940 3723
rect 11888 3680 11940 3689
rect 10692 3612 10744 3664
rect 14096 3655 14148 3664
rect 14096 3621 14105 3655
rect 14105 3621 14139 3655
rect 14139 3621 14148 3655
rect 14096 3612 14148 3621
rect 16580 3680 16632 3732
rect 16764 3680 16816 3732
rect 16488 3612 16540 3664
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 6276 3544 6328 3596
rect 6828 3587 6880 3596
rect 6828 3553 6837 3587
rect 6837 3553 6871 3587
rect 6871 3553 6880 3587
rect 6828 3544 6880 3553
rect 5632 3476 5684 3528
rect 6184 3476 6236 3528
rect 9128 3544 9180 3596
rect 12808 3544 12860 3596
rect 14280 3587 14332 3596
rect 14280 3553 14289 3587
rect 14289 3553 14323 3587
rect 14323 3553 14332 3587
rect 14280 3544 14332 3553
rect 15476 3587 15528 3596
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 15752 3544 15804 3596
rect 17316 3544 17368 3596
rect 19432 3612 19484 3664
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 9772 3476 9824 3528
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 7472 3408 7524 3460
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 14004 3476 14056 3528
rect 15292 3476 15344 3528
rect 12164 3408 12216 3460
rect 12716 3408 12768 3460
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 10140 3340 10192 3392
rect 11428 3340 11480 3392
rect 15936 3451 15988 3460
rect 15936 3417 15945 3451
rect 15945 3417 15979 3451
rect 15979 3417 15988 3451
rect 15936 3408 15988 3417
rect 13728 3340 13780 3392
rect 16212 3383 16264 3392
rect 16212 3349 16221 3383
rect 16221 3349 16255 3383
rect 16255 3349 16264 3383
rect 16212 3340 16264 3349
rect 16396 3383 16448 3392
rect 16396 3349 16405 3383
rect 16405 3349 16439 3383
rect 16439 3349 16448 3383
rect 16396 3340 16448 3349
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 18236 3519 18288 3528
rect 18236 3485 18245 3519
rect 18245 3485 18279 3519
rect 18279 3485 18288 3519
rect 18236 3476 18288 3485
rect 16856 3408 16908 3460
rect 17960 3408 18012 3460
rect 22100 3680 22152 3732
rect 20076 3612 20128 3664
rect 21456 3612 21508 3664
rect 24216 3612 24268 3664
rect 20812 3587 20864 3596
rect 20812 3553 20821 3587
rect 20821 3553 20855 3587
rect 20855 3553 20864 3587
rect 20812 3544 20864 3553
rect 22836 3587 22888 3596
rect 22836 3553 22845 3587
rect 22845 3553 22879 3587
rect 22879 3553 22888 3587
rect 22836 3544 22888 3553
rect 20352 3519 20404 3528
rect 20352 3485 20361 3519
rect 20361 3485 20395 3519
rect 20395 3485 20404 3519
rect 20352 3476 20404 3485
rect 20444 3476 20496 3528
rect 23204 3476 23256 3528
rect 24400 3476 24452 3528
rect 24676 3476 24728 3528
rect 25596 3655 25648 3664
rect 25596 3621 25605 3655
rect 25605 3621 25639 3655
rect 25639 3621 25648 3655
rect 25596 3612 25648 3621
rect 26148 3587 26200 3596
rect 26148 3553 26157 3587
rect 26157 3553 26191 3587
rect 26191 3553 26200 3587
rect 26148 3544 26200 3553
rect 27620 3544 27672 3596
rect 18604 3340 18656 3392
rect 20076 3340 20128 3392
rect 21824 3340 21876 3392
rect 22100 3408 22152 3460
rect 22468 3408 22520 3460
rect 24124 3408 24176 3460
rect 26608 3476 26660 3528
rect 28356 3680 28408 3732
rect 28724 3723 28776 3732
rect 28724 3689 28733 3723
rect 28733 3689 28767 3723
rect 28767 3689 28776 3723
rect 28724 3680 28776 3689
rect 30288 3680 30340 3732
rect 33324 3680 33376 3732
rect 34244 3723 34296 3732
rect 34244 3689 34253 3723
rect 34253 3689 34287 3723
rect 34287 3689 34296 3723
rect 34244 3680 34296 3689
rect 34796 3680 34848 3732
rect 35716 3680 35768 3732
rect 36452 3680 36504 3732
rect 40316 3680 40368 3732
rect 31852 3612 31904 3664
rect 32036 3612 32088 3664
rect 28356 3544 28408 3596
rect 30380 3544 30432 3596
rect 31300 3544 31352 3596
rect 32772 3544 32824 3596
rect 38936 3612 38988 3664
rect 29092 3519 29144 3528
rect 29092 3485 29101 3519
rect 29101 3485 29135 3519
rect 29135 3485 29144 3519
rect 29092 3476 29144 3485
rect 30288 3476 30340 3528
rect 30748 3476 30800 3528
rect 31208 3476 31260 3528
rect 34428 3519 34480 3528
rect 34428 3485 34437 3519
rect 34437 3485 34471 3519
rect 34471 3485 34480 3519
rect 34428 3476 34480 3485
rect 35164 3544 35216 3596
rect 35440 3544 35492 3596
rect 22744 3340 22796 3392
rect 23388 3340 23440 3392
rect 24492 3340 24544 3392
rect 25412 3383 25464 3392
rect 25412 3349 25421 3383
rect 25421 3349 25455 3383
rect 25455 3349 25464 3383
rect 25412 3340 25464 3349
rect 25688 3383 25740 3392
rect 25688 3349 25697 3383
rect 25697 3349 25731 3383
rect 25731 3349 25740 3383
rect 25688 3340 25740 3349
rect 26884 3408 26936 3460
rect 26148 3340 26200 3392
rect 26332 3340 26384 3392
rect 26700 3340 26752 3392
rect 26792 3340 26844 3392
rect 28540 3408 28592 3460
rect 30196 3408 30248 3460
rect 30380 3408 30432 3460
rect 30564 3408 30616 3460
rect 31852 3408 31904 3460
rect 32404 3408 32456 3460
rect 32956 3408 33008 3460
rect 27988 3340 28040 3392
rect 30472 3340 30524 3392
rect 30656 3340 30708 3392
rect 34980 3408 35032 3460
rect 35072 3451 35124 3460
rect 35072 3417 35081 3451
rect 35081 3417 35115 3451
rect 35115 3417 35124 3451
rect 35072 3408 35124 3417
rect 35716 3451 35768 3460
rect 35716 3417 35725 3451
rect 35725 3417 35759 3451
rect 35759 3417 35768 3451
rect 35716 3408 35768 3417
rect 36636 3476 36688 3528
rect 36820 3587 36872 3596
rect 36820 3553 36829 3587
rect 36829 3553 36863 3587
rect 36863 3553 36872 3587
rect 36820 3544 36872 3553
rect 38660 3587 38712 3596
rect 38660 3553 38669 3587
rect 38669 3553 38703 3587
rect 38703 3553 38712 3587
rect 38660 3544 38712 3553
rect 37924 3408 37976 3460
rect 34612 3340 34664 3392
rect 37096 3340 37148 3392
rect 38752 3340 38804 3392
rect 39764 3544 39816 3596
rect 46940 3680 46992 3732
rect 48780 3680 48832 3732
rect 67916 3723 67968 3732
rect 67916 3689 67925 3723
rect 67925 3689 67959 3723
rect 67959 3689 67968 3723
rect 67916 3680 67968 3689
rect 71688 3723 71740 3732
rect 71688 3689 71697 3723
rect 71697 3689 71731 3723
rect 71731 3689 71740 3723
rect 71688 3680 71740 3689
rect 77576 3723 77628 3732
rect 77576 3689 77585 3723
rect 77585 3689 77619 3723
rect 77619 3689 77628 3723
rect 77576 3680 77628 3689
rect 40316 3476 40368 3528
rect 42248 3587 42300 3596
rect 42248 3553 42257 3587
rect 42257 3553 42291 3587
rect 42291 3553 42300 3587
rect 42248 3544 42300 3553
rect 46388 3612 46440 3664
rect 39948 3340 40000 3392
rect 41144 3383 41196 3392
rect 41144 3349 41153 3383
rect 41153 3349 41187 3383
rect 41187 3349 41196 3383
rect 41144 3340 41196 3349
rect 41236 3383 41288 3392
rect 41236 3349 41245 3383
rect 41245 3349 41279 3383
rect 41279 3349 41288 3383
rect 41236 3340 41288 3349
rect 42064 3476 42116 3528
rect 44272 3587 44324 3596
rect 44272 3553 44281 3587
rect 44281 3553 44315 3587
rect 44315 3553 44324 3587
rect 44272 3544 44324 3553
rect 45560 3544 45612 3596
rect 45744 3544 45796 3596
rect 46296 3476 46348 3528
rect 46480 3519 46532 3528
rect 46480 3485 46489 3519
rect 46489 3485 46523 3519
rect 46523 3485 46532 3519
rect 46480 3476 46532 3485
rect 46664 3476 46716 3528
rect 72424 3587 72476 3596
rect 72424 3553 72433 3587
rect 72433 3553 72467 3587
rect 72467 3553 72476 3587
rect 72424 3544 72476 3553
rect 77024 3587 77076 3596
rect 77024 3553 77033 3587
rect 77033 3553 77067 3587
rect 77067 3553 77076 3587
rect 77024 3544 77076 3553
rect 46940 3476 46992 3528
rect 49792 3519 49844 3528
rect 49792 3485 49801 3519
rect 49801 3485 49835 3519
rect 49835 3485 49844 3519
rect 49792 3476 49844 3485
rect 51264 3476 51316 3528
rect 52460 3519 52512 3528
rect 52460 3485 52469 3519
rect 52469 3485 52503 3519
rect 52503 3485 52512 3519
rect 52460 3476 52512 3485
rect 53656 3519 53708 3528
rect 53656 3485 53665 3519
rect 53665 3485 53699 3519
rect 53699 3485 53708 3519
rect 53656 3476 53708 3485
rect 57336 3476 57388 3528
rect 58072 3476 58124 3528
rect 60924 3476 60976 3528
rect 62120 3519 62172 3528
rect 62120 3485 62129 3519
rect 62129 3485 62163 3519
rect 62163 3485 62172 3519
rect 62120 3476 62172 3485
rect 64696 3476 64748 3528
rect 67088 3476 67140 3528
rect 69112 3519 69164 3528
rect 69112 3485 69121 3519
rect 69121 3485 69155 3519
rect 69155 3485 69164 3519
rect 69112 3476 69164 3485
rect 72240 3519 72292 3528
rect 72240 3485 72249 3519
rect 72249 3485 72283 3519
rect 72283 3485 72292 3519
rect 72240 3476 72292 3485
rect 74448 3476 74500 3528
rect 76656 3519 76708 3528
rect 76656 3485 76665 3519
rect 76665 3485 76699 3519
rect 76699 3485 76708 3519
rect 76656 3476 76708 3485
rect 41696 3408 41748 3460
rect 42800 3408 42852 3460
rect 42984 3408 43036 3460
rect 46848 3408 46900 3460
rect 75460 3451 75512 3460
rect 75460 3417 75469 3451
rect 75469 3417 75503 3451
rect 75503 3417 75512 3451
rect 75460 3408 75512 3417
rect 44272 3340 44324 3392
rect 44916 3383 44968 3392
rect 44916 3349 44925 3383
rect 44925 3349 44959 3383
rect 44959 3349 44968 3383
rect 44916 3340 44968 3349
rect 48596 3340 48648 3392
rect 50620 3383 50672 3392
rect 50620 3349 50629 3383
rect 50629 3349 50663 3383
rect 50663 3349 50672 3383
rect 50620 3340 50672 3349
rect 51448 3340 51500 3392
rect 53012 3340 53064 3392
rect 56048 3340 56100 3392
rect 57428 3383 57480 3392
rect 57428 3349 57437 3383
rect 57437 3349 57471 3383
rect 57471 3349 57480 3383
rect 57428 3340 57480 3349
rect 58624 3340 58676 3392
rect 61108 3340 61160 3392
rect 62764 3383 62816 3392
rect 62764 3349 62773 3383
rect 62773 3349 62807 3383
rect 62807 3349 62816 3383
rect 62764 3340 62816 3349
rect 64880 3340 64932 3392
rect 71504 3340 71556 3392
rect 73068 3383 73120 3392
rect 73068 3349 73077 3383
rect 73077 3349 73111 3383
rect 73111 3349 73120 3383
rect 73068 3340 73120 3349
rect 74540 3383 74592 3392
rect 74540 3349 74549 3383
rect 74549 3349 74583 3383
rect 74583 3349 74592 3383
rect 74540 3340 74592 3349
rect 5794 3238 5846 3290
rect 5858 3238 5910 3290
rect 5922 3238 5974 3290
rect 5986 3238 6038 3290
rect 6050 3238 6102 3290
rect 36514 3238 36566 3290
rect 36578 3238 36630 3290
rect 36642 3238 36694 3290
rect 36706 3238 36758 3290
rect 36770 3238 36822 3290
rect 67234 3238 67286 3290
rect 67298 3238 67350 3290
rect 67362 3238 67414 3290
rect 67426 3238 67478 3290
rect 67490 3238 67542 3290
rect 4896 3179 4948 3188
rect 4896 3145 4905 3179
rect 4905 3145 4939 3179
rect 4939 3145 4948 3179
rect 4896 3136 4948 3145
rect 7840 3136 7892 3188
rect 9128 3136 9180 3188
rect 9404 3136 9456 3188
rect 6736 3068 6788 3120
rect 10600 3136 10652 3188
rect 12164 3136 12216 3188
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 5540 3000 5592 3052
rect 7012 3000 7064 3052
rect 8300 3000 8352 3052
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9680 3000 9732 3052
rect 11336 3068 11388 3120
rect 12900 3136 12952 3188
rect 10416 3000 10468 3052
rect 10508 3043 10560 3052
rect 10508 3009 10517 3043
rect 10517 3009 10551 3043
rect 10551 3009 10560 3043
rect 10508 3000 10560 3009
rect 7564 2932 7616 2984
rect 8852 2932 8904 2984
rect 11428 2932 11480 2984
rect 11520 2932 11572 2984
rect 8024 2864 8076 2916
rect 10508 2864 10560 2916
rect 7656 2796 7708 2848
rect 12716 2796 12768 2848
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 13360 3111 13412 3120
rect 13360 3077 13369 3111
rect 13369 3077 13403 3111
rect 13403 3077 13412 3111
rect 13360 3068 13412 3077
rect 13636 3068 13688 3120
rect 15384 3136 15436 3188
rect 18144 3136 18196 3188
rect 15660 3068 15712 3120
rect 17776 3068 17828 3120
rect 16488 3000 16540 3052
rect 18604 3111 18656 3120
rect 18604 3077 18613 3111
rect 18613 3077 18647 3111
rect 18647 3077 18656 3111
rect 18604 3068 18656 3077
rect 19892 3136 19944 3188
rect 19984 3136 20036 3188
rect 20168 3136 20220 3188
rect 19064 3068 19116 3120
rect 21732 3068 21784 3120
rect 22008 3111 22060 3120
rect 22008 3077 22017 3111
rect 22017 3077 22051 3111
rect 22051 3077 22060 3111
rect 22008 3068 22060 3077
rect 22100 3068 22152 3120
rect 22376 3111 22428 3120
rect 22376 3077 22385 3111
rect 22385 3077 22419 3111
rect 22419 3077 22428 3111
rect 22376 3068 22428 3077
rect 22744 3111 22796 3120
rect 22744 3077 22753 3111
rect 22753 3077 22787 3111
rect 22787 3077 22796 3111
rect 22744 3068 22796 3077
rect 23204 3136 23256 3188
rect 25228 3136 25280 3188
rect 26608 3136 26660 3188
rect 26884 3136 26936 3188
rect 27344 3136 27396 3188
rect 28172 3136 28224 3188
rect 28264 3136 28316 3188
rect 30472 3179 30524 3188
rect 30472 3145 30481 3179
rect 30481 3145 30515 3179
rect 30515 3145 30524 3179
rect 30472 3136 30524 3145
rect 32680 3179 32732 3188
rect 32680 3145 32689 3179
rect 32689 3145 32723 3179
rect 32723 3145 32732 3179
rect 32680 3136 32732 3145
rect 33324 3136 33376 3188
rect 33508 3179 33560 3188
rect 33508 3145 33517 3179
rect 33517 3145 33551 3179
rect 33551 3145 33560 3179
rect 33508 3136 33560 3145
rect 34060 3179 34112 3188
rect 34060 3145 34069 3179
rect 34069 3145 34103 3179
rect 34103 3145 34112 3179
rect 34060 3136 34112 3145
rect 34612 3136 34664 3188
rect 13452 2932 13504 2984
rect 13820 2932 13872 2984
rect 15568 2932 15620 2984
rect 16948 2932 17000 2984
rect 17500 2932 17552 2984
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 22284 3000 22336 3009
rect 23112 3000 23164 3052
rect 23572 3068 23624 3120
rect 25872 3068 25924 3120
rect 27804 3068 27856 3120
rect 24584 3000 24636 3052
rect 25044 3043 25096 3052
rect 25044 3009 25053 3043
rect 25053 3009 25087 3043
rect 25087 3009 25096 3043
rect 25044 3000 25096 3009
rect 25228 3000 25280 3052
rect 27252 3043 27304 3052
rect 27252 3009 27261 3043
rect 27261 3009 27295 3043
rect 27295 3009 27304 3043
rect 27252 3000 27304 3009
rect 27344 3043 27396 3052
rect 27344 3009 27353 3043
rect 27353 3009 27387 3043
rect 27387 3009 27396 3043
rect 27344 3000 27396 3009
rect 27988 3000 28040 3052
rect 28724 3068 28776 3120
rect 30012 3111 30064 3120
rect 30012 3077 30021 3111
rect 30021 3077 30055 3111
rect 30055 3077 30064 3111
rect 30012 3068 30064 3077
rect 14556 2796 14608 2848
rect 15292 2796 15344 2848
rect 16856 2796 16908 2848
rect 21456 2864 21508 2916
rect 23572 2932 23624 2984
rect 27160 2932 27212 2984
rect 28080 2932 28132 2984
rect 28540 3000 28592 3052
rect 29276 2932 29328 2984
rect 24676 2864 24728 2916
rect 20536 2796 20588 2848
rect 21088 2796 21140 2848
rect 22928 2839 22980 2848
rect 22928 2805 22937 2839
rect 22937 2805 22971 2839
rect 22971 2805 22980 2839
rect 22928 2796 22980 2805
rect 24860 2796 24912 2848
rect 25136 2796 25188 2848
rect 25228 2839 25280 2848
rect 25228 2805 25237 2839
rect 25237 2805 25271 2839
rect 25271 2805 25280 2839
rect 25228 2796 25280 2805
rect 31116 3068 31168 3120
rect 31208 3111 31260 3120
rect 31208 3077 31217 3111
rect 31217 3077 31251 3111
rect 31251 3077 31260 3111
rect 31208 3068 31260 3077
rect 32956 3068 33008 3120
rect 33140 3068 33192 3120
rect 35808 3136 35860 3188
rect 31300 2932 31352 2984
rect 32220 2932 32272 2984
rect 33784 3000 33836 3052
rect 33876 3043 33928 3052
rect 33876 3009 33885 3043
rect 33885 3009 33919 3043
rect 33919 3009 33928 3043
rect 33876 3000 33928 3009
rect 35624 3111 35676 3120
rect 35624 3077 35633 3111
rect 35633 3077 35667 3111
rect 35667 3077 35676 3111
rect 35624 3068 35676 3077
rect 37832 3136 37884 3188
rect 37556 3068 37608 3120
rect 37648 3111 37700 3120
rect 37648 3077 37657 3111
rect 37657 3077 37691 3111
rect 37691 3077 37700 3111
rect 37648 3068 37700 3077
rect 38476 3136 38528 3188
rect 41144 3136 41196 3188
rect 41696 3136 41748 3188
rect 42340 3136 42392 3188
rect 44824 3136 44876 3188
rect 45376 3179 45428 3188
rect 45376 3145 45385 3179
rect 45385 3145 45419 3179
rect 45419 3145 45428 3179
rect 45376 3136 45428 3145
rect 45928 3136 45980 3188
rect 48044 3179 48096 3188
rect 48044 3145 48053 3179
rect 48053 3145 48087 3179
rect 48087 3145 48096 3179
rect 48044 3136 48096 3145
rect 50068 3179 50120 3188
rect 50068 3145 50077 3179
rect 50077 3145 50111 3179
rect 50111 3145 50120 3179
rect 50068 3136 50120 3145
rect 51264 3179 51316 3188
rect 51264 3145 51273 3179
rect 51273 3145 51307 3179
rect 51307 3145 51316 3179
rect 51264 3136 51316 3145
rect 52460 3136 52512 3188
rect 53656 3179 53708 3188
rect 53656 3145 53665 3179
rect 53665 3145 53699 3179
rect 53699 3145 53708 3179
rect 53656 3136 53708 3145
rect 57336 3179 57388 3188
rect 57336 3145 57345 3179
rect 57345 3145 57379 3179
rect 57379 3145 57388 3179
rect 57336 3136 57388 3145
rect 58072 3179 58124 3188
rect 58072 3145 58081 3179
rect 58081 3145 58115 3179
rect 58115 3145 58124 3179
rect 58072 3136 58124 3145
rect 60924 3179 60976 3188
rect 60924 3145 60933 3179
rect 60933 3145 60967 3179
rect 60967 3145 60976 3179
rect 60924 3136 60976 3145
rect 62120 3136 62172 3188
rect 64696 3179 64748 3188
rect 64696 3145 64705 3179
rect 64705 3145 64739 3179
rect 64739 3145 64748 3179
rect 64696 3136 64748 3145
rect 65432 3179 65484 3188
rect 65432 3145 65441 3179
rect 65441 3145 65475 3179
rect 65475 3145 65484 3179
rect 65432 3136 65484 3145
rect 67088 3136 67140 3188
rect 69112 3179 69164 3188
rect 69112 3145 69121 3179
rect 69121 3145 69155 3179
rect 69155 3145 69164 3179
rect 69112 3136 69164 3145
rect 74448 3179 74500 3188
rect 74448 3145 74457 3179
rect 74457 3145 74491 3179
rect 74491 3145 74500 3179
rect 74448 3136 74500 3145
rect 35992 3000 36044 3052
rect 36268 3000 36320 3052
rect 29920 2796 29972 2848
rect 30380 2796 30432 2848
rect 30564 2796 30616 2848
rect 30840 2839 30892 2848
rect 30840 2805 30849 2839
rect 30849 2805 30883 2839
rect 30883 2805 30892 2839
rect 30840 2796 30892 2805
rect 33048 2907 33100 2916
rect 33048 2873 33057 2907
rect 33057 2873 33091 2907
rect 33091 2873 33100 2907
rect 33048 2864 33100 2873
rect 34612 2932 34664 2984
rect 40040 3000 40092 3052
rect 40960 3043 41012 3052
rect 40960 3009 40969 3043
rect 40969 3009 41003 3043
rect 41003 3009 41012 3043
rect 40960 3000 41012 3009
rect 42984 3068 43036 3120
rect 43812 3111 43864 3120
rect 43812 3077 43821 3111
rect 43821 3077 43855 3111
rect 43855 3077 43864 3111
rect 43812 3068 43864 3077
rect 45100 3068 45152 3120
rect 46940 3068 46992 3120
rect 43352 3000 43404 3052
rect 38384 2932 38436 2984
rect 40316 2932 40368 2984
rect 42156 2932 42208 2984
rect 45652 3000 45704 3052
rect 45836 3043 45888 3052
rect 45836 3009 45845 3043
rect 45845 3009 45879 3043
rect 45879 3009 45888 3043
rect 45836 3000 45888 3009
rect 46112 3043 46164 3052
rect 46112 3009 46121 3043
rect 46121 3009 46155 3043
rect 46155 3009 46164 3043
rect 46112 3000 46164 3009
rect 47492 3043 47544 3052
rect 47492 3009 47501 3043
rect 47501 3009 47535 3043
rect 47535 3009 47544 3043
rect 47492 3000 47544 3009
rect 49240 3000 49292 3052
rect 49792 3043 49844 3052
rect 49792 3009 49801 3043
rect 49801 3009 49835 3043
rect 49835 3009 49844 3043
rect 49792 3000 49844 3009
rect 50620 3043 50672 3052
rect 50620 3009 50629 3043
rect 50629 3009 50663 3043
rect 50663 3009 50672 3043
rect 50620 3000 50672 3009
rect 51080 3043 51132 3052
rect 51080 3009 51089 3043
rect 51089 3009 51123 3043
rect 51123 3009 51132 3043
rect 51080 3000 51132 3009
rect 51448 3043 51500 3052
rect 51448 3009 51457 3043
rect 51457 3009 51491 3043
rect 51491 3009 51500 3043
rect 51448 3000 51500 3009
rect 52092 3043 52144 3052
rect 52092 3009 52101 3043
rect 52101 3009 52135 3043
rect 52135 3009 52144 3043
rect 52092 3000 52144 3009
rect 52368 3000 52420 3052
rect 54024 3043 54076 3052
rect 54024 3009 54033 3043
rect 54033 3009 54067 3043
rect 54067 3009 54076 3043
rect 54024 3000 54076 3009
rect 56048 3043 56100 3052
rect 56048 3009 56057 3043
rect 56057 3009 56091 3043
rect 56091 3009 56100 3043
rect 56048 3000 56100 3009
rect 57428 3043 57480 3052
rect 57428 3009 57437 3043
rect 57437 3009 57471 3043
rect 57471 3009 57480 3043
rect 57428 3000 57480 3009
rect 61108 3043 61160 3052
rect 61108 3009 61117 3043
rect 61117 3009 61151 3043
rect 61151 3009 61160 3043
rect 61108 3000 61160 3009
rect 61752 3043 61804 3052
rect 61752 3009 61761 3043
rect 61761 3009 61795 3043
rect 61795 3009 61804 3043
rect 61752 3000 61804 3009
rect 64880 3043 64932 3052
rect 64880 3009 64889 3043
rect 64889 3009 64923 3043
rect 64923 3009 64932 3043
rect 64880 3000 64932 3009
rect 65524 3043 65576 3052
rect 65524 3009 65533 3043
rect 65533 3009 65567 3043
rect 65567 3009 65576 3043
rect 65524 3000 65576 3009
rect 67640 3043 67692 3052
rect 67640 3009 67649 3043
rect 67649 3009 67683 3043
rect 67683 3009 67692 3043
rect 67640 3000 67692 3009
rect 70308 3068 70360 3120
rect 69480 3043 69532 3052
rect 69480 3009 69489 3043
rect 69489 3009 69523 3043
rect 69523 3009 69532 3043
rect 69480 3000 69532 3009
rect 71504 3043 71556 3052
rect 71504 3009 71513 3043
rect 71513 3009 71547 3043
rect 71547 3009 71556 3043
rect 71504 3000 71556 3009
rect 72608 3000 72660 3052
rect 74080 3000 74132 3052
rect 74540 3043 74592 3052
rect 74540 3009 74549 3043
rect 74549 3009 74583 3043
rect 74583 3009 74592 3043
rect 74540 3000 74592 3009
rect 76656 3043 76708 3052
rect 76656 3009 76665 3043
rect 76665 3009 76699 3043
rect 76699 3009 76708 3043
rect 76656 3000 76708 3009
rect 34428 2864 34480 2916
rect 34888 2796 34940 2848
rect 35072 2796 35124 2848
rect 35532 2796 35584 2848
rect 36176 2839 36228 2848
rect 36176 2805 36185 2839
rect 36185 2805 36219 2839
rect 36219 2805 36228 2839
rect 36176 2796 36228 2805
rect 41420 2864 41472 2916
rect 44916 2932 44968 2984
rect 45928 2932 45980 2984
rect 46480 2975 46532 2984
rect 46480 2941 46489 2975
rect 46489 2941 46523 2975
rect 46523 2941 46532 2975
rect 46480 2932 46532 2941
rect 47676 2932 47728 2984
rect 51540 2932 51592 2984
rect 53472 2932 53524 2984
rect 61200 2932 61252 2984
rect 65064 2932 65116 2984
rect 68928 2932 68980 2984
rect 70860 2932 70912 2984
rect 74724 2932 74776 2984
rect 45468 2864 45520 2916
rect 66996 2864 67048 2916
rect 42800 2796 42852 2848
rect 43536 2839 43588 2848
rect 43536 2805 43545 2839
rect 43545 2805 43579 2839
rect 43579 2805 43588 2839
rect 43536 2796 43588 2805
rect 55312 2796 55364 2848
rect 59268 2796 59320 2848
rect 70492 2796 70544 2848
rect 76196 2796 76248 2848
rect 5134 2694 5186 2746
rect 5198 2694 5250 2746
rect 5262 2694 5314 2746
rect 5326 2694 5378 2746
rect 5390 2694 5442 2746
rect 35854 2694 35906 2746
rect 35918 2694 35970 2746
rect 35982 2694 36034 2746
rect 36046 2694 36098 2746
rect 36110 2694 36162 2746
rect 66574 2694 66626 2746
rect 66638 2694 66690 2746
rect 66702 2694 66754 2746
rect 66766 2694 66818 2746
rect 66830 2694 66882 2746
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 4528 2635 4580 2644
rect 4528 2601 4537 2635
rect 4537 2601 4571 2635
rect 4571 2601 4580 2635
rect 4528 2592 4580 2601
rect 5632 2592 5684 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 9772 2592 9824 2644
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 8852 2524 8904 2576
rect 12716 2592 12768 2644
rect 11244 2567 11296 2576
rect 11244 2533 11253 2567
rect 11253 2533 11287 2567
rect 11287 2533 11296 2567
rect 11244 2524 11296 2533
rect 3976 2499 4028 2508
rect 3976 2465 3985 2499
rect 3985 2465 4019 2499
rect 4019 2465 4028 2499
rect 3976 2456 4028 2465
rect 5816 2499 5868 2508
rect 5816 2465 5825 2499
rect 5825 2465 5859 2499
rect 5859 2465 5868 2499
rect 5816 2456 5868 2465
rect 7932 2456 7984 2508
rect 10784 2456 10836 2508
rect 11060 2456 11112 2508
rect 11796 2499 11848 2508
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 3608 2431 3660 2440
rect 3608 2397 3617 2431
rect 3617 2397 3651 2431
rect 3651 2397 3660 2431
rect 3608 2388 3660 2397
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 6184 2388 6236 2440
rect 7656 2431 7708 2440
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 10416 2388 10468 2440
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 11520 2388 11572 2440
rect 13912 2524 13964 2576
rect 16856 2592 16908 2644
rect 17132 2592 17184 2644
rect 12624 2456 12676 2508
rect 12808 2431 12860 2440
rect 12808 2397 12817 2431
rect 12817 2397 12851 2431
rect 12851 2397 12860 2431
rect 12808 2388 12860 2397
rect 5632 2363 5684 2372
rect 5632 2329 5641 2363
rect 5641 2329 5675 2363
rect 5675 2329 5684 2363
rect 5632 2320 5684 2329
rect 10968 2320 11020 2372
rect 12992 2320 13044 2372
rect 8944 2295 8996 2304
rect 8944 2261 8953 2295
rect 8953 2261 8987 2295
rect 8987 2261 8996 2295
rect 8944 2252 8996 2261
rect 11704 2295 11756 2304
rect 11704 2261 11713 2295
rect 11713 2261 11747 2295
rect 11747 2261 11756 2295
rect 11704 2252 11756 2261
rect 11796 2252 11848 2304
rect 13544 2320 13596 2372
rect 14648 2431 14700 2440
rect 14648 2397 14657 2431
rect 14657 2397 14691 2431
rect 14691 2397 14700 2431
rect 14648 2388 14700 2397
rect 14832 2456 14884 2508
rect 16028 2524 16080 2576
rect 20260 2592 20312 2644
rect 24308 2592 24360 2644
rect 26516 2592 26568 2644
rect 34612 2592 34664 2644
rect 15752 2388 15804 2440
rect 19340 2499 19392 2508
rect 19340 2465 19349 2499
rect 19349 2465 19383 2499
rect 19383 2465 19392 2499
rect 19340 2456 19392 2465
rect 20720 2499 20772 2508
rect 20720 2465 20729 2499
rect 20729 2465 20763 2499
rect 20763 2465 20772 2499
rect 20720 2456 20772 2465
rect 22192 2456 22244 2508
rect 22836 2456 22888 2508
rect 23940 2456 23992 2508
rect 24400 2499 24452 2508
rect 24400 2465 24409 2499
rect 24409 2465 24443 2499
rect 24443 2465 24452 2499
rect 24400 2456 24452 2465
rect 24768 2456 24820 2508
rect 17868 2388 17920 2440
rect 20168 2431 20220 2440
rect 20168 2397 20177 2431
rect 20177 2397 20211 2431
rect 20211 2397 20220 2431
rect 20168 2388 20220 2397
rect 20352 2388 20404 2440
rect 16948 2320 17000 2372
rect 21548 2431 21600 2440
rect 21548 2397 21557 2431
rect 21557 2397 21591 2431
rect 21591 2397 21600 2431
rect 21548 2388 21600 2397
rect 22284 2388 22336 2440
rect 22560 2431 22612 2440
rect 22560 2397 22569 2431
rect 22569 2397 22603 2431
rect 22603 2397 22612 2431
rect 22560 2388 22612 2397
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 25320 2431 25372 2440
rect 25320 2397 25329 2431
rect 25329 2397 25363 2431
rect 25363 2397 25372 2431
rect 25320 2388 25372 2397
rect 26240 2499 26292 2508
rect 26240 2465 26249 2499
rect 26249 2465 26283 2499
rect 26283 2465 26292 2499
rect 26240 2456 26292 2465
rect 26424 2456 26476 2508
rect 34152 2524 34204 2576
rect 35808 2567 35860 2576
rect 35808 2533 35817 2567
rect 35817 2533 35851 2567
rect 35851 2533 35860 2567
rect 35808 2524 35860 2533
rect 30288 2456 30340 2508
rect 32220 2499 32272 2508
rect 32220 2465 32229 2499
rect 32229 2465 32263 2499
rect 32263 2465 32272 2499
rect 32220 2456 32272 2465
rect 41604 2592 41656 2644
rect 43536 2592 43588 2644
rect 44732 2592 44784 2644
rect 45836 2592 45888 2644
rect 46848 2592 46900 2644
rect 49976 2635 50028 2644
rect 49976 2601 49985 2635
rect 49985 2601 50019 2635
rect 50019 2601 50028 2635
rect 49976 2592 50028 2601
rect 72240 2592 72292 2644
rect 74632 2592 74684 2644
rect 76656 2592 76708 2644
rect 39856 2456 39908 2508
rect 40040 2456 40092 2508
rect 27896 2431 27948 2440
rect 27896 2397 27905 2431
rect 27905 2397 27939 2431
rect 27939 2397 27948 2431
rect 27896 2388 27948 2397
rect 26976 2320 27028 2372
rect 15200 2295 15252 2304
rect 15200 2261 15209 2295
rect 15209 2261 15243 2295
rect 15243 2261 15252 2295
rect 15200 2252 15252 2261
rect 15568 2295 15620 2304
rect 15568 2261 15577 2295
rect 15577 2261 15611 2295
rect 15611 2261 15620 2295
rect 15568 2252 15620 2261
rect 16396 2252 16448 2304
rect 18052 2295 18104 2304
rect 18052 2261 18061 2295
rect 18061 2261 18095 2295
rect 18095 2261 18104 2295
rect 18052 2252 18104 2261
rect 20352 2295 20404 2304
rect 20352 2261 20361 2295
rect 20361 2261 20395 2295
rect 20395 2261 20404 2295
rect 20352 2252 20404 2261
rect 20628 2295 20680 2304
rect 20628 2261 20637 2295
rect 20637 2261 20671 2295
rect 20671 2261 20680 2295
rect 20628 2252 20680 2261
rect 22100 2295 22152 2304
rect 22100 2261 22109 2295
rect 22109 2261 22143 2295
rect 22143 2261 22152 2295
rect 22100 2252 22152 2261
rect 22836 2252 22888 2304
rect 23848 2252 23900 2304
rect 30104 2388 30156 2440
rect 30380 2388 30432 2440
rect 32772 2388 32824 2440
rect 33324 2388 33376 2440
rect 35256 2431 35308 2440
rect 35256 2397 35265 2431
rect 35265 2397 35299 2431
rect 35299 2397 35308 2431
rect 35256 2388 35308 2397
rect 35624 2431 35676 2440
rect 35624 2397 35633 2431
rect 35633 2397 35667 2431
rect 35667 2397 35676 2431
rect 35624 2388 35676 2397
rect 35992 2431 36044 2440
rect 35992 2397 36001 2431
rect 36001 2397 36035 2431
rect 36035 2397 36044 2431
rect 35992 2388 36044 2397
rect 28816 2363 28868 2372
rect 28816 2329 28825 2363
rect 28825 2329 28859 2363
rect 28859 2329 28868 2363
rect 28816 2320 28868 2329
rect 34152 2320 34204 2372
rect 38016 2388 38068 2440
rect 38844 2431 38896 2440
rect 38844 2397 38853 2431
rect 38853 2397 38887 2431
rect 38887 2397 38896 2431
rect 38844 2388 38896 2397
rect 38936 2431 38988 2440
rect 38936 2397 38945 2431
rect 38945 2397 38979 2431
rect 38979 2397 38988 2431
rect 38936 2388 38988 2397
rect 41972 2524 42024 2576
rect 44640 2524 44692 2576
rect 49608 2524 49660 2576
rect 41144 2499 41196 2508
rect 41144 2465 41153 2499
rect 41153 2465 41187 2499
rect 41187 2465 41196 2499
rect 41144 2456 41196 2465
rect 41880 2456 41932 2508
rect 44272 2456 44324 2508
rect 38752 2320 38804 2372
rect 44824 2388 44876 2440
rect 45836 2388 45888 2440
rect 45928 2431 45980 2440
rect 45928 2397 45937 2431
rect 45937 2397 45971 2431
rect 45971 2397 45980 2431
rect 45928 2388 45980 2397
rect 42708 2320 42760 2372
rect 43812 2320 43864 2372
rect 47032 2456 47084 2508
rect 49792 2456 49844 2508
rect 52092 2499 52144 2508
rect 52092 2465 52101 2499
rect 52101 2465 52135 2499
rect 52135 2465 52144 2499
rect 52092 2456 52144 2465
rect 54024 2499 54076 2508
rect 54024 2465 54033 2499
rect 54033 2465 54067 2499
rect 54067 2465 54076 2499
rect 54024 2456 54076 2465
rect 48320 2431 48372 2440
rect 48320 2397 48329 2431
rect 48329 2397 48363 2431
rect 48363 2397 48372 2431
rect 48320 2388 48372 2397
rect 49884 2431 49936 2440
rect 49884 2397 49893 2431
rect 49893 2397 49927 2431
rect 49927 2397 49936 2431
rect 49884 2388 49936 2397
rect 50528 2431 50580 2440
rect 50528 2397 50537 2431
rect 50537 2397 50571 2431
rect 50571 2397 50580 2431
rect 50528 2388 50580 2397
rect 53012 2431 53064 2440
rect 53012 2397 53021 2431
rect 53021 2397 53055 2431
rect 53055 2397 53064 2431
rect 53012 2388 53064 2397
rect 55312 2388 55364 2440
rect 55404 2388 55456 2440
rect 58624 2431 58676 2440
rect 58624 2397 58633 2431
rect 58633 2397 58667 2431
rect 58667 2397 58676 2431
rect 58624 2388 58676 2397
rect 57336 2320 57388 2372
rect 61752 2499 61804 2508
rect 61752 2465 61761 2499
rect 61761 2465 61795 2499
rect 61795 2465 61804 2499
rect 61752 2456 61804 2465
rect 65524 2499 65576 2508
rect 65524 2465 65533 2499
rect 65533 2465 65567 2499
rect 65567 2465 65576 2499
rect 65524 2456 65576 2465
rect 67640 2499 67692 2508
rect 67640 2465 67649 2499
rect 67649 2465 67683 2499
rect 67683 2465 67692 2499
rect 67640 2456 67692 2465
rect 69480 2499 69532 2508
rect 69480 2465 69489 2499
rect 69489 2465 69523 2499
rect 69523 2465 69532 2499
rect 69480 2456 69532 2465
rect 70308 2456 70360 2508
rect 62764 2431 62816 2440
rect 62764 2397 62773 2431
rect 62773 2397 62807 2431
rect 62807 2397 62816 2431
rect 62764 2388 62816 2397
rect 63132 2388 63184 2440
rect 66260 2431 66312 2440
rect 66260 2397 66269 2431
rect 66269 2397 66303 2431
rect 66303 2397 66312 2431
rect 66260 2388 66312 2397
rect 68284 2431 68336 2440
rect 68284 2397 68293 2431
rect 68293 2397 68327 2431
rect 68327 2397 68336 2431
rect 68284 2388 68336 2397
rect 70492 2431 70544 2440
rect 70492 2397 70501 2431
rect 70501 2397 70535 2431
rect 70535 2397 70544 2431
rect 70492 2388 70544 2397
rect 72608 2499 72660 2508
rect 72608 2465 72617 2499
rect 72617 2465 72651 2499
rect 72651 2465 72660 2499
rect 72608 2456 72660 2465
rect 72792 2456 72844 2508
rect 75460 2456 75512 2508
rect 73068 2431 73120 2440
rect 73068 2397 73077 2431
rect 73077 2397 73111 2431
rect 73111 2397 73120 2431
rect 73068 2388 73120 2397
rect 76196 2431 76248 2440
rect 76196 2397 76205 2431
rect 76205 2397 76239 2431
rect 76239 2397 76248 2431
rect 76196 2388 76248 2397
rect 28080 2295 28132 2304
rect 28080 2261 28089 2295
rect 28089 2261 28123 2295
rect 28123 2261 28132 2295
rect 28080 2252 28132 2261
rect 31392 2295 31444 2304
rect 31392 2261 31401 2295
rect 31401 2261 31435 2295
rect 31435 2261 31444 2295
rect 31392 2252 31444 2261
rect 34980 2252 35032 2304
rect 47400 2295 47452 2304
rect 47400 2261 47409 2295
rect 47409 2261 47443 2295
rect 47443 2261 47452 2295
rect 47400 2252 47452 2261
rect 5794 2150 5846 2202
rect 5858 2150 5910 2202
rect 5922 2150 5974 2202
rect 5986 2150 6038 2202
rect 6050 2150 6102 2202
rect 36514 2150 36566 2202
rect 36578 2150 36630 2202
rect 36642 2150 36694 2202
rect 36706 2150 36758 2202
rect 36770 2150 36822 2202
rect 67234 2150 67286 2202
rect 67298 2150 67350 2202
rect 67362 2150 67414 2202
rect 67426 2150 67478 2202
rect 67490 2150 67542 2202
rect 6276 2048 6328 2100
rect 11612 2048 11664 2100
rect 12992 2048 13044 2100
rect 9128 1980 9180 2032
rect 16396 1980 16448 2032
rect 10600 1912 10652 1964
rect 13360 1912 13412 1964
rect 20628 2048 20680 2100
rect 27528 2048 27580 2100
rect 35992 2048 36044 2100
rect 47400 2048 47452 2100
rect 22100 1980 22152 2032
rect 23572 1912 23624 1964
rect 23848 1912 23900 1964
rect 30472 1912 30524 1964
rect 5724 1844 5776 1896
rect 11704 1844 11756 1896
rect 16304 1844 16356 1896
rect 8300 1776 8352 1828
rect 18052 1776 18104 1828
rect 20168 1776 20220 1828
rect 26332 1776 26384 1828
rect 8944 1708 8996 1760
rect 18144 1708 18196 1760
rect 8576 1640 8628 1692
rect 13360 1640 13412 1692
rect 25688 1640 25740 1692
rect 15200 1572 15252 1624
rect 20352 1572 20404 1624
rect 25780 1572 25832 1624
rect 31576 1980 31628 2032
rect 38936 1980 38988 2032
rect 44456 1980 44508 2032
rect 50528 1980 50580 2032
rect 35624 1912 35676 1964
rect 40684 1912 40736 1964
rect 35808 1844 35860 1896
rect 40500 1844 40552 1896
rect 32772 1776 32824 1828
rect 39212 1776 39264 1828
rect 31392 1708 31444 1760
rect 41236 1708 41288 1760
rect 36912 1640 36964 1692
rect 35716 1572 35768 1624
rect 14924 1300 14976 1352
rect 16120 1300 16172 1352
rect 42524 1300 42576 1352
rect 47124 1300 47176 1352
rect 40592 1096 40644 1148
rect 45192 1096 45244 1148
rect 7656 280 7708 332
rect 18604 280 18656 332
rect 21732 280 21784 332
rect 31484 280 31536 332
rect 10140 212 10192 264
rect 21180 212 21232 264
rect 21640 212 21692 264
rect 32772 212 32824 264
rect 8392 144 8444 196
rect 23112 144 23164 196
rect 9128 76 9180 128
rect 23480 76 23532 128
<< metal2 >>
rect 2226 39200 2282 40000
rect 4066 39200 4122 40000
rect 5906 39200 5962 40000
rect 7746 39200 7802 40000
rect 9586 39200 9642 40000
rect 11426 39200 11482 40000
rect 13266 39200 13322 40000
rect 15106 39200 15162 40000
rect 16946 39200 17002 40000
rect 18786 39200 18842 40000
rect 20626 39200 20682 40000
rect 22466 39200 22522 40000
rect 24306 39200 24362 40000
rect 26146 39200 26202 40000
rect 27986 39200 28042 40000
rect 29826 39200 29882 40000
rect 31666 39200 31722 40000
rect 33506 39200 33562 40000
rect 35346 39200 35402 40000
rect 37186 39200 37242 40000
rect 39026 39200 39082 40000
rect 40866 39200 40922 40000
rect 42706 39200 42762 40000
rect 44546 39200 44602 40000
rect 46386 39200 46442 40000
rect 48226 39200 48282 40000
rect 50066 39200 50122 40000
rect 51906 39200 51962 40000
rect 53746 39200 53802 40000
rect 55586 39200 55642 40000
rect 57426 39200 57482 40000
rect 59266 39200 59322 40000
rect 2240 37330 2268 39200
rect 2228 37324 2280 37330
rect 2228 37266 2280 37272
rect 3516 37256 3568 37262
rect 3516 37198 3568 37204
rect 3528 24177 3556 37198
rect 4080 36854 4108 39200
rect 5134 37564 5442 37573
rect 5134 37562 5140 37564
rect 5196 37562 5220 37564
rect 5276 37562 5300 37564
rect 5356 37562 5380 37564
rect 5436 37562 5442 37564
rect 5196 37510 5198 37562
rect 5378 37510 5380 37562
rect 5134 37508 5140 37510
rect 5196 37508 5220 37510
rect 5276 37508 5300 37510
rect 5356 37508 5380 37510
rect 5436 37508 5442 37510
rect 5134 37499 5442 37508
rect 5920 37262 5948 39200
rect 7760 37618 7788 39200
rect 7760 37590 7972 37618
rect 7944 37262 7972 37590
rect 5908 37256 5960 37262
rect 5908 37198 5960 37204
rect 7012 37256 7064 37262
rect 7012 37198 7064 37204
rect 7748 37256 7800 37262
rect 7748 37198 7800 37204
rect 7932 37256 7984 37262
rect 7932 37198 7984 37204
rect 5794 37020 6102 37029
rect 5794 37018 5800 37020
rect 5856 37018 5880 37020
rect 5936 37018 5960 37020
rect 6016 37018 6040 37020
rect 6096 37018 6102 37020
rect 5856 36966 5858 37018
rect 6038 36966 6040 37018
rect 5794 36964 5800 36966
rect 5856 36964 5880 36966
rect 5936 36964 5960 36966
rect 6016 36964 6040 36966
rect 6096 36964 6102 36966
rect 5794 36955 6102 36964
rect 4068 36848 4120 36854
rect 4068 36790 4120 36796
rect 7024 36553 7052 37198
rect 7760 36922 7788 37198
rect 7748 36916 7800 36922
rect 7748 36858 7800 36864
rect 9600 36854 9628 39200
rect 11440 37262 11468 39200
rect 13280 37330 13308 39200
rect 15120 37346 15148 39200
rect 13268 37324 13320 37330
rect 13268 37266 13320 37272
rect 15028 37318 15148 37346
rect 11428 37256 11480 37262
rect 11428 37198 11480 37204
rect 11888 37256 11940 37262
rect 11888 37198 11940 37204
rect 14556 37256 14608 37262
rect 14556 37198 14608 37204
rect 11900 36922 11928 37198
rect 11888 36916 11940 36922
rect 11888 36858 11940 36864
rect 9588 36848 9640 36854
rect 9588 36790 9640 36796
rect 10876 36780 10928 36786
rect 10876 36722 10928 36728
rect 11796 36780 11848 36786
rect 11796 36722 11848 36728
rect 7010 36544 7066 36553
rect 5134 36476 5442 36485
rect 7010 36479 7066 36488
rect 5134 36474 5140 36476
rect 5196 36474 5220 36476
rect 5276 36474 5300 36476
rect 5356 36474 5380 36476
rect 5436 36474 5442 36476
rect 5196 36422 5198 36474
rect 5378 36422 5380 36474
rect 5134 36420 5140 36422
rect 5196 36420 5220 36422
rect 5276 36420 5300 36422
rect 5356 36420 5380 36422
rect 5436 36420 5442 36422
rect 5134 36411 5442 36420
rect 5794 35932 6102 35941
rect 5794 35930 5800 35932
rect 5856 35930 5880 35932
rect 5936 35930 5960 35932
rect 6016 35930 6040 35932
rect 6096 35930 6102 35932
rect 5856 35878 5858 35930
rect 6038 35878 6040 35930
rect 5794 35876 5800 35878
rect 5856 35876 5880 35878
rect 5936 35876 5960 35878
rect 6016 35876 6040 35878
rect 6096 35876 6102 35878
rect 5794 35867 6102 35876
rect 5134 35388 5442 35397
rect 5134 35386 5140 35388
rect 5196 35386 5220 35388
rect 5276 35386 5300 35388
rect 5356 35386 5380 35388
rect 5436 35386 5442 35388
rect 5196 35334 5198 35386
rect 5378 35334 5380 35386
rect 5134 35332 5140 35334
rect 5196 35332 5220 35334
rect 5276 35332 5300 35334
rect 5356 35332 5380 35334
rect 5436 35332 5442 35334
rect 5134 35323 5442 35332
rect 5794 34844 6102 34853
rect 5794 34842 5800 34844
rect 5856 34842 5880 34844
rect 5936 34842 5960 34844
rect 6016 34842 6040 34844
rect 6096 34842 6102 34844
rect 5856 34790 5858 34842
rect 6038 34790 6040 34842
rect 5794 34788 5800 34790
rect 5856 34788 5880 34790
rect 5936 34788 5960 34790
rect 6016 34788 6040 34790
rect 6096 34788 6102 34790
rect 5794 34779 6102 34788
rect 5134 34300 5442 34309
rect 5134 34298 5140 34300
rect 5196 34298 5220 34300
rect 5276 34298 5300 34300
rect 5356 34298 5380 34300
rect 5436 34298 5442 34300
rect 5196 34246 5198 34298
rect 5378 34246 5380 34298
rect 5134 34244 5140 34246
rect 5196 34244 5220 34246
rect 5276 34244 5300 34246
rect 5356 34244 5380 34246
rect 5436 34244 5442 34246
rect 5134 34235 5442 34244
rect 5794 33756 6102 33765
rect 5794 33754 5800 33756
rect 5856 33754 5880 33756
rect 5936 33754 5960 33756
rect 6016 33754 6040 33756
rect 6096 33754 6102 33756
rect 5856 33702 5858 33754
rect 6038 33702 6040 33754
rect 5794 33700 5800 33702
rect 5856 33700 5880 33702
rect 5936 33700 5960 33702
rect 6016 33700 6040 33702
rect 6096 33700 6102 33702
rect 5794 33691 6102 33700
rect 5134 33212 5442 33221
rect 5134 33210 5140 33212
rect 5196 33210 5220 33212
rect 5276 33210 5300 33212
rect 5356 33210 5380 33212
rect 5436 33210 5442 33212
rect 5196 33158 5198 33210
rect 5378 33158 5380 33210
rect 5134 33156 5140 33158
rect 5196 33156 5220 33158
rect 5276 33156 5300 33158
rect 5356 33156 5380 33158
rect 5436 33156 5442 33158
rect 5134 33147 5442 33156
rect 5794 32668 6102 32677
rect 5794 32666 5800 32668
rect 5856 32666 5880 32668
rect 5936 32666 5960 32668
rect 6016 32666 6040 32668
rect 6096 32666 6102 32668
rect 5856 32614 5858 32666
rect 6038 32614 6040 32666
rect 5794 32612 5800 32614
rect 5856 32612 5880 32614
rect 5936 32612 5960 32614
rect 6016 32612 6040 32614
rect 6096 32612 6102 32614
rect 5794 32603 6102 32612
rect 5134 32124 5442 32133
rect 5134 32122 5140 32124
rect 5196 32122 5220 32124
rect 5276 32122 5300 32124
rect 5356 32122 5380 32124
rect 5436 32122 5442 32124
rect 5196 32070 5198 32122
rect 5378 32070 5380 32122
rect 5134 32068 5140 32070
rect 5196 32068 5220 32070
rect 5276 32068 5300 32070
rect 5356 32068 5380 32070
rect 5436 32068 5442 32070
rect 5134 32059 5442 32068
rect 5794 31580 6102 31589
rect 5794 31578 5800 31580
rect 5856 31578 5880 31580
rect 5936 31578 5960 31580
rect 6016 31578 6040 31580
rect 6096 31578 6102 31580
rect 5856 31526 5858 31578
rect 6038 31526 6040 31578
rect 5794 31524 5800 31526
rect 5856 31524 5880 31526
rect 5936 31524 5960 31526
rect 6016 31524 6040 31526
rect 6096 31524 6102 31526
rect 5794 31515 6102 31524
rect 5134 31036 5442 31045
rect 5134 31034 5140 31036
rect 5196 31034 5220 31036
rect 5276 31034 5300 31036
rect 5356 31034 5380 31036
rect 5436 31034 5442 31036
rect 5196 30982 5198 31034
rect 5378 30982 5380 31034
rect 5134 30980 5140 30982
rect 5196 30980 5220 30982
rect 5276 30980 5300 30982
rect 5356 30980 5380 30982
rect 5436 30980 5442 30982
rect 5134 30971 5442 30980
rect 5794 30492 6102 30501
rect 5794 30490 5800 30492
rect 5856 30490 5880 30492
rect 5936 30490 5960 30492
rect 6016 30490 6040 30492
rect 6096 30490 6102 30492
rect 5856 30438 5858 30490
rect 6038 30438 6040 30490
rect 5794 30436 5800 30438
rect 5856 30436 5880 30438
rect 5936 30436 5960 30438
rect 6016 30436 6040 30438
rect 6096 30436 6102 30438
rect 5794 30427 6102 30436
rect 5134 29948 5442 29957
rect 5134 29946 5140 29948
rect 5196 29946 5220 29948
rect 5276 29946 5300 29948
rect 5356 29946 5380 29948
rect 5436 29946 5442 29948
rect 5196 29894 5198 29946
rect 5378 29894 5380 29946
rect 5134 29892 5140 29894
rect 5196 29892 5220 29894
rect 5276 29892 5300 29894
rect 5356 29892 5380 29894
rect 5436 29892 5442 29894
rect 5134 29883 5442 29892
rect 5794 29404 6102 29413
rect 5794 29402 5800 29404
rect 5856 29402 5880 29404
rect 5936 29402 5960 29404
rect 6016 29402 6040 29404
rect 6096 29402 6102 29404
rect 5856 29350 5858 29402
rect 6038 29350 6040 29402
rect 5794 29348 5800 29350
rect 5856 29348 5880 29350
rect 5936 29348 5960 29350
rect 6016 29348 6040 29350
rect 6096 29348 6102 29350
rect 5794 29339 6102 29348
rect 5134 28860 5442 28869
rect 5134 28858 5140 28860
rect 5196 28858 5220 28860
rect 5276 28858 5300 28860
rect 5356 28858 5380 28860
rect 5436 28858 5442 28860
rect 5196 28806 5198 28858
rect 5378 28806 5380 28858
rect 5134 28804 5140 28806
rect 5196 28804 5220 28806
rect 5276 28804 5300 28806
rect 5356 28804 5380 28806
rect 5436 28804 5442 28806
rect 5134 28795 5442 28804
rect 5794 28316 6102 28325
rect 5794 28314 5800 28316
rect 5856 28314 5880 28316
rect 5936 28314 5960 28316
rect 6016 28314 6040 28316
rect 6096 28314 6102 28316
rect 5856 28262 5858 28314
rect 6038 28262 6040 28314
rect 5794 28260 5800 28262
rect 5856 28260 5880 28262
rect 5936 28260 5960 28262
rect 6016 28260 6040 28262
rect 6096 28260 6102 28262
rect 5794 28251 6102 28260
rect 5134 27772 5442 27781
rect 5134 27770 5140 27772
rect 5196 27770 5220 27772
rect 5276 27770 5300 27772
rect 5356 27770 5380 27772
rect 5436 27770 5442 27772
rect 5196 27718 5198 27770
rect 5378 27718 5380 27770
rect 5134 27716 5140 27718
rect 5196 27716 5220 27718
rect 5276 27716 5300 27718
rect 5356 27716 5380 27718
rect 5436 27716 5442 27718
rect 5134 27707 5442 27716
rect 5794 27228 6102 27237
rect 5794 27226 5800 27228
rect 5856 27226 5880 27228
rect 5936 27226 5960 27228
rect 6016 27226 6040 27228
rect 6096 27226 6102 27228
rect 5856 27174 5858 27226
rect 6038 27174 6040 27226
rect 5794 27172 5800 27174
rect 5856 27172 5880 27174
rect 5936 27172 5960 27174
rect 6016 27172 6040 27174
rect 6096 27172 6102 27174
rect 5794 27163 6102 27172
rect 10888 26897 10916 36722
rect 11808 36650 11836 36722
rect 11796 36644 11848 36650
rect 11796 36586 11848 36592
rect 10874 26888 10930 26897
rect 10874 26823 10930 26832
rect 5134 26684 5442 26693
rect 5134 26682 5140 26684
rect 5196 26682 5220 26684
rect 5276 26682 5300 26684
rect 5356 26682 5380 26684
rect 5436 26682 5442 26684
rect 5196 26630 5198 26682
rect 5378 26630 5380 26682
rect 5134 26628 5140 26630
rect 5196 26628 5220 26630
rect 5276 26628 5300 26630
rect 5356 26628 5380 26630
rect 5436 26628 5442 26630
rect 5134 26619 5442 26628
rect 5794 26140 6102 26149
rect 5794 26138 5800 26140
rect 5856 26138 5880 26140
rect 5936 26138 5960 26140
rect 6016 26138 6040 26140
rect 6096 26138 6102 26140
rect 5856 26086 5858 26138
rect 6038 26086 6040 26138
rect 5794 26084 5800 26086
rect 5856 26084 5880 26086
rect 5936 26084 5960 26086
rect 6016 26084 6040 26086
rect 6096 26084 6102 26086
rect 5794 26075 6102 26084
rect 5134 25596 5442 25605
rect 5134 25594 5140 25596
rect 5196 25594 5220 25596
rect 5276 25594 5300 25596
rect 5356 25594 5380 25596
rect 5436 25594 5442 25596
rect 5196 25542 5198 25594
rect 5378 25542 5380 25594
rect 5134 25540 5140 25542
rect 5196 25540 5220 25542
rect 5276 25540 5300 25542
rect 5356 25540 5380 25542
rect 5436 25540 5442 25542
rect 5134 25531 5442 25540
rect 5794 25052 6102 25061
rect 5794 25050 5800 25052
rect 5856 25050 5880 25052
rect 5936 25050 5960 25052
rect 6016 25050 6040 25052
rect 6096 25050 6102 25052
rect 5856 24998 5858 25050
rect 6038 24998 6040 25050
rect 5794 24996 5800 24998
rect 5856 24996 5880 24998
rect 5936 24996 5960 24998
rect 6016 24996 6040 24998
rect 6096 24996 6102 24998
rect 5794 24987 6102 24996
rect 5134 24508 5442 24517
rect 5134 24506 5140 24508
rect 5196 24506 5220 24508
rect 5276 24506 5300 24508
rect 5356 24506 5380 24508
rect 5436 24506 5442 24508
rect 5196 24454 5198 24506
rect 5378 24454 5380 24506
rect 5134 24452 5140 24454
rect 5196 24452 5220 24454
rect 5276 24452 5300 24454
rect 5356 24452 5380 24454
rect 5436 24452 5442 24454
rect 5134 24443 5442 24452
rect 3514 24168 3570 24177
rect 3514 24103 3570 24112
rect 5794 23964 6102 23973
rect 5794 23962 5800 23964
rect 5856 23962 5880 23964
rect 5936 23962 5960 23964
rect 6016 23962 6040 23964
rect 6096 23962 6102 23964
rect 5856 23910 5858 23962
rect 6038 23910 6040 23962
rect 5794 23908 5800 23910
rect 5856 23908 5880 23910
rect 5936 23908 5960 23910
rect 6016 23908 6040 23910
rect 6096 23908 6102 23910
rect 5794 23899 6102 23908
rect 5134 23420 5442 23429
rect 5134 23418 5140 23420
rect 5196 23418 5220 23420
rect 5276 23418 5300 23420
rect 5356 23418 5380 23420
rect 5436 23418 5442 23420
rect 5196 23366 5198 23418
rect 5378 23366 5380 23418
rect 5134 23364 5140 23366
rect 5196 23364 5220 23366
rect 5276 23364 5300 23366
rect 5356 23364 5380 23366
rect 5436 23364 5442 23366
rect 5134 23355 5442 23364
rect 5794 22876 6102 22885
rect 5794 22874 5800 22876
rect 5856 22874 5880 22876
rect 5936 22874 5960 22876
rect 6016 22874 6040 22876
rect 6096 22874 6102 22876
rect 5856 22822 5858 22874
rect 6038 22822 6040 22874
rect 5794 22820 5800 22822
rect 5856 22820 5880 22822
rect 5936 22820 5960 22822
rect 6016 22820 6040 22822
rect 6096 22820 6102 22822
rect 5794 22811 6102 22820
rect 5134 22332 5442 22341
rect 5134 22330 5140 22332
rect 5196 22330 5220 22332
rect 5276 22330 5300 22332
rect 5356 22330 5380 22332
rect 5436 22330 5442 22332
rect 5196 22278 5198 22330
rect 5378 22278 5380 22330
rect 5134 22276 5140 22278
rect 5196 22276 5220 22278
rect 5276 22276 5300 22278
rect 5356 22276 5380 22278
rect 5436 22276 5442 22278
rect 5134 22267 5442 22276
rect 5794 21788 6102 21797
rect 5794 21786 5800 21788
rect 5856 21786 5880 21788
rect 5936 21786 5960 21788
rect 6016 21786 6040 21788
rect 6096 21786 6102 21788
rect 5856 21734 5858 21786
rect 6038 21734 6040 21786
rect 5794 21732 5800 21734
rect 5856 21732 5880 21734
rect 5936 21732 5960 21734
rect 6016 21732 6040 21734
rect 6096 21732 6102 21734
rect 5794 21723 6102 21732
rect 5134 21244 5442 21253
rect 5134 21242 5140 21244
rect 5196 21242 5220 21244
rect 5276 21242 5300 21244
rect 5356 21242 5380 21244
rect 5436 21242 5442 21244
rect 5196 21190 5198 21242
rect 5378 21190 5380 21242
rect 5134 21188 5140 21190
rect 5196 21188 5220 21190
rect 5276 21188 5300 21190
rect 5356 21188 5380 21190
rect 5436 21188 5442 21190
rect 5134 21179 5442 21188
rect 5794 20700 6102 20709
rect 5794 20698 5800 20700
rect 5856 20698 5880 20700
rect 5936 20698 5960 20700
rect 6016 20698 6040 20700
rect 6096 20698 6102 20700
rect 5856 20646 5858 20698
rect 6038 20646 6040 20698
rect 5794 20644 5800 20646
rect 5856 20644 5880 20646
rect 5936 20644 5960 20646
rect 6016 20644 6040 20646
rect 6096 20644 6102 20646
rect 5794 20635 6102 20644
rect 5134 20156 5442 20165
rect 5134 20154 5140 20156
rect 5196 20154 5220 20156
rect 5276 20154 5300 20156
rect 5356 20154 5380 20156
rect 5436 20154 5442 20156
rect 5196 20102 5198 20154
rect 5378 20102 5380 20154
rect 5134 20100 5140 20102
rect 5196 20100 5220 20102
rect 5276 20100 5300 20102
rect 5356 20100 5380 20102
rect 5436 20100 5442 20102
rect 5134 20091 5442 20100
rect 5794 19612 6102 19621
rect 5794 19610 5800 19612
rect 5856 19610 5880 19612
rect 5936 19610 5960 19612
rect 6016 19610 6040 19612
rect 6096 19610 6102 19612
rect 5856 19558 5858 19610
rect 6038 19558 6040 19610
rect 5794 19556 5800 19558
rect 5856 19556 5880 19558
rect 5936 19556 5960 19558
rect 6016 19556 6040 19558
rect 6096 19556 6102 19558
rect 5794 19547 6102 19556
rect 5134 19068 5442 19077
rect 5134 19066 5140 19068
rect 5196 19066 5220 19068
rect 5276 19066 5300 19068
rect 5356 19066 5380 19068
rect 5436 19066 5442 19068
rect 5196 19014 5198 19066
rect 5378 19014 5380 19066
rect 5134 19012 5140 19014
rect 5196 19012 5220 19014
rect 5276 19012 5300 19014
rect 5356 19012 5380 19014
rect 5436 19012 5442 19014
rect 5134 19003 5442 19012
rect 5794 18524 6102 18533
rect 5794 18522 5800 18524
rect 5856 18522 5880 18524
rect 5936 18522 5960 18524
rect 6016 18522 6040 18524
rect 6096 18522 6102 18524
rect 5856 18470 5858 18522
rect 6038 18470 6040 18522
rect 5794 18468 5800 18470
rect 5856 18468 5880 18470
rect 5936 18468 5960 18470
rect 6016 18468 6040 18470
rect 6096 18468 6102 18470
rect 5794 18459 6102 18468
rect 5134 17980 5442 17989
rect 5134 17978 5140 17980
rect 5196 17978 5220 17980
rect 5276 17978 5300 17980
rect 5356 17978 5380 17980
rect 5436 17978 5442 17980
rect 5196 17926 5198 17978
rect 5378 17926 5380 17978
rect 5134 17924 5140 17926
rect 5196 17924 5220 17926
rect 5276 17924 5300 17926
rect 5356 17924 5380 17926
rect 5436 17924 5442 17926
rect 5134 17915 5442 17924
rect 5794 17436 6102 17445
rect 5794 17434 5800 17436
rect 5856 17434 5880 17436
rect 5936 17434 5960 17436
rect 6016 17434 6040 17436
rect 6096 17434 6102 17436
rect 5856 17382 5858 17434
rect 6038 17382 6040 17434
rect 5794 17380 5800 17382
rect 5856 17380 5880 17382
rect 5936 17380 5960 17382
rect 6016 17380 6040 17382
rect 6096 17380 6102 17382
rect 5794 17371 6102 17380
rect 5134 16892 5442 16901
rect 5134 16890 5140 16892
rect 5196 16890 5220 16892
rect 5276 16890 5300 16892
rect 5356 16890 5380 16892
rect 5436 16890 5442 16892
rect 5196 16838 5198 16890
rect 5378 16838 5380 16890
rect 5134 16836 5140 16838
rect 5196 16836 5220 16838
rect 5276 16836 5300 16838
rect 5356 16836 5380 16838
rect 5436 16836 5442 16838
rect 5134 16827 5442 16836
rect 5794 16348 6102 16357
rect 5794 16346 5800 16348
rect 5856 16346 5880 16348
rect 5936 16346 5960 16348
rect 6016 16346 6040 16348
rect 6096 16346 6102 16348
rect 5856 16294 5858 16346
rect 6038 16294 6040 16346
rect 5794 16292 5800 16294
rect 5856 16292 5880 16294
rect 5936 16292 5960 16294
rect 6016 16292 6040 16294
rect 6096 16292 6102 16294
rect 5794 16283 6102 16292
rect 5134 15804 5442 15813
rect 5134 15802 5140 15804
rect 5196 15802 5220 15804
rect 5276 15802 5300 15804
rect 5356 15802 5380 15804
rect 5436 15802 5442 15804
rect 5196 15750 5198 15802
rect 5378 15750 5380 15802
rect 5134 15748 5140 15750
rect 5196 15748 5220 15750
rect 5276 15748 5300 15750
rect 5356 15748 5380 15750
rect 5436 15748 5442 15750
rect 5134 15739 5442 15748
rect 5794 15260 6102 15269
rect 5794 15258 5800 15260
rect 5856 15258 5880 15260
rect 5936 15258 5960 15260
rect 6016 15258 6040 15260
rect 6096 15258 6102 15260
rect 5856 15206 5858 15258
rect 6038 15206 6040 15258
rect 5794 15204 5800 15206
rect 5856 15204 5880 15206
rect 5936 15204 5960 15206
rect 6016 15204 6040 15206
rect 6096 15204 6102 15206
rect 5794 15195 6102 15204
rect 5134 14716 5442 14725
rect 5134 14714 5140 14716
rect 5196 14714 5220 14716
rect 5276 14714 5300 14716
rect 5356 14714 5380 14716
rect 5436 14714 5442 14716
rect 5196 14662 5198 14714
rect 5378 14662 5380 14714
rect 5134 14660 5140 14662
rect 5196 14660 5220 14662
rect 5276 14660 5300 14662
rect 5356 14660 5380 14662
rect 5436 14660 5442 14662
rect 5134 14651 5442 14660
rect 5794 14172 6102 14181
rect 5794 14170 5800 14172
rect 5856 14170 5880 14172
rect 5936 14170 5960 14172
rect 6016 14170 6040 14172
rect 6096 14170 6102 14172
rect 5856 14118 5858 14170
rect 6038 14118 6040 14170
rect 5794 14116 5800 14118
rect 5856 14116 5880 14118
rect 5936 14116 5960 14118
rect 6016 14116 6040 14118
rect 6096 14116 6102 14118
rect 5794 14107 6102 14116
rect 5134 13628 5442 13637
rect 5134 13626 5140 13628
rect 5196 13626 5220 13628
rect 5276 13626 5300 13628
rect 5356 13626 5380 13628
rect 5436 13626 5442 13628
rect 5196 13574 5198 13626
rect 5378 13574 5380 13626
rect 5134 13572 5140 13574
rect 5196 13572 5220 13574
rect 5276 13572 5300 13574
rect 5356 13572 5380 13574
rect 5436 13572 5442 13574
rect 5134 13563 5442 13572
rect 5794 13084 6102 13093
rect 5794 13082 5800 13084
rect 5856 13082 5880 13084
rect 5936 13082 5960 13084
rect 6016 13082 6040 13084
rect 6096 13082 6102 13084
rect 5856 13030 5858 13082
rect 6038 13030 6040 13082
rect 5794 13028 5800 13030
rect 5856 13028 5880 13030
rect 5936 13028 5960 13030
rect 6016 13028 6040 13030
rect 6096 13028 6102 13030
rect 5794 13019 6102 13028
rect 5134 12540 5442 12549
rect 5134 12538 5140 12540
rect 5196 12538 5220 12540
rect 5276 12538 5300 12540
rect 5356 12538 5380 12540
rect 5436 12538 5442 12540
rect 5196 12486 5198 12538
rect 5378 12486 5380 12538
rect 5134 12484 5140 12486
rect 5196 12484 5220 12486
rect 5276 12484 5300 12486
rect 5356 12484 5380 12486
rect 5436 12484 5442 12486
rect 5134 12475 5442 12484
rect 5794 11996 6102 12005
rect 5794 11994 5800 11996
rect 5856 11994 5880 11996
rect 5936 11994 5960 11996
rect 6016 11994 6040 11996
rect 6096 11994 6102 11996
rect 5856 11942 5858 11994
rect 6038 11942 6040 11994
rect 5794 11940 5800 11942
rect 5856 11940 5880 11942
rect 5936 11940 5960 11942
rect 6016 11940 6040 11942
rect 6096 11940 6102 11942
rect 5794 11931 6102 11940
rect 5134 11452 5442 11461
rect 5134 11450 5140 11452
rect 5196 11450 5220 11452
rect 5276 11450 5300 11452
rect 5356 11450 5380 11452
rect 5436 11450 5442 11452
rect 5196 11398 5198 11450
rect 5378 11398 5380 11450
rect 5134 11396 5140 11398
rect 5196 11396 5220 11398
rect 5276 11396 5300 11398
rect 5356 11396 5380 11398
rect 5436 11396 5442 11398
rect 5134 11387 5442 11396
rect 5794 10908 6102 10917
rect 5794 10906 5800 10908
rect 5856 10906 5880 10908
rect 5936 10906 5960 10908
rect 6016 10906 6040 10908
rect 6096 10906 6102 10908
rect 5856 10854 5858 10906
rect 6038 10854 6040 10906
rect 5794 10852 5800 10854
rect 5856 10852 5880 10854
rect 5936 10852 5960 10854
rect 6016 10852 6040 10854
rect 6096 10852 6102 10854
rect 5794 10843 6102 10852
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 5134 10364 5442 10373
rect 5134 10362 5140 10364
rect 5196 10362 5220 10364
rect 5276 10362 5300 10364
rect 5356 10362 5380 10364
rect 5436 10362 5442 10364
rect 5196 10310 5198 10362
rect 5378 10310 5380 10362
rect 5134 10308 5140 10310
rect 5196 10308 5220 10310
rect 5276 10308 5300 10310
rect 5356 10308 5380 10310
rect 5436 10308 5442 10310
rect 5134 10299 5442 10308
rect 9034 9888 9090 9897
rect 5794 9820 6102 9829
rect 9034 9823 9090 9832
rect 5794 9818 5800 9820
rect 5856 9818 5880 9820
rect 5936 9818 5960 9820
rect 6016 9818 6040 9820
rect 6096 9818 6102 9820
rect 5856 9766 5858 9818
rect 6038 9766 6040 9818
rect 5794 9764 5800 9766
rect 5856 9764 5880 9766
rect 5936 9764 5960 9766
rect 6016 9764 6040 9766
rect 6096 9764 6102 9766
rect 5794 9755 6102 9764
rect 5134 9276 5442 9285
rect 5134 9274 5140 9276
rect 5196 9274 5220 9276
rect 5276 9274 5300 9276
rect 5356 9274 5380 9276
rect 5436 9274 5442 9276
rect 5196 9222 5198 9274
rect 5378 9222 5380 9274
rect 5134 9220 5140 9222
rect 5196 9220 5220 9222
rect 5276 9220 5300 9222
rect 5356 9220 5380 9222
rect 5436 9220 5442 9222
rect 5134 9211 5442 9220
rect 5794 8732 6102 8741
rect 5794 8730 5800 8732
rect 5856 8730 5880 8732
rect 5936 8730 5960 8732
rect 6016 8730 6040 8732
rect 6096 8730 6102 8732
rect 5856 8678 5858 8730
rect 6038 8678 6040 8730
rect 5794 8676 5800 8678
rect 5856 8676 5880 8678
rect 5936 8676 5960 8678
rect 6016 8676 6040 8678
rect 6096 8676 6102 8678
rect 5794 8667 6102 8676
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3620 2446 3648 5850
rect 3804 2650 3832 6122
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3988 2514 4016 8298
rect 5134 8188 5442 8197
rect 5134 8186 5140 8188
rect 5196 8186 5220 8188
rect 5276 8186 5300 8188
rect 5356 8186 5380 8188
rect 5436 8186 5442 8188
rect 5196 8134 5198 8186
rect 5378 8134 5380 8186
rect 5134 8132 5140 8134
rect 5196 8132 5220 8134
rect 5276 8132 5300 8134
rect 5356 8132 5380 8134
rect 5436 8132 5442 8134
rect 5134 8123 5442 8132
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 5794 7644 6102 7653
rect 5794 7642 5800 7644
rect 5856 7642 5880 7644
rect 5936 7642 5960 7644
rect 6016 7642 6040 7644
rect 6096 7642 6102 7644
rect 5856 7590 5858 7642
rect 6038 7590 6040 7642
rect 5794 7588 5800 7590
rect 5856 7588 5880 7590
rect 5936 7588 5960 7590
rect 6016 7588 6040 7590
rect 6096 7588 6102 7590
rect 5794 7579 6102 7588
rect 5134 7100 5442 7109
rect 5134 7098 5140 7100
rect 5196 7098 5220 7100
rect 5276 7098 5300 7100
rect 5356 7098 5380 7100
rect 5436 7098 5442 7100
rect 5196 7046 5198 7098
rect 5378 7046 5380 7098
rect 5134 7044 5140 7046
rect 5196 7044 5220 7046
rect 5276 7044 5300 7046
rect 5356 7044 5380 7046
rect 5436 7044 5442 7046
rect 5134 7035 5442 7044
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4356 3058 4384 6802
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4540 2650 4568 6870
rect 5794 6556 6102 6565
rect 5794 6554 5800 6556
rect 5856 6554 5880 6556
rect 5936 6554 5960 6556
rect 6016 6554 6040 6556
rect 6096 6554 6102 6556
rect 5856 6502 5858 6554
rect 6038 6502 6040 6554
rect 5794 6500 5800 6502
rect 5856 6500 5880 6502
rect 5936 6500 5960 6502
rect 6016 6500 6040 6502
rect 6096 6500 6102 6502
rect 5794 6491 6102 6500
rect 5134 6012 5442 6021
rect 5134 6010 5140 6012
rect 5196 6010 5220 6012
rect 5276 6010 5300 6012
rect 5356 6010 5380 6012
rect 5436 6010 5442 6012
rect 5196 5958 5198 6010
rect 5378 5958 5380 6010
rect 5134 5956 5140 5958
rect 5196 5956 5220 5958
rect 5276 5956 5300 5958
rect 5356 5956 5380 5958
rect 5436 5956 5442 5958
rect 5134 5947 5442 5956
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4724 2446 4752 5510
rect 5794 5468 6102 5477
rect 5794 5466 5800 5468
rect 5856 5466 5880 5468
rect 5936 5466 5960 5468
rect 6016 5466 6040 5468
rect 6096 5466 6102 5468
rect 5856 5414 5858 5466
rect 6038 5414 6040 5466
rect 5794 5412 5800 5414
rect 5856 5412 5880 5414
rect 5936 5412 5960 5414
rect 6016 5412 6040 5414
rect 6096 5412 6102 5414
rect 5794 5403 6102 5412
rect 5134 4924 5442 4933
rect 5134 4922 5140 4924
rect 5196 4922 5220 4924
rect 5276 4922 5300 4924
rect 5356 4922 5380 4924
rect 5436 4922 5442 4924
rect 5196 4870 5198 4922
rect 5378 4870 5380 4922
rect 5134 4868 5140 4870
rect 5196 4868 5220 4870
rect 5276 4868 5300 4870
rect 5356 4868 5380 4870
rect 5436 4868 5442 4870
rect 5134 4859 5442 4868
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 5794 4380 6102 4389
rect 5794 4378 5800 4380
rect 5856 4378 5880 4380
rect 5936 4378 5960 4380
rect 6016 4378 6040 4380
rect 6096 4378 6102 4380
rect 5856 4326 5858 4378
rect 6038 4326 6040 4378
rect 5794 4324 5800 4326
rect 5856 4324 5880 4326
rect 5936 4324 5960 4326
rect 6016 4324 6040 4326
rect 6096 4324 6102 4326
rect 5794 4315 6102 4324
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4908 3194 4936 3946
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5134 3836 5442 3845
rect 5134 3834 5140 3836
rect 5196 3834 5220 3836
rect 5276 3834 5300 3836
rect 5356 3834 5380 3836
rect 5436 3834 5442 3836
rect 5196 3782 5198 3834
rect 5378 3782 5380 3834
rect 5134 3780 5140 3782
rect 5196 3780 5220 3782
rect 5276 3780 5300 3782
rect 5356 3780 5380 3782
rect 5436 3780 5442 3782
rect 5134 3771 5442 3780
rect 5078 3632 5134 3641
rect 5078 3567 5134 3576
rect 5092 3534 5120 3567
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5552 3058 5580 3878
rect 6012 3738 6040 4082
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5134 2748 5442 2757
rect 5134 2746 5140 2748
rect 5196 2746 5220 2748
rect 5276 2746 5300 2748
rect 5356 2746 5380 2748
rect 5436 2746 5442 2748
rect 5196 2694 5198 2746
rect 5378 2694 5380 2746
rect 5134 2692 5140 2694
rect 5196 2692 5220 2694
rect 5276 2692 5300 2694
rect 5356 2692 5380 2694
rect 5436 2692 5442 2694
rect 5134 2683 5442 2692
rect 5644 2650 5672 3470
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 5630 2408 5686 2417
rect 5630 2343 5632 2352
rect 5684 2343 5686 2352
rect 5632 2314 5684 2320
rect 5736 1902 5764 3674
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 5794 3292 6102 3301
rect 5794 3290 5800 3292
rect 5856 3290 5880 3292
rect 5936 3290 5960 3292
rect 6016 3290 6040 3292
rect 6096 3290 6102 3292
rect 5856 3238 5858 3290
rect 6038 3238 6040 3290
rect 5794 3236 5800 3238
rect 5856 3236 5880 3238
rect 5936 3236 5960 3238
rect 6016 3236 6040 3238
rect 6096 3236 6102 3238
rect 5794 3227 6102 3236
rect 5814 2544 5870 2553
rect 5814 2479 5816 2488
rect 5868 2479 5870 2488
rect 5816 2450 5868 2456
rect 6196 2446 6224 3470
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 5794 2204 6102 2213
rect 5794 2202 5800 2204
rect 5856 2202 5880 2204
rect 5936 2202 5960 2204
rect 6016 2202 6040 2204
rect 6096 2202 6102 2204
rect 5856 2150 5858 2202
rect 6038 2150 6040 2202
rect 5794 2148 5800 2150
rect 5856 2148 5880 2150
rect 5936 2148 5960 2150
rect 6016 2148 6040 2150
rect 6096 2148 6102 2150
rect 5794 2139 6102 2148
rect 6288 2106 6316 3538
rect 6380 2650 6408 4150
rect 6840 3602 6868 4422
rect 6932 4214 6960 7822
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 3126 6776 3334
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 7024 3058 7052 6394
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7392 4282 7420 4558
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7470 3632 7526 3641
rect 7470 3567 7526 3576
rect 7484 3466 7512 3567
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7576 2990 7604 5782
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 3233 7696 3470
rect 7654 3224 7710 3233
rect 7852 3194 7880 5714
rect 7654 3159 7710 3168
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 7668 2446 7696 2790
rect 7944 2514 7972 6054
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 8036 2922 8064 5578
rect 8128 4010 8156 6258
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8220 3534 8248 8434
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8312 3670 8340 5646
rect 8300 3664 8352 3670
rect 8300 3606 8352 3612
rect 8404 3534 8432 6598
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8956 4826 8984 6190
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8390 3088 8446 3097
rect 8300 3052 8352 3058
rect 8390 3023 8392 3032
rect 8300 2994 8352 3000
rect 8444 3023 8446 3032
rect 8392 2994 8444 3000
rect 8024 2916 8076 2922
rect 8024 2858 8076 2864
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 6276 2100 6328 2106
rect 6276 2042 6328 2048
rect 5724 1896 5776 1902
rect 5724 1838 5776 1844
rect 7668 338 7696 2382
rect 8312 1834 8340 2994
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8300 1828 8352 1834
rect 8300 1770 8352 1776
rect 7656 332 7708 338
rect 7656 274 7708 280
rect 8404 202 8432 2382
rect 8588 1698 8616 4014
rect 9048 3058 9076 9823
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 10414 8936 10470 8945
rect 9678 7576 9734 7585
rect 9678 7511 9734 7520
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9140 3194 9168 3538
rect 9416 3194 9444 4422
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9692 3058 9720 7511
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9784 5914 9812 6054
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9876 5846 9904 6054
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9784 4690 9812 5510
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9784 3618 9812 4218
rect 9876 3738 9904 5170
rect 9968 5030 9996 8910
rect 10414 8871 10470 8880
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10138 6216 10194 6225
rect 10138 6151 10194 6160
rect 10152 5914 10180 6151
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10244 5234 10272 7686
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9968 4690 9996 4966
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 9968 4282 9996 4490
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9784 3590 9904 3618
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8864 2582 8892 2926
rect 9784 2650 9812 3470
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8956 1766 8984 2246
rect 9140 2038 9168 2382
rect 9876 2360 9904 3590
rect 9968 2825 9996 3946
rect 9954 2816 10010 2825
rect 9954 2751 10010 2760
rect 10060 2650 10088 4490
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10152 3398 10180 4014
rect 10244 3618 10272 4150
rect 10336 4146 10364 5646
rect 10428 5234 10456 8871
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10428 4078 10456 5034
rect 10520 4468 10548 10474
rect 11808 9178 11836 36586
rect 14568 14521 14596 37198
rect 15028 37194 15056 37318
rect 15108 37256 15160 37262
rect 15108 37198 15160 37204
rect 15016 37188 15068 37194
rect 15016 37130 15068 37136
rect 15120 36922 15148 37198
rect 15108 36916 15160 36922
rect 15108 36858 15160 36864
rect 16960 36854 16988 39200
rect 18800 37262 18828 39200
rect 20640 37262 20668 39200
rect 22480 37346 22508 39200
rect 22480 37318 22600 37346
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 18788 37256 18840 37262
rect 18788 37198 18840 37204
rect 20628 37256 20680 37262
rect 20628 37198 20680 37204
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 18708 36922 18736 37198
rect 18696 36916 18748 36922
rect 18696 36858 18748 36864
rect 16948 36848 17000 36854
rect 16948 36790 17000 36796
rect 18972 36780 19024 36786
rect 18972 36722 19024 36728
rect 18984 29617 19012 36722
rect 18970 29608 19026 29617
rect 18970 29543 19026 29552
rect 21928 18057 21956 37198
rect 22480 36922 22508 37198
rect 22572 37194 22600 37318
rect 22560 37188 22612 37194
rect 22560 37130 22612 37136
rect 22468 36916 22520 36922
rect 22468 36858 22520 36864
rect 24320 36854 24348 39200
rect 26056 37256 26108 37262
rect 26056 37198 26108 37204
rect 26068 36922 26096 37198
rect 26160 37194 26188 39200
rect 28000 37262 28028 39200
rect 27988 37256 28040 37262
rect 27988 37198 28040 37204
rect 29276 37256 29328 37262
rect 29276 37198 29328 37204
rect 26148 37188 26200 37194
rect 26148 37130 26200 37136
rect 26056 36916 26108 36922
rect 26056 36858 26108 36864
rect 24308 36848 24360 36854
rect 24308 36790 24360 36796
rect 25780 36780 25832 36786
rect 25780 36722 25832 36728
rect 25792 33114 25820 36722
rect 25780 33108 25832 33114
rect 25780 33050 25832 33056
rect 27344 33108 27396 33114
rect 27344 33050 27396 33056
rect 26332 32428 26384 32434
rect 26332 32370 26384 32376
rect 26056 29640 26108 29646
rect 26056 29582 26108 29588
rect 25688 26920 25740 26926
rect 25688 26862 25740 26868
rect 25504 24132 25556 24138
rect 25504 24074 25556 24080
rect 21914 18048 21970 18057
rect 21914 17983 21970 17992
rect 14554 14512 14610 14521
rect 14554 14447 14610 14456
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11978 9072 12034 9081
rect 10876 9036 10928 9042
rect 11978 9007 12034 9016
rect 10876 8978 10928 8984
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10612 6390 10640 6734
rect 10704 6458 10732 6734
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10704 5370 10732 5646
rect 10796 5370 10824 7482
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10704 4468 10732 4558
rect 10520 4440 10732 4468
rect 10888 4162 10916 8978
rect 11702 8664 11758 8673
rect 11702 8599 11758 8608
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10796 4134 10916 4162
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10692 3664 10744 3670
rect 10244 3590 10364 3618
rect 10692 3606 10744 3612
rect 10232 3528 10284 3534
rect 10230 3496 10232 3505
rect 10284 3496 10286 3505
rect 10230 3431 10286 3440
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9692 2332 9904 2360
rect 9128 2032 9180 2038
rect 9128 1974 9180 1980
rect 8944 1760 8996 1766
rect 8944 1702 8996 1708
rect 8576 1692 8628 1698
rect 8576 1634 8628 1640
rect 9048 870 9168 898
rect 9048 800 9076 870
rect 8392 196 8444 202
rect 8392 138 8444 144
rect 9034 0 9090 800
rect 9140 134 9168 870
rect 9692 800 9720 2332
rect 9128 128 9180 134
rect 9128 70 9180 76
rect 9678 0 9734 800
rect 10152 270 10180 3334
rect 10336 800 10364 3590
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10612 3074 10640 3130
rect 10520 3058 10640 3074
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10508 3052 10640 3058
rect 10560 3046 10640 3052
rect 10508 2994 10560 3000
rect 10428 2689 10456 2994
rect 10506 2952 10562 2961
rect 10506 2887 10508 2896
rect 10560 2887 10562 2896
rect 10508 2858 10560 2864
rect 10414 2680 10470 2689
rect 10414 2615 10470 2624
rect 10428 2446 10456 2615
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10612 1970 10640 2382
rect 10600 1964 10652 1970
rect 10600 1906 10652 1912
rect 10140 264 10192 270
rect 10140 206 10192 212
rect 10322 0 10378 800
rect 10704 762 10732 3606
rect 10796 2514 10824 4134
rect 10876 4072 10928 4078
rect 10874 4040 10876 4049
rect 10928 4040 10930 4049
rect 10874 3975 10930 3984
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10980 2378 11008 6870
rect 11072 4826 11100 7346
rect 11164 5914 11192 7890
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11348 5710 11376 6666
rect 11624 6458 11652 6734
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11244 4684 11296 4690
rect 11296 4644 11376 4672
rect 11244 4626 11296 4632
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 11072 2514 11100 4490
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 4146 11192 4422
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11256 2582 11284 4218
rect 11348 3369 11376 4644
rect 11440 4486 11468 5646
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11428 3392 11480 3398
rect 11334 3360 11390 3369
rect 11428 3334 11480 3340
rect 11334 3295 11390 3304
rect 11348 3126 11376 3295
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 11440 2990 11468 3334
rect 11532 2990 11560 5646
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11624 4690 11652 5170
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11716 4162 11744 8599
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11808 6186 11836 6734
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11888 6180 11940 6186
rect 11888 6122 11940 6128
rect 11900 5370 11928 6122
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11992 4826 12020 9007
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12162 5672 12218 5681
rect 12162 5607 12218 5616
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11624 4134 11744 4162
rect 11624 4078 11652 4134
rect 11612 4072 11664 4078
rect 11704 4072 11756 4078
rect 11612 4014 11664 4020
rect 11702 4040 11704 4049
rect 11888 4072 11940 4078
rect 11756 4040 11758 4049
rect 11888 4014 11940 4020
rect 11702 3975 11758 3984
rect 11702 3904 11758 3913
rect 11702 3839 11758 3848
rect 11716 3534 11744 3839
rect 11900 3738 11928 4014
rect 11980 4004 12032 4010
rect 12084 3992 12112 5510
rect 12176 4690 12204 5607
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12032 3964 12112 3992
rect 11980 3946 12032 3952
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12176 3194 12204 3402
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11532 2446 11560 2926
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 11808 2310 11836 2450
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 11612 2100 11664 2106
rect 11612 2042 11664 2048
rect 10888 870 11008 898
rect 10888 762 10916 870
rect 10980 800 11008 870
rect 11624 800 11652 2042
rect 11716 1902 11744 2246
rect 11704 1896 11756 1902
rect 11704 1838 11756 1844
rect 12268 800 12296 6190
rect 12360 5234 12388 7142
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12452 5914 12480 6734
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12440 5636 12492 5642
rect 12544 5624 12572 6598
rect 12714 6352 12770 6361
rect 12714 6287 12716 6296
rect 12768 6287 12770 6296
rect 12716 6258 12768 6264
rect 12716 6112 12768 6118
rect 12714 6080 12716 6089
rect 12768 6080 12770 6089
rect 12714 6015 12770 6024
rect 12492 5596 12572 5624
rect 12440 5578 12492 5584
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12452 4758 12480 4966
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12544 2774 12572 5238
rect 12622 4856 12678 4865
rect 12622 4791 12624 4800
rect 12676 4791 12678 4800
rect 12624 4762 12676 4768
rect 12622 4720 12678 4729
rect 12622 4655 12678 4664
rect 12636 4146 12664 4655
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12820 3602 12848 4422
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12728 3369 12756 3402
rect 12714 3360 12770 3369
rect 12714 3295 12770 3304
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12544 2746 12664 2774
rect 12636 2514 12664 2746
rect 12728 2650 12756 2790
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12820 2446 12848 3538
rect 12912 3194 12940 8366
rect 13004 5302 13032 11494
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13542 9752 13598 9761
rect 13542 9687 13598 9696
rect 13450 9344 13506 9353
rect 13450 9279 13506 9288
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 13174 5264 13230 5273
rect 13174 5199 13230 5208
rect 13188 5166 13216 5199
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 12990 3904 13046 3913
rect 12990 3839 13046 3848
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 13004 3058 13032 3839
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 12992 2372 13044 2378
rect 12992 2314 13044 2320
rect 13004 2106 13032 2314
rect 12992 2100 13044 2106
rect 12992 2042 13044 2048
rect 12912 870 13032 898
rect 12912 800 12940 870
rect 10704 734 10916 762
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13004 762 13032 870
rect 13188 762 13216 4694
rect 13280 3942 13308 5510
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13372 3126 13400 6394
rect 13464 4622 13492 9279
rect 13556 4826 13584 9687
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13464 2990 13492 4218
rect 13556 3641 13584 4558
rect 13542 3632 13598 3641
rect 13542 3567 13598 3576
rect 13648 3482 13676 6326
rect 13740 4146 13768 9930
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13832 5710 13860 9318
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13924 5556 13952 8502
rect 14094 5944 14150 5953
rect 14094 5879 14150 5888
rect 14108 5710 14136 5879
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 13832 5528 13952 5556
rect 13832 5166 13860 5528
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13648 3454 13768 3482
rect 13740 3398 13768 3454
rect 13728 3392 13780 3398
rect 13634 3360 13690 3369
rect 13728 3334 13780 3340
rect 13634 3295 13690 3304
rect 13648 3126 13676 3295
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 13832 2990 13860 3946
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13820 2984 13872 2990
rect 13924 2961 13952 5102
rect 14094 4992 14150 5001
rect 14094 4927 14150 4936
rect 14108 3670 14136 4927
rect 14200 4758 14228 12650
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14292 7002 14320 7346
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14292 4554 14320 6598
rect 14384 4690 14412 6598
rect 14476 5914 14504 7346
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 6322 14596 7142
rect 14648 6928 14700 6934
rect 14648 6870 14700 6876
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14660 6118 14688 6870
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14752 5930 14780 10406
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14660 5902 14780 5930
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14280 4548 14332 4554
rect 14280 4490 14332 4496
rect 14476 4282 14504 4626
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14476 3942 14504 4218
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14278 3768 14334 3777
rect 14278 3703 14334 3712
rect 14096 3664 14148 3670
rect 14002 3632 14058 3641
rect 14096 3606 14148 3612
rect 14292 3602 14320 3703
rect 14002 3567 14058 3576
rect 14280 3596 14332 3602
rect 14016 3534 14044 3567
rect 14280 3538 14332 3544
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 13820 2926 13872 2932
rect 13910 2952 13966 2961
rect 13910 2887 13966 2896
rect 14016 2774 14044 3470
rect 14568 2854 14596 4966
rect 14660 4146 14688 5902
rect 14740 5636 14792 5642
rect 14740 5578 14792 5584
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14648 4004 14700 4010
rect 14648 3946 14700 3952
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 13924 2746 14044 2774
rect 13924 2582 13952 2746
rect 13912 2576 13964 2582
rect 13912 2518 13964 2524
rect 14660 2446 14688 3946
rect 14752 2774 14780 5578
rect 14844 4146 14872 7686
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14752 2746 14872 2774
rect 14844 2514 14872 2746
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 13360 1964 13412 1970
rect 13360 1906 13412 1912
rect 13372 1698 13400 1906
rect 13360 1692 13412 1698
rect 13360 1634 13412 1640
rect 13556 800 13584 2314
rect 14936 1358 14964 6734
rect 15028 5370 15056 7142
rect 15120 5914 15148 8570
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15212 6254 15240 7210
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15106 5672 15162 5681
rect 15290 5672 15346 5681
rect 15162 5630 15240 5658
rect 15106 5607 15162 5616
rect 15212 5574 15240 5630
rect 15290 5607 15292 5616
rect 15344 5607 15346 5616
rect 15292 5578 15344 5584
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15198 5400 15254 5409
rect 15016 5364 15068 5370
rect 15198 5335 15200 5344
rect 15016 5306 15068 5312
rect 15252 5335 15254 5344
rect 15200 5306 15252 5312
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 15028 4457 15056 5170
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15014 4448 15070 4457
rect 15014 4383 15070 4392
rect 15028 4146 15056 4383
rect 15120 4282 15148 4558
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 15106 4176 15162 4185
rect 15016 4140 15068 4146
rect 15106 4111 15162 4120
rect 15016 4082 15068 4088
rect 15120 4078 15148 4111
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15304 3534 15332 5102
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15304 2854 15332 3470
rect 15396 3194 15424 7822
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15488 7206 15516 7346
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15488 3602 15516 6666
rect 15580 6361 15608 9590
rect 15658 9480 15714 9489
rect 15658 9415 15714 9424
rect 15672 6905 15700 9415
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15750 8392 15806 8401
rect 15750 8327 15806 8336
rect 15658 6896 15714 6905
rect 15658 6831 15714 6840
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15672 6458 15700 6734
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15566 6352 15622 6361
rect 15566 6287 15622 6296
rect 15580 5930 15608 6287
rect 15580 5902 15700 5930
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15474 3224 15530 3233
rect 15384 3188 15436 3194
rect 15474 3159 15530 3168
rect 15384 3130 15436 3136
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15212 1630 15240 2246
rect 15200 1624 15252 1630
rect 15200 1566 15252 1572
rect 14924 1352 14976 1358
rect 14924 1294 14976 1300
rect 15488 800 15516 3159
rect 15580 2990 15608 5782
rect 15672 4622 15700 5902
rect 15764 5166 15792 8327
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15856 7002 15884 7142
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15842 6896 15898 6905
rect 15842 6831 15898 6840
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15856 4622 15884 6831
rect 15948 5370 15976 9114
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 16040 5778 16068 7142
rect 16132 6458 16160 8434
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16316 7546 16344 7822
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16118 6352 16174 6361
rect 16118 6287 16174 6296
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 16132 4486 16160 6287
rect 16224 5302 16252 7142
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16316 5817 16344 6802
rect 16408 6322 16436 8298
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16500 6934 16528 7414
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16394 6080 16450 6089
rect 16394 6015 16450 6024
rect 16302 5808 16358 5817
rect 16302 5743 16304 5752
rect 16356 5743 16358 5752
rect 16304 5714 16356 5720
rect 16408 5658 16436 6015
rect 16500 5846 16528 6734
rect 16592 6254 16620 11154
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16684 6458 16712 10542
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 16316 5630 16436 5658
rect 16580 5636 16632 5642
rect 16316 5574 16344 5630
rect 16580 5578 16632 5584
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16316 4486 16344 5102
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16408 4146 16436 5510
rect 16592 4826 16620 5578
rect 16868 5234 16896 10134
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16684 4282 16712 4422
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16776 4214 16804 5102
rect 17038 4856 17094 4865
rect 17038 4791 17040 4800
rect 17092 4791 17094 4800
rect 17040 4762 17092 4768
rect 16854 4584 16910 4593
rect 16854 4519 16910 4528
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16592 3738 16620 4082
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15658 3360 15714 3369
rect 15658 3295 15714 3304
rect 15672 3126 15700 3295
rect 15660 3120 15712 3126
rect 15660 3062 15712 3068
rect 15568 2984 15620 2990
rect 15764 2972 15792 3538
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15948 3369 15976 3402
rect 16212 3392 16264 3398
rect 15934 3360 15990 3369
rect 16212 3334 16264 3340
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 15934 3295 15990 3304
rect 15568 2926 15620 2932
rect 15672 2944 15792 2972
rect 15580 2310 15608 2926
rect 15672 2428 15700 2944
rect 16224 2774 16252 3334
rect 16224 2746 16344 2774
rect 16028 2576 16080 2582
rect 16028 2518 16080 2524
rect 15752 2440 15804 2446
rect 15672 2400 15752 2428
rect 16040 2428 16068 2518
rect 15804 2400 16068 2428
rect 15752 2382 15804 2388
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 16316 1902 16344 2746
rect 16408 2310 16436 3334
rect 16500 3058 16528 3606
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16408 2038 16436 2246
rect 16396 2032 16448 2038
rect 16396 1974 16448 1980
rect 16304 1896 16356 1902
rect 16304 1838 16356 1844
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 16132 800 16160 1294
rect 16776 800 16804 3674
rect 16868 3466 16896 4519
rect 16946 3904 17002 3913
rect 16946 3839 17002 3848
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16868 3233 16896 3402
rect 16854 3224 16910 3233
rect 16854 3159 16910 3168
rect 16960 2990 16988 3839
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16868 2650 16896 2790
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 16960 2378 16988 2926
rect 17144 2650 17172 8366
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 4146 17264 6598
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17328 3602 17356 8298
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 17420 1329 17448 7822
rect 17512 2990 17540 10678
rect 17604 9178 17632 12582
rect 24674 12200 24730 12209
rect 24674 12135 24730 12144
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17592 6180 17644 6186
rect 17592 6122 17644 6128
rect 17604 5234 17632 6122
rect 17696 5710 17724 9114
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17788 6866 17816 8978
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17972 8090 18000 8910
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 18064 6866 18092 8842
rect 18156 8634 18184 8842
rect 18248 8809 18276 10950
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18420 8832 18472 8838
rect 18234 8800 18290 8809
rect 18420 8774 18472 8780
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18234 8735 18290 8744
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17868 6792 17920 6798
rect 17920 6740 18092 6746
rect 17868 6734 18092 6740
rect 17880 6718 18092 6734
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17788 5630 18000 5658
rect 17682 5264 17738 5273
rect 17592 5228 17644 5234
rect 17682 5199 17684 5208
rect 17592 5170 17644 5176
rect 17736 5199 17738 5208
rect 17684 5170 17736 5176
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17604 4214 17632 4966
rect 17682 4856 17738 4865
rect 17682 4791 17738 4800
rect 17696 4758 17724 4791
rect 17684 4752 17736 4758
rect 17684 4694 17736 4700
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 17788 3126 17816 5630
rect 17972 5574 18000 5630
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17880 2446 17908 5510
rect 17960 3460 18012 3466
rect 18064 3448 18092 6718
rect 18156 6662 18184 8366
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18156 5370 18184 6190
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18156 4010 18184 5170
rect 18248 5166 18276 7686
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18156 3534 18184 3946
rect 18248 3534 18276 4014
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18012 3420 18092 3448
rect 17960 3402 18012 3408
rect 18156 3194 18184 3470
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 17958 2816 18014 2825
rect 18340 2774 18368 7890
rect 18432 6458 18460 8774
rect 18616 8537 18644 8774
rect 18602 8528 18658 8537
rect 18602 8463 18658 8472
rect 18708 8401 18736 9522
rect 18892 8430 18920 9590
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 18880 8424 18932 8430
rect 18694 8392 18750 8401
rect 18880 8366 18932 8372
rect 18694 8327 18750 8336
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18604 7812 18656 7818
rect 18604 7754 18656 7760
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 17958 2751 18014 2760
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17406 1320 17462 1329
rect 17406 1255 17462 1264
rect 17972 1034 18000 2751
rect 18156 2746 18368 2774
rect 18432 2774 18460 5850
rect 18524 5302 18552 6598
rect 18616 6254 18644 7754
rect 18800 7206 18828 7822
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18696 6112 18748 6118
rect 18602 6080 18658 6089
rect 18696 6054 18748 6060
rect 18602 6015 18658 6024
rect 18616 5914 18644 6015
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18708 5710 18736 6054
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 18602 5536 18658 5545
rect 18602 5471 18658 5480
rect 18512 5296 18564 5302
rect 18512 5238 18564 5244
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18524 5030 18552 5102
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18512 4752 18564 4758
rect 18512 4694 18564 4700
rect 18524 4321 18552 4694
rect 18616 4622 18644 5471
rect 18694 5128 18750 5137
rect 18694 5063 18750 5072
rect 18708 4622 18736 5063
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18510 4312 18566 4321
rect 18510 4247 18566 4256
rect 18800 4078 18828 6938
rect 18984 5370 19012 9046
rect 19076 6798 19104 9454
rect 19168 8090 19196 9522
rect 19260 8634 19288 10610
rect 19444 10062 19472 11630
rect 21916 11620 21968 11626
rect 21916 11562 21968 11568
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 19982 10568 20038 10577
rect 19982 10503 20038 10512
rect 19996 10266 20024 10503
rect 19892 10260 19944 10266
rect 19892 10202 19944 10208
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19904 10146 19932 10202
rect 20088 10146 20116 10746
rect 19904 10118 20116 10146
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19340 9648 19392 9654
rect 19444 9620 19472 9998
rect 19720 9674 19748 9998
rect 19720 9646 19840 9674
rect 19340 9590 19392 9596
rect 19432 9614 19484 9620
rect 19352 9081 19380 9590
rect 19432 9556 19484 9562
rect 19616 9614 19668 9620
rect 19616 9556 19668 9562
rect 19338 9072 19394 9081
rect 19338 9007 19394 9016
rect 19444 8634 19472 9556
rect 19628 9081 19656 9556
rect 19614 9072 19670 9081
rect 19614 9007 19670 9016
rect 19616 8900 19668 8906
rect 19616 8842 19668 8848
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19260 6474 19288 8298
rect 19352 6798 19380 8366
rect 19432 8356 19484 8362
rect 19432 8298 19484 8304
rect 19444 7954 19472 8298
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19432 7336 19484 7342
rect 19430 7304 19432 7313
rect 19484 7304 19486 7313
rect 19430 7239 19486 7248
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19076 6446 19288 6474
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 19076 4264 19104 6446
rect 19246 6352 19302 6361
rect 19352 6322 19380 6598
rect 19246 6287 19302 6296
rect 19340 6316 19392 6322
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19168 5778 19196 6190
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19168 4593 19196 5306
rect 19260 4758 19288 6287
rect 19340 6258 19392 6264
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19338 6216 19394 6225
rect 19338 6151 19394 6160
rect 19352 5778 19380 6151
rect 19444 5914 19472 6258
rect 19536 5914 19564 8774
rect 19628 6798 19656 8842
rect 19812 8378 19840 9646
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19904 8673 19932 8910
rect 19890 8664 19946 8673
rect 19890 8599 19946 8608
rect 19892 8560 19944 8566
rect 19996 8537 20024 9522
rect 19892 8502 19944 8508
rect 19982 8528 20038 8537
rect 19720 8350 19840 8378
rect 19720 7478 19748 8350
rect 19800 8288 19852 8294
rect 19800 8230 19852 8236
rect 19812 8090 19840 8230
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19708 7472 19760 7478
rect 19708 7414 19760 7420
rect 19616 6792 19668 6798
rect 19614 6760 19616 6769
rect 19668 6760 19670 6769
rect 19614 6695 19670 6704
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19430 5808 19486 5817
rect 19340 5772 19392 5778
rect 19430 5743 19486 5752
rect 19340 5714 19392 5720
rect 19444 5574 19472 5743
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19536 5409 19564 5850
rect 19522 5400 19578 5409
rect 19522 5335 19578 5344
rect 19430 4856 19486 4865
rect 19430 4791 19486 4800
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 19444 4622 19472 4791
rect 19432 4616 19484 4622
rect 19154 4584 19210 4593
rect 19432 4558 19484 4564
rect 19154 4519 19210 4528
rect 19536 4486 19564 5335
rect 19628 4758 19656 6695
rect 19720 6066 19748 7414
rect 19812 6254 19840 7686
rect 19904 7002 19932 8502
rect 19982 8463 20038 8472
rect 20088 8072 20116 10118
rect 20272 8974 20300 11018
rect 20260 8968 20312 8974
rect 20180 8928 20260 8956
rect 20180 8838 20208 8928
rect 20260 8910 20312 8916
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 19996 8044 20116 8072
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 19720 6038 19932 6066
rect 19616 4752 19668 4758
rect 19616 4694 19668 4700
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19706 4584 19762 4593
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19076 4236 19196 4264
rect 19062 4176 19118 4185
rect 19168 4146 19196 4236
rect 19340 4208 19392 4214
rect 19338 4176 19340 4185
rect 19524 4208 19576 4214
rect 19392 4176 19394 4185
rect 19062 4111 19118 4120
rect 19156 4140 19208 4146
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 3126 18644 3334
rect 19076 3126 19104 4111
rect 19628 4185 19656 4558
rect 19706 4519 19762 4528
rect 19524 4150 19576 4156
rect 19614 4176 19670 4185
rect 19338 4111 19394 4120
rect 19156 4082 19208 4088
rect 19536 4060 19564 4150
rect 19614 4111 19670 4120
rect 19720 4060 19748 4519
rect 19904 4282 19932 6038
rect 19996 4622 20024 8044
rect 20074 7984 20130 7993
rect 20074 7919 20130 7928
rect 20088 5273 20116 7919
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20074 5264 20130 5273
rect 20074 5199 20130 5208
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19984 4480 20036 4486
rect 19982 4448 19984 4457
rect 20036 4448 20038 4457
rect 19982 4383 20038 4392
rect 19892 4276 19944 4282
rect 19944 4236 20024 4264
rect 19892 4218 19944 4224
rect 19536 4032 19748 4060
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19444 3670 19472 3878
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 19064 3120 19116 3126
rect 19536 3097 19564 3878
rect 19996 3194 20024 4236
rect 20088 3942 20116 5199
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20076 3664 20128 3670
rect 20076 3606 20128 3612
rect 20088 3398 20116 3606
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 20180 3194 20208 6734
rect 20272 6254 20300 8774
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 20272 6118 20300 6190
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20364 5574 20392 11290
rect 21928 11150 21956 11562
rect 22100 11280 22152 11286
rect 22100 11222 22152 11228
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20732 10674 20760 10746
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20824 10130 20852 11086
rect 21638 10976 21694 10985
rect 21638 10911 21694 10920
rect 21652 10742 21680 10911
rect 21640 10736 21692 10742
rect 21640 10678 21692 10684
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20442 8936 20498 8945
rect 20442 8871 20444 8880
rect 20496 8871 20498 8880
rect 20444 8842 20496 8848
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20456 5778 20484 8366
rect 20548 7002 20576 9862
rect 20824 8906 20852 10066
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20732 7410 20760 8774
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20536 6724 20588 6730
rect 20536 6666 20588 6672
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20350 5264 20406 5273
rect 20350 5199 20352 5208
rect 20404 5199 20406 5208
rect 20352 5170 20404 5176
rect 20456 5098 20484 5714
rect 20548 5370 20576 6666
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20444 5092 20496 5098
rect 20444 5034 20496 5040
rect 20444 4752 20496 4758
rect 20444 4694 20496 4700
rect 20260 4548 20312 4554
rect 20260 4490 20312 4496
rect 20272 4162 20300 4490
rect 20456 4214 20484 4694
rect 20640 4214 20668 7278
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20732 6905 20760 7142
rect 20718 6896 20774 6905
rect 20718 6831 20774 6840
rect 20732 5794 20760 6831
rect 20824 6458 20852 8366
rect 20916 8265 20944 9998
rect 21088 9988 21140 9994
rect 21088 9930 21140 9936
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20902 8256 20958 8265
rect 20902 8191 20958 8200
rect 20916 7041 20944 8191
rect 20902 7032 20958 7041
rect 20902 6967 20958 6976
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20732 5766 20852 5794
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20444 4208 20496 4214
rect 20272 4134 20392 4162
rect 20628 4208 20680 4214
rect 20444 4150 20496 4156
rect 20534 4176 20590 4185
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 19904 3097 19932 3130
rect 19064 3062 19116 3068
rect 19522 3088 19578 3097
rect 19522 3023 19578 3032
rect 19890 3088 19946 3097
rect 19890 3023 19946 3032
rect 18432 2746 18644 2774
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18064 1834 18092 2246
rect 18052 1828 18104 1834
rect 18052 1770 18104 1776
rect 18156 1766 18184 2746
rect 18144 1760 18196 1766
rect 18144 1702 18196 1708
rect 18616 1193 18644 2746
rect 20272 2650 20300 4014
rect 20364 3618 20392 4134
rect 20628 4150 20680 4156
rect 20534 4111 20590 4120
rect 20364 3590 20484 3618
rect 20456 3534 20484 3590
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 19338 2544 19394 2553
rect 19338 2479 19340 2488
rect 19392 2479 19394 2488
rect 19340 2450 19392 2456
rect 20364 2446 20392 3470
rect 20548 2854 20576 4111
rect 20732 4026 20760 5646
rect 20824 5234 20852 5766
rect 20904 5704 20956 5710
rect 20904 5646 20956 5652
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20916 4729 20944 5646
rect 21008 5302 21036 9318
rect 21100 8514 21128 9930
rect 21284 9081 21312 10610
rect 22112 10554 22140 11222
rect 22204 11082 22232 11766
rect 22466 11248 22522 11257
rect 22466 11183 22522 11192
rect 22480 11150 22508 11183
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22192 11076 22244 11082
rect 22192 11018 22244 11024
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22112 10526 22232 10554
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21376 10033 21404 10406
rect 21560 10305 21588 10406
rect 21546 10296 21602 10305
rect 21456 10260 21508 10266
rect 21546 10231 21602 10240
rect 21456 10202 21508 10208
rect 21468 10130 21496 10202
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21824 10056 21876 10062
rect 21362 10024 21418 10033
rect 21824 9998 21876 10004
rect 21362 9959 21418 9968
rect 21364 9920 21416 9926
rect 21362 9888 21364 9897
rect 21416 9888 21418 9897
rect 21362 9823 21418 9832
rect 21836 9518 21864 9998
rect 22008 9988 22060 9994
rect 22008 9930 22060 9936
rect 22020 9586 22048 9930
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21732 9444 21784 9450
rect 21732 9386 21784 9392
rect 21270 9072 21326 9081
rect 21270 9007 21326 9016
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21456 8832 21508 8838
rect 21456 8774 21508 8780
rect 21100 8486 21404 8514
rect 21178 8392 21234 8401
rect 21088 8356 21140 8362
rect 21178 8327 21180 8336
rect 21088 8298 21140 8304
rect 21232 8327 21234 8336
rect 21180 8298 21232 8304
rect 21100 6458 21128 8298
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 20996 5296 21048 5302
rect 20996 5238 21048 5244
rect 20902 4720 20958 4729
rect 20902 4655 20958 4664
rect 21100 4214 21128 6054
rect 21192 5914 21220 7346
rect 21376 6118 21404 8486
rect 21468 7585 21496 8774
rect 21454 7576 21510 7585
rect 21454 7511 21510 7520
rect 21560 7410 21588 8842
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21652 7954 21680 8434
rect 21744 7954 21772 9386
rect 21836 7970 21864 9454
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 21928 8566 21956 9046
rect 22112 9042 22140 9862
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 21916 8560 21968 8566
rect 21916 8502 21968 8508
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 21916 8424 21968 8430
rect 21916 8366 21968 8372
rect 21928 8090 21956 8366
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21732 7948 21784 7954
rect 21836 7942 21956 7970
rect 21732 7890 21784 7896
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21730 7576 21786 7585
rect 21730 7511 21786 7520
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21468 6118 21496 7346
rect 21652 7290 21680 7346
rect 21744 7342 21772 7511
rect 21836 7478 21864 7686
rect 21824 7472 21876 7478
rect 21824 7414 21876 7420
rect 21560 7262 21680 7290
rect 21732 7336 21784 7342
rect 21732 7278 21784 7284
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21456 6112 21508 6118
rect 21456 6054 21508 6060
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 21284 5642 21312 6054
rect 21362 5808 21418 5817
rect 21362 5743 21418 5752
rect 21272 5636 21324 5642
rect 21272 5578 21324 5584
rect 21376 5574 21404 5743
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21178 4856 21234 4865
rect 21178 4791 21234 4800
rect 21192 4622 21220 4791
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 21088 4208 21140 4214
rect 21088 4150 21140 4156
rect 20732 3998 21036 4026
rect 20732 3942 20760 3998
rect 21008 3942 21036 3998
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 20352 2440 20404 2446
rect 20352 2382 20404 2388
rect 20180 1834 20208 2382
rect 20352 2304 20404 2310
rect 20352 2246 20404 2252
rect 20628 2304 20680 2310
rect 20732 2281 20760 2450
rect 20628 2246 20680 2252
rect 20718 2272 20774 2281
rect 20168 1828 20220 1834
rect 20168 1770 20220 1776
rect 20364 1630 20392 2246
rect 20640 2106 20668 2246
rect 20718 2207 20774 2216
rect 20628 2100 20680 2106
rect 20628 2042 20680 2048
rect 20352 1624 20404 1630
rect 20352 1566 20404 1572
rect 20824 1465 20852 3538
rect 20916 3505 20944 3878
rect 20902 3496 20958 3505
rect 20902 3431 20958 3440
rect 21100 2854 21128 4150
rect 21376 3913 21404 5510
rect 21454 5400 21510 5409
rect 21560 5370 21588 7262
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 21836 6934 21864 7142
rect 21824 6928 21876 6934
rect 21824 6870 21876 6876
rect 21822 6624 21878 6633
rect 21822 6559 21878 6568
rect 21640 6384 21692 6390
rect 21692 6344 21772 6372
rect 21640 6326 21692 6332
rect 21640 6112 21692 6118
rect 21640 6054 21692 6060
rect 21652 5692 21680 6054
rect 21744 5846 21772 6344
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 21836 5778 21864 6559
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21652 5664 21772 5692
rect 21744 5370 21772 5664
rect 21454 5335 21510 5344
rect 21548 5364 21600 5370
rect 21468 5234 21496 5335
rect 21548 5306 21600 5312
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 21836 5250 21864 5306
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 21652 5222 21864 5250
rect 21652 4060 21680 5222
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21560 4049 21680 4060
rect 21546 4040 21680 4049
rect 21602 4032 21680 4040
rect 21744 3992 21772 5102
rect 21824 5092 21876 5098
rect 21824 5034 21876 5040
rect 21836 4593 21864 5034
rect 21822 4584 21878 4593
rect 21822 4519 21878 4528
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21546 3975 21602 3984
rect 21652 3964 21772 3992
rect 21362 3904 21418 3913
rect 21362 3839 21418 3848
rect 21456 3664 21508 3670
rect 21456 3606 21508 3612
rect 21468 2922 21496 3606
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 21548 2440 21600 2446
rect 21548 2382 21600 2388
rect 21560 1737 21588 2382
rect 21546 1728 21602 1737
rect 21546 1663 21602 1672
rect 19982 1456 20038 1465
rect 19982 1391 20038 1400
rect 20810 1456 20866 1465
rect 20810 1391 20866 1400
rect 19338 1320 19394 1329
rect 19338 1255 19394 1264
rect 18602 1184 18658 1193
rect 18602 1119 18658 1128
rect 17972 1006 18092 1034
rect 18064 800 18092 1006
rect 18616 870 18736 898
rect 13004 734 13216 762
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18616 338 18644 870
rect 18708 800 18736 870
rect 19352 800 19380 1255
rect 19996 800 20024 1391
rect 21192 870 21312 898
rect 18604 332 18656 338
rect 18604 274 18656 280
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21192 270 21220 870
rect 21284 800 21312 870
rect 21180 264 21232 270
rect 21180 206 21232 212
rect 21270 0 21326 800
rect 21652 270 21680 3964
rect 21836 3398 21864 4014
rect 21824 3392 21876 3398
rect 21824 3334 21876 3340
rect 21732 3120 21784 3126
rect 21730 3088 21732 3097
rect 21784 3088 21786 3097
rect 21730 3023 21786 3032
rect 21836 2774 21864 3334
rect 21744 2746 21864 2774
rect 21744 338 21772 2746
rect 21928 800 21956 7942
rect 22020 7426 22048 8502
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 22112 7528 22140 8434
rect 22204 8090 22232 10526
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22296 7546 22324 10610
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22388 8498 22416 9862
rect 22572 9654 22600 11086
rect 22744 10804 22796 10810
rect 22744 10746 22796 10752
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 22756 10674 22784 10746
rect 22836 10736 22888 10742
rect 22836 10678 22888 10684
rect 22744 10668 22796 10674
rect 22744 10610 22796 10616
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22664 10130 22692 10406
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22756 10062 22784 10406
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22848 9586 22876 10678
rect 22928 10056 22980 10062
rect 22928 9998 22980 10004
rect 22940 9625 22968 9998
rect 22926 9616 22982 9625
rect 22836 9580 22888 9586
rect 22756 9540 22836 9568
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22388 7818 22416 8230
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22376 7812 22428 7818
rect 22376 7754 22428 7760
rect 22284 7540 22336 7546
rect 22112 7500 22232 7528
rect 22020 7398 22140 7426
rect 22008 7336 22060 7342
rect 22006 7304 22008 7313
rect 22060 7304 22062 7313
rect 22006 7239 22062 7248
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22020 6497 22048 7142
rect 22112 6730 22140 7398
rect 22204 7206 22232 7500
rect 22284 7482 22336 7488
rect 22374 7440 22430 7449
rect 22374 7375 22430 7384
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22388 6905 22416 7375
rect 22374 6896 22430 6905
rect 22374 6831 22376 6840
rect 22428 6831 22430 6840
rect 22376 6802 22428 6808
rect 22192 6792 22244 6798
rect 22190 6760 22192 6769
rect 22244 6760 22246 6769
rect 22100 6724 22152 6730
rect 22190 6695 22246 6704
rect 22374 6760 22430 6769
rect 22374 6695 22430 6704
rect 22100 6666 22152 6672
rect 22006 6488 22062 6497
rect 22006 6423 22062 6432
rect 22020 6254 22048 6423
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22020 3369 22048 6054
rect 22112 5409 22140 6666
rect 22282 6488 22338 6497
rect 22282 6423 22338 6432
rect 22192 6248 22244 6254
rect 22192 6190 22244 6196
rect 22204 6118 22232 6190
rect 22296 6118 22324 6423
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 22296 5574 22324 6054
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22284 5568 22336 5574
rect 22284 5510 22336 5516
rect 22098 5400 22154 5409
rect 22098 5335 22154 5344
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 22112 4622 22140 4762
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22100 4480 22152 4486
rect 22098 4448 22100 4457
rect 22152 4448 22154 4457
rect 22098 4383 22154 4392
rect 22098 4040 22154 4049
rect 22098 3975 22154 3984
rect 22112 3738 22140 3975
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 22006 3360 22062 3369
rect 22006 3295 22062 3304
rect 22020 3126 22048 3295
rect 22112 3126 22140 3402
rect 22008 3120 22060 3126
rect 22008 3062 22060 3068
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 22204 2514 22232 5510
rect 22282 5400 22338 5409
rect 22282 5335 22338 5344
rect 22296 5302 22324 5335
rect 22284 5296 22336 5302
rect 22284 5238 22336 5244
rect 22284 4616 22336 4622
rect 22282 4584 22284 4593
rect 22336 4584 22338 4593
rect 22282 4519 22338 4528
rect 22282 3224 22338 3233
rect 22282 3159 22338 3168
rect 22296 3058 22324 3159
rect 22388 3126 22416 6695
rect 22480 5778 22508 8026
rect 22558 7984 22614 7993
rect 22558 7919 22614 7928
rect 22572 7342 22600 7919
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22572 7041 22600 7142
rect 22558 7032 22614 7041
rect 22756 7002 22784 9540
rect 23032 9586 23060 10746
rect 23124 10470 23152 11834
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23400 10962 23428 11222
rect 23492 11121 23520 11222
rect 23952 11150 23980 11630
rect 23940 11144 23992 11150
rect 23478 11112 23534 11121
rect 23940 11086 23992 11092
rect 23478 11047 23534 11056
rect 24216 11076 24268 11082
rect 24216 11018 24268 11024
rect 23400 10934 23796 10962
rect 23296 10736 23348 10742
rect 23296 10678 23348 10684
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23112 10464 23164 10470
rect 23112 10406 23164 10412
rect 23204 10464 23256 10470
rect 23204 10406 23256 10412
rect 23124 9926 23152 10406
rect 23216 10266 23244 10406
rect 23308 10266 23336 10678
rect 23400 10577 23428 10678
rect 23386 10568 23442 10577
rect 23386 10503 23442 10512
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23296 9988 23348 9994
rect 23296 9930 23348 9936
rect 23112 9920 23164 9926
rect 23112 9862 23164 9868
rect 23308 9761 23336 9930
rect 23400 9897 23428 10503
rect 23480 10056 23532 10062
rect 23478 10024 23480 10033
rect 23532 10024 23534 10033
rect 23478 9959 23534 9968
rect 23480 9920 23532 9926
rect 23386 9888 23442 9897
rect 23480 9862 23532 9868
rect 23386 9823 23442 9832
rect 23294 9752 23350 9761
rect 23492 9738 23520 9862
rect 23294 9687 23350 9696
rect 23400 9710 23520 9738
rect 23572 9716 23624 9722
rect 22926 9551 22982 9560
rect 23020 9580 23072 9586
rect 22836 9522 22888 9528
rect 23020 9522 23072 9528
rect 23296 9512 23348 9518
rect 23296 9454 23348 9460
rect 23112 9444 23164 9450
rect 23112 9386 23164 9392
rect 22928 9036 22980 9042
rect 22928 8978 22980 8984
rect 22834 8936 22890 8945
rect 22834 8871 22890 8880
rect 22848 7449 22876 8871
rect 22834 7440 22890 7449
rect 22834 7375 22890 7384
rect 22836 7200 22888 7206
rect 22836 7142 22888 7148
rect 22558 6967 22614 6976
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22652 6928 22704 6934
rect 22652 6870 22704 6876
rect 22742 6896 22798 6905
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22572 6254 22600 6734
rect 22664 6390 22692 6870
rect 22742 6831 22798 6840
rect 22652 6384 22704 6390
rect 22652 6326 22704 6332
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22652 6248 22704 6254
rect 22652 6190 22704 6196
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 22572 5574 22600 6054
rect 22664 5710 22692 6190
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 22560 5568 22612 5574
rect 22560 5510 22612 5516
rect 22480 3466 22508 5510
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 22376 3120 22428 3126
rect 22376 3062 22428 3068
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22296 2446 22324 2994
rect 22572 2446 22600 5510
rect 22756 4826 22784 6831
rect 22744 4820 22796 4826
rect 22744 4762 22796 4768
rect 22848 4706 22876 7142
rect 22940 6866 22968 8978
rect 23020 7472 23072 7478
rect 23020 7414 23072 7420
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 22928 5908 22980 5914
rect 22928 5850 22980 5856
rect 22940 4826 22968 5850
rect 23032 5778 23060 7414
rect 23124 6662 23152 9386
rect 23308 9382 23336 9454
rect 23204 9376 23256 9382
rect 23204 9318 23256 9324
rect 23296 9376 23348 9382
rect 23400 9353 23428 9710
rect 23572 9658 23624 9664
rect 23584 9382 23612 9658
rect 23572 9376 23624 9382
rect 23296 9318 23348 9324
rect 23386 9344 23442 9353
rect 23216 9178 23244 9318
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 23308 9110 23336 9318
rect 23572 9318 23624 9324
rect 23386 9279 23442 9288
rect 23570 9208 23626 9217
rect 23570 9143 23626 9152
rect 23296 9104 23348 9110
rect 23296 9046 23348 9052
rect 23584 9042 23612 9143
rect 23572 9036 23624 9042
rect 23572 8978 23624 8984
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23204 7268 23256 7274
rect 23204 7210 23256 7216
rect 23112 6656 23164 6662
rect 23112 6598 23164 6604
rect 23020 5772 23072 5778
rect 23020 5714 23072 5720
rect 23112 5160 23164 5166
rect 23112 5102 23164 5108
rect 23020 5024 23072 5030
rect 23020 4966 23072 4972
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 22848 4678 22968 4706
rect 23032 4690 23060 4966
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22652 4072 22704 4078
rect 22650 4040 22652 4049
rect 22704 4040 22706 4049
rect 22650 3975 22706 3984
rect 22848 3602 22876 4082
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22756 3126 22784 3334
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 22940 2854 22968 4678
rect 23020 4684 23072 4690
rect 23020 4626 23072 4632
rect 23124 3058 23152 5102
rect 23216 4729 23244 7210
rect 23308 6866 23336 8570
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23400 7546 23428 8366
rect 23492 7721 23520 8774
rect 23664 8560 23716 8566
rect 23664 8502 23716 8508
rect 23572 8016 23624 8022
rect 23572 7958 23624 7964
rect 23478 7712 23534 7721
rect 23478 7647 23534 7656
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 23388 6996 23440 7002
rect 23388 6938 23440 6944
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 23296 6248 23348 6254
rect 23296 6190 23348 6196
rect 23202 4720 23258 4729
rect 23202 4655 23258 4664
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23216 3194 23244 3470
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23308 2961 23336 6190
rect 23400 3398 23428 6938
rect 23492 6866 23520 7142
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23584 6798 23612 7958
rect 23676 7818 23704 8502
rect 23768 8362 23796 10934
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 10130 23888 10406
rect 24136 10146 24164 10542
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 23952 10118 24164 10146
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23664 7812 23716 7818
rect 23664 7754 23716 7760
rect 23664 7336 23716 7342
rect 23768 7324 23796 8298
rect 23716 7296 23796 7324
rect 23664 7278 23716 7284
rect 23664 7200 23716 7206
rect 23664 7142 23716 7148
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23480 6248 23532 6254
rect 23480 6190 23532 6196
rect 23492 5846 23520 6190
rect 23480 5840 23532 5846
rect 23480 5782 23532 5788
rect 23572 5772 23624 5778
rect 23572 5714 23624 5720
rect 23480 5636 23532 5642
rect 23480 5578 23532 5584
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 23294 2952 23350 2961
rect 23294 2887 23350 2896
rect 22928 2848 22980 2854
rect 22928 2790 22980 2796
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 22848 2310 22876 2450
rect 22100 2304 22152 2310
rect 22100 2246 22152 2252
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 22112 2038 22140 2246
rect 22100 2032 22152 2038
rect 22100 1974 22152 1980
rect 22558 1456 22614 1465
rect 22558 1391 22614 1400
rect 22572 800 22600 1391
rect 23124 870 23244 898
rect 21732 332 21784 338
rect 21732 274 21784 280
rect 21640 264 21692 270
rect 21640 206 21692 212
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23124 202 23152 870
rect 23216 800 23244 870
rect 23112 196 23164 202
rect 23112 138 23164 144
rect 23202 0 23258 800
rect 23492 134 23520 5578
rect 23584 5302 23612 5714
rect 23676 5370 23704 7142
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23768 6322 23796 6734
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23754 5944 23810 5953
rect 23754 5879 23810 5888
rect 23768 5846 23796 5879
rect 23860 5846 23888 9318
rect 23952 8294 23980 10118
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 24136 9722 24164 9998
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 24228 9450 24256 11018
rect 24216 9444 24268 9450
rect 24216 9386 24268 9392
rect 24320 9058 24348 11698
rect 24688 11354 24716 12135
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 24768 11756 24820 11762
rect 24768 11698 24820 11704
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 24492 11212 24544 11218
rect 24492 11154 24544 11160
rect 24398 10568 24454 10577
rect 24398 10503 24454 10512
rect 24228 9030 24348 9058
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 23940 8288 23992 8294
rect 23940 8230 23992 8236
rect 23940 8016 23992 8022
rect 23940 7958 23992 7964
rect 23952 7886 23980 7958
rect 24044 7954 24072 8366
rect 24228 8022 24256 9030
rect 24308 8968 24360 8974
rect 24308 8910 24360 8916
rect 24320 8537 24348 8910
rect 24306 8528 24362 8537
rect 24306 8463 24362 8472
rect 24308 8424 24360 8430
rect 24308 8366 24360 8372
rect 24216 8016 24268 8022
rect 24122 7984 24178 7993
rect 24032 7948 24084 7954
rect 24216 7958 24268 7964
rect 24122 7919 24124 7928
rect 24032 7890 24084 7896
rect 24176 7919 24178 7928
rect 24124 7890 24176 7896
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23952 7721 23980 7822
rect 23938 7712 23994 7721
rect 23938 7647 23994 7656
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 23952 6798 23980 7278
rect 24044 6934 24072 7890
rect 24032 6928 24084 6934
rect 24032 6870 24084 6876
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23756 5840 23808 5846
rect 23756 5782 23808 5788
rect 23848 5840 23900 5846
rect 23848 5782 23900 5788
rect 23756 5704 23808 5710
rect 23754 5672 23756 5681
rect 23848 5704 23900 5710
rect 23808 5672 23810 5681
rect 23848 5646 23900 5652
rect 23754 5607 23810 5616
rect 23664 5364 23716 5370
rect 23664 5306 23716 5312
rect 23860 5302 23888 5646
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23848 5296 23900 5302
rect 23848 5238 23900 5244
rect 23756 5024 23808 5030
rect 23860 5001 23888 5238
rect 23756 4966 23808 4972
rect 23846 4992 23902 5001
rect 23662 4720 23718 4729
rect 23662 4655 23718 4664
rect 23676 4486 23704 4655
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23584 3126 23612 4082
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23572 3120 23624 3126
rect 23572 3062 23624 3068
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23584 1970 23612 2926
rect 23572 1964 23624 1970
rect 23572 1906 23624 1912
rect 23676 1465 23704 4014
rect 23768 3777 23796 4966
rect 23846 4927 23902 4936
rect 23754 3768 23810 3777
rect 23754 3703 23810 3712
rect 23952 2514 23980 6598
rect 24044 5370 24072 6870
rect 24124 6860 24176 6866
rect 24228 6848 24256 7958
rect 24176 6820 24256 6848
rect 24320 6848 24348 8366
rect 24412 7342 24440 10503
rect 24504 9654 24532 11154
rect 24688 11150 24716 11290
rect 24780 11150 24808 11698
rect 24860 11620 24912 11626
rect 24860 11562 24912 11568
rect 24872 11218 24900 11562
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 25332 11150 25360 11834
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24768 11144 24820 11150
rect 24952 11144 25004 11150
rect 24768 11086 24820 11092
rect 24950 11112 24952 11121
rect 25320 11144 25372 11150
rect 25004 11112 25006 11121
rect 24860 11076 24912 11082
rect 25320 11086 25372 11092
rect 24950 11047 25006 11056
rect 24860 11018 24912 11024
rect 24584 11008 24636 11014
rect 24584 10950 24636 10956
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 24596 10606 24624 10950
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24688 10470 24716 10950
rect 24584 10464 24636 10470
rect 24584 10406 24636 10412
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 24492 9648 24544 9654
rect 24492 9590 24544 9596
rect 24504 9353 24532 9590
rect 24490 9344 24546 9353
rect 24490 9279 24546 9288
rect 24492 8968 24544 8974
rect 24492 8910 24544 8916
rect 24504 8129 24532 8910
rect 24490 8120 24546 8129
rect 24490 8055 24546 8064
rect 24492 7472 24544 7478
rect 24492 7414 24544 7420
rect 24400 7336 24452 7342
rect 24400 7278 24452 7284
rect 24504 7002 24532 7414
rect 24492 6996 24544 7002
rect 24492 6938 24544 6944
rect 24492 6860 24544 6866
rect 24320 6820 24492 6848
rect 24124 6802 24176 6808
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 24044 4146 24072 5306
rect 24136 5098 24164 6258
rect 24124 5092 24176 5098
rect 24124 5034 24176 5040
rect 24124 4684 24176 4690
rect 24124 4626 24176 4632
rect 24136 4214 24164 4626
rect 24124 4208 24176 4214
rect 24124 4150 24176 4156
rect 24032 4140 24084 4146
rect 24032 4082 24084 4088
rect 24136 3466 24164 4150
rect 24228 3670 24256 6820
rect 24492 6802 24544 6808
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24412 6254 24440 6394
rect 24400 6248 24452 6254
rect 24400 6190 24452 6196
rect 24308 5840 24360 5846
rect 24360 5800 24440 5828
rect 24308 5782 24360 5788
rect 24308 5092 24360 5098
rect 24308 5034 24360 5040
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24124 3460 24176 3466
rect 24124 3402 24176 3408
rect 24320 2650 24348 5034
rect 24412 4758 24440 5800
rect 24492 5704 24544 5710
rect 24492 5646 24544 5652
rect 24400 4752 24452 4758
rect 24400 4694 24452 4700
rect 24412 3534 24440 4694
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 24504 3482 24532 5646
rect 24596 4842 24624 10406
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24688 9654 24716 10202
rect 24676 9648 24728 9654
rect 24676 9590 24728 9596
rect 24674 9480 24730 9489
rect 24674 9415 24676 9424
rect 24728 9415 24730 9424
rect 24676 9386 24728 9392
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 24688 6458 24716 8366
rect 24780 8022 24808 10950
rect 24768 8016 24820 8022
rect 24768 7958 24820 7964
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24780 7274 24808 7686
rect 24768 7268 24820 7274
rect 24768 7210 24820 7216
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24768 5908 24820 5914
rect 24768 5850 24820 5856
rect 24780 5250 24808 5850
rect 24872 5370 24900 11018
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 25148 10146 25176 10542
rect 25424 10470 25452 10542
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25056 10118 25176 10146
rect 25056 9926 25084 10118
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 25148 8974 25176 9998
rect 25424 9926 25452 10406
rect 25516 10062 25544 24074
rect 25700 12209 25728 26862
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 25686 12200 25742 12209
rect 25608 12158 25686 12186
rect 25608 10062 25636 12158
rect 25686 12135 25742 12144
rect 25688 12096 25740 12102
rect 25688 12038 25740 12044
rect 25700 11150 25728 12038
rect 25976 11626 26004 14418
rect 25964 11620 26016 11626
rect 25884 11580 25964 11608
rect 25688 11144 25740 11150
rect 25688 11086 25740 11092
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25792 10577 25820 11086
rect 25778 10568 25834 10577
rect 25778 10503 25834 10512
rect 25504 10056 25556 10062
rect 25504 9998 25556 10004
rect 25596 10056 25648 10062
rect 25596 9998 25648 10004
rect 25228 9920 25280 9926
rect 25228 9862 25280 9868
rect 25412 9920 25464 9926
rect 25412 9862 25464 9868
rect 25240 9518 25268 9862
rect 25516 9518 25544 9998
rect 25608 9761 25636 9998
rect 25884 9994 25912 11580
rect 25964 11562 26016 11568
rect 26068 10606 26096 29582
rect 26240 11756 26292 11762
rect 26240 11698 26292 11704
rect 26252 11150 26280 11698
rect 26344 11150 26372 32370
rect 27356 16574 27384 33050
rect 29288 17882 29316 37198
rect 29840 36854 29868 39200
rect 31680 37262 31708 39200
rect 33520 37330 33548 39200
rect 33508 37324 33560 37330
rect 33508 37266 33560 37272
rect 31668 37256 31720 37262
rect 31668 37198 31720 37204
rect 32772 37256 32824 37262
rect 32772 37198 32824 37204
rect 33784 37256 33836 37262
rect 33784 37198 33836 37204
rect 29828 36848 29880 36854
rect 29828 36790 29880 36796
rect 32784 36553 32812 37198
rect 33796 36922 33824 37198
rect 33784 36916 33836 36922
rect 33784 36858 33836 36864
rect 35360 36718 35388 39200
rect 35854 37564 36162 37573
rect 35854 37562 35860 37564
rect 35916 37562 35940 37564
rect 35996 37562 36020 37564
rect 36076 37562 36100 37564
rect 36156 37562 36162 37564
rect 35916 37510 35918 37562
rect 36098 37510 36100 37562
rect 35854 37508 35860 37510
rect 35916 37508 35940 37510
rect 35996 37508 36020 37510
rect 36076 37508 36100 37510
rect 36156 37508 36162 37510
rect 35854 37499 36162 37508
rect 37200 37262 37228 39200
rect 39040 37330 39068 39200
rect 40880 37618 40908 39200
rect 40880 37590 41092 37618
rect 39028 37324 39080 37330
rect 39028 37266 39080 37272
rect 41064 37262 41092 37590
rect 37004 37256 37056 37262
rect 37004 37198 37056 37204
rect 37188 37256 37240 37262
rect 37188 37198 37240 37204
rect 39120 37256 39172 37262
rect 39120 37198 39172 37204
rect 40868 37256 40920 37262
rect 40868 37198 40920 37204
rect 41052 37256 41104 37262
rect 41052 37198 41104 37204
rect 36514 37020 36822 37029
rect 36514 37018 36520 37020
rect 36576 37018 36600 37020
rect 36656 37018 36680 37020
rect 36736 37018 36760 37020
rect 36816 37018 36822 37020
rect 36576 36966 36578 37018
rect 36758 36966 36760 37018
rect 36514 36964 36520 36966
rect 36576 36964 36600 36966
rect 36656 36964 36680 36966
rect 36736 36964 36760 36966
rect 36816 36964 36822 36966
rect 36514 36955 36822 36964
rect 37016 36922 37044 37198
rect 37004 36916 37056 36922
rect 37004 36858 37056 36864
rect 35440 36780 35492 36786
rect 35440 36722 35492 36728
rect 35348 36712 35400 36718
rect 35348 36654 35400 36660
rect 32770 36544 32826 36553
rect 32770 36479 32826 36488
rect 35452 17882 35480 36722
rect 35854 36476 36162 36485
rect 35854 36474 35860 36476
rect 35916 36474 35940 36476
rect 35996 36474 36020 36476
rect 36076 36474 36100 36476
rect 36156 36474 36162 36476
rect 35916 36422 35918 36474
rect 36098 36422 36100 36474
rect 35854 36420 35860 36422
rect 35916 36420 35940 36422
rect 35996 36420 36020 36422
rect 36076 36420 36100 36422
rect 36156 36420 36162 36422
rect 35854 36411 36162 36420
rect 36514 35932 36822 35941
rect 36514 35930 36520 35932
rect 36576 35930 36600 35932
rect 36656 35930 36680 35932
rect 36736 35930 36760 35932
rect 36816 35930 36822 35932
rect 36576 35878 36578 35930
rect 36758 35878 36760 35930
rect 36514 35876 36520 35878
rect 36576 35876 36600 35878
rect 36656 35876 36680 35878
rect 36736 35876 36760 35878
rect 36816 35876 36822 35878
rect 36514 35867 36822 35876
rect 35854 35388 36162 35397
rect 35854 35386 35860 35388
rect 35916 35386 35940 35388
rect 35996 35386 36020 35388
rect 36076 35386 36100 35388
rect 36156 35386 36162 35388
rect 35916 35334 35918 35386
rect 36098 35334 36100 35386
rect 35854 35332 35860 35334
rect 35916 35332 35940 35334
rect 35996 35332 36020 35334
rect 36076 35332 36100 35334
rect 36156 35332 36162 35334
rect 35854 35323 36162 35332
rect 36514 34844 36822 34853
rect 36514 34842 36520 34844
rect 36576 34842 36600 34844
rect 36656 34842 36680 34844
rect 36736 34842 36760 34844
rect 36816 34842 36822 34844
rect 36576 34790 36578 34842
rect 36758 34790 36760 34842
rect 36514 34788 36520 34790
rect 36576 34788 36600 34790
rect 36656 34788 36680 34790
rect 36736 34788 36760 34790
rect 36816 34788 36822 34790
rect 36514 34779 36822 34788
rect 35854 34300 36162 34309
rect 35854 34298 35860 34300
rect 35916 34298 35940 34300
rect 35996 34298 36020 34300
rect 36076 34298 36100 34300
rect 36156 34298 36162 34300
rect 35916 34246 35918 34298
rect 36098 34246 36100 34298
rect 35854 34244 35860 34246
rect 35916 34244 35940 34246
rect 35996 34244 36020 34246
rect 36076 34244 36100 34246
rect 36156 34244 36162 34246
rect 35854 34235 36162 34244
rect 36514 33756 36822 33765
rect 36514 33754 36520 33756
rect 36576 33754 36600 33756
rect 36656 33754 36680 33756
rect 36736 33754 36760 33756
rect 36816 33754 36822 33756
rect 36576 33702 36578 33754
rect 36758 33702 36760 33754
rect 36514 33700 36520 33702
rect 36576 33700 36600 33702
rect 36656 33700 36680 33702
rect 36736 33700 36760 33702
rect 36816 33700 36822 33702
rect 36514 33691 36822 33700
rect 35854 33212 36162 33221
rect 35854 33210 35860 33212
rect 35916 33210 35940 33212
rect 35996 33210 36020 33212
rect 36076 33210 36100 33212
rect 36156 33210 36162 33212
rect 35916 33158 35918 33210
rect 36098 33158 36100 33210
rect 35854 33156 35860 33158
rect 35916 33156 35940 33158
rect 35996 33156 36020 33158
rect 36076 33156 36100 33158
rect 36156 33156 36162 33158
rect 35854 33147 36162 33156
rect 36514 32668 36822 32677
rect 36514 32666 36520 32668
rect 36576 32666 36600 32668
rect 36656 32666 36680 32668
rect 36736 32666 36760 32668
rect 36816 32666 36822 32668
rect 36576 32614 36578 32666
rect 36758 32614 36760 32666
rect 36514 32612 36520 32614
rect 36576 32612 36600 32614
rect 36656 32612 36680 32614
rect 36736 32612 36760 32614
rect 36816 32612 36822 32614
rect 36514 32603 36822 32612
rect 35854 32124 36162 32133
rect 35854 32122 35860 32124
rect 35916 32122 35940 32124
rect 35996 32122 36020 32124
rect 36076 32122 36100 32124
rect 36156 32122 36162 32124
rect 35916 32070 35918 32122
rect 36098 32070 36100 32122
rect 35854 32068 35860 32070
rect 35916 32068 35940 32070
rect 35996 32068 36020 32070
rect 36076 32068 36100 32070
rect 36156 32068 36162 32070
rect 35854 32059 36162 32068
rect 36514 31580 36822 31589
rect 36514 31578 36520 31580
rect 36576 31578 36600 31580
rect 36656 31578 36680 31580
rect 36736 31578 36760 31580
rect 36816 31578 36822 31580
rect 36576 31526 36578 31578
rect 36758 31526 36760 31578
rect 36514 31524 36520 31526
rect 36576 31524 36600 31526
rect 36656 31524 36680 31526
rect 36736 31524 36760 31526
rect 36816 31524 36822 31526
rect 36514 31515 36822 31524
rect 35854 31036 36162 31045
rect 35854 31034 35860 31036
rect 35916 31034 35940 31036
rect 35996 31034 36020 31036
rect 36076 31034 36100 31036
rect 36156 31034 36162 31036
rect 35916 30982 35918 31034
rect 36098 30982 36100 31034
rect 35854 30980 35860 30982
rect 35916 30980 35940 30982
rect 35996 30980 36020 30982
rect 36076 30980 36100 30982
rect 36156 30980 36162 30982
rect 35854 30971 36162 30980
rect 36514 30492 36822 30501
rect 36514 30490 36520 30492
rect 36576 30490 36600 30492
rect 36656 30490 36680 30492
rect 36736 30490 36760 30492
rect 36816 30490 36822 30492
rect 36576 30438 36578 30490
rect 36758 30438 36760 30490
rect 36514 30436 36520 30438
rect 36576 30436 36600 30438
rect 36656 30436 36680 30438
rect 36736 30436 36760 30438
rect 36816 30436 36822 30438
rect 36514 30427 36822 30436
rect 35854 29948 36162 29957
rect 35854 29946 35860 29948
rect 35916 29946 35940 29948
rect 35996 29946 36020 29948
rect 36076 29946 36100 29948
rect 36156 29946 36162 29948
rect 35916 29894 35918 29946
rect 36098 29894 36100 29946
rect 35854 29892 35860 29894
rect 35916 29892 35940 29894
rect 35996 29892 36020 29894
rect 36076 29892 36100 29894
rect 36156 29892 36162 29894
rect 35854 29883 36162 29892
rect 36514 29404 36822 29413
rect 36514 29402 36520 29404
rect 36576 29402 36600 29404
rect 36656 29402 36680 29404
rect 36736 29402 36760 29404
rect 36816 29402 36822 29404
rect 36576 29350 36578 29402
rect 36758 29350 36760 29402
rect 36514 29348 36520 29350
rect 36576 29348 36600 29350
rect 36656 29348 36680 29350
rect 36736 29348 36760 29350
rect 36816 29348 36822 29350
rect 36514 29339 36822 29348
rect 35854 28860 36162 28869
rect 35854 28858 35860 28860
rect 35916 28858 35940 28860
rect 35996 28858 36020 28860
rect 36076 28858 36100 28860
rect 36156 28858 36162 28860
rect 35916 28806 35918 28858
rect 36098 28806 36100 28858
rect 35854 28804 35860 28806
rect 35916 28804 35940 28806
rect 35996 28804 36020 28806
rect 36076 28804 36100 28806
rect 36156 28804 36162 28806
rect 35854 28795 36162 28804
rect 36514 28316 36822 28325
rect 36514 28314 36520 28316
rect 36576 28314 36600 28316
rect 36656 28314 36680 28316
rect 36736 28314 36760 28316
rect 36816 28314 36822 28316
rect 36576 28262 36578 28314
rect 36758 28262 36760 28314
rect 36514 28260 36520 28262
rect 36576 28260 36600 28262
rect 36656 28260 36680 28262
rect 36736 28260 36760 28262
rect 36816 28260 36822 28262
rect 36514 28251 36822 28260
rect 35854 27772 36162 27781
rect 35854 27770 35860 27772
rect 35916 27770 35940 27772
rect 35996 27770 36020 27772
rect 36076 27770 36100 27772
rect 36156 27770 36162 27772
rect 35916 27718 35918 27770
rect 36098 27718 36100 27770
rect 35854 27716 35860 27718
rect 35916 27716 35940 27718
rect 35996 27716 36020 27718
rect 36076 27716 36100 27718
rect 36156 27716 36162 27718
rect 35854 27707 36162 27716
rect 36514 27228 36822 27237
rect 36514 27226 36520 27228
rect 36576 27226 36600 27228
rect 36656 27226 36680 27228
rect 36736 27226 36760 27228
rect 36816 27226 36822 27228
rect 36576 27174 36578 27226
rect 36758 27174 36760 27226
rect 36514 27172 36520 27174
rect 36576 27172 36600 27174
rect 36656 27172 36680 27174
rect 36736 27172 36760 27174
rect 36816 27172 36822 27174
rect 36514 27163 36822 27172
rect 35854 26684 36162 26693
rect 35854 26682 35860 26684
rect 35916 26682 35940 26684
rect 35996 26682 36020 26684
rect 36076 26682 36100 26684
rect 36156 26682 36162 26684
rect 35916 26630 35918 26682
rect 36098 26630 36100 26682
rect 35854 26628 35860 26630
rect 35916 26628 35940 26630
rect 35996 26628 36020 26630
rect 36076 26628 36100 26630
rect 36156 26628 36162 26630
rect 35854 26619 36162 26628
rect 36514 26140 36822 26149
rect 36514 26138 36520 26140
rect 36576 26138 36600 26140
rect 36656 26138 36680 26140
rect 36736 26138 36760 26140
rect 36816 26138 36822 26140
rect 36576 26086 36578 26138
rect 36758 26086 36760 26138
rect 36514 26084 36520 26086
rect 36576 26084 36600 26086
rect 36656 26084 36680 26086
rect 36736 26084 36760 26086
rect 36816 26084 36822 26086
rect 36514 26075 36822 26084
rect 35854 25596 36162 25605
rect 35854 25594 35860 25596
rect 35916 25594 35940 25596
rect 35996 25594 36020 25596
rect 36076 25594 36100 25596
rect 36156 25594 36162 25596
rect 35916 25542 35918 25594
rect 36098 25542 36100 25594
rect 35854 25540 35860 25542
rect 35916 25540 35940 25542
rect 35996 25540 36020 25542
rect 36076 25540 36100 25542
rect 36156 25540 36162 25542
rect 35854 25531 36162 25540
rect 36514 25052 36822 25061
rect 36514 25050 36520 25052
rect 36576 25050 36600 25052
rect 36656 25050 36680 25052
rect 36736 25050 36760 25052
rect 36816 25050 36822 25052
rect 36576 24998 36578 25050
rect 36758 24998 36760 25050
rect 36514 24996 36520 24998
rect 36576 24996 36600 24998
rect 36656 24996 36680 24998
rect 36736 24996 36760 24998
rect 36816 24996 36822 24998
rect 36514 24987 36822 24996
rect 35854 24508 36162 24517
rect 35854 24506 35860 24508
rect 35916 24506 35940 24508
rect 35996 24506 36020 24508
rect 36076 24506 36100 24508
rect 36156 24506 36162 24508
rect 35916 24454 35918 24506
rect 36098 24454 36100 24506
rect 35854 24452 35860 24454
rect 35916 24452 35940 24454
rect 35996 24452 36020 24454
rect 36076 24452 36100 24454
rect 36156 24452 36162 24454
rect 35854 24443 36162 24452
rect 36514 23964 36822 23973
rect 36514 23962 36520 23964
rect 36576 23962 36600 23964
rect 36656 23962 36680 23964
rect 36736 23962 36760 23964
rect 36816 23962 36822 23964
rect 36576 23910 36578 23962
rect 36758 23910 36760 23962
rect 36514 23908 36520 23910
rect 36576 23908 36600 23910
rect 36656 23908 36680 23910
rect 36736 23908 36760 23910
rect 36816 23908 36822 23910
rect 36514 23899 36822 23908
rect 35854 23420 36162 23429
rect 35854 23418 35860 23420
rect 35916 23418 35940 23420
rect 35996 23418 36020 23420
rect 36076 23418 36100 23420
rect 36156 23418 36162 23420
rect 35916 23366 35918 23418
rect 36098 23366 36100 23418
rect 35854 23364 35860 23366
rect 35916 23364 35940 23366
rect 35996 23364 36020 23366
rect 36076 23364 36100 23366
rect 36156 23364 36162 23366
rect 35854 23355 36162 23364
rect 36514 22876 36822 22885
rect 36514 22874 36520 22876
rect 36576 22874 36600 22876
rect 36656 22874 36680 22876
rect 36736 22874 36760 22876
rect 36816 22874 36822 22876
rect 36576 22822 36578 22874
rect 36758 22822 36760 22874
rect 36514 22820 36520 22822
rect 36576 22820 36600 22822
rect 36656 22820 36680 22822
rect 36736 22820 36760 22822
rect 36816 22820 36822 22822
rect 36514 22811 36822 22820
rect 35854 22332 36162 22341
rect 35854 22330 35860 22332
rect 35916 22330 35940 22332
rect 35996 22330 36020 22332
rect 36076 22330 36100 22332
rect 36156 22330 36162 22332
rect 35916 22278 35918 22330
rect 36098 22278 36100 22330
rect 35854 22276 35860 22278
rect 35916 22276 35940 22278
rect 35996 22276 36020 22278
rect 36076 22276 36100 22278
rect 36156 22276 36162 22278
rect 35854 22267 36162 22276
rect 36514 21788 36822 21797
rect 36514 21786 36520 21788
rect 36576 21786 36600 21788
rect 36656 21786 36680 21788
rect 36736 21786 36760 21788
rect 36816 21786 36822 21788
rect 36576 21734 36578 21786
rect 36758 21734 36760 21786
rect 36514 21732 36520 21734
rect 36576 21732 36600 21734
rect 36656 21732 36680 21734
rect 36736 21732 36760 21734
rect 36816 21732 36822 21734
rect 36514 21723 36822 21732
rect 35854 21244 36162 21253
rect 35854 21242 35860 21244
rect 35916 21242 35940 21244
rect 35996 21242 36020 21244
rect 36076 21242 36100 21244
rect 36156 21242 36162 21244
rect 35916 21190 35918 21242
rect 36098 21190 36100 21242
rect 35854 21188 35860 21190
rect 35916 21188 35940 21190
rect 35996 21188 36020 21190
rect 36076 21188 36100 21190
rect 36156 21188 36162 21190
rect 35854 21179 36162 21188
rect 36514 20700 36822 20709
rect 36514 20698 36520 20700
rect 36576 20698 36600 20700
rect 36656 20698 36680 20700
rect 36736 20698 36760 20700
rect 36816 20698 36822 20700
rect 36576 20646 36578 20698
rect 36758 20646 36760 20698
rect 36514 20644 36520 20646
rect 36576 20644 36600 20646
rect 36656 20644 36680 20646
rect 36736 20644 36760 20646
rect 36816 20644 36822 20646
rect 36514 20635 36822 20644
rect 35854 20156 36162 20165
rect 35854 20154 35860 20156
rect 35916 20154 35940 20156
rect 35996 20154 36020 20156
rect 36076 20154 36100 20156
rect 36156 20154 36162 20156
rect 35916 20102 35918 20154
rect 36098 20102 36100 20154
rect 35854 20100 35860 20102
rect 35916 20100 35940 20102
rect 35996 20100 36020 20102
rect 36076 20100 36100 20102
rect 36156 20100 36162 20102
rect 35854 20091 36162 20100
rect 36514 19612 36822 19621
rect 36514 19610 36520 19612
rect 36576 19610 36600 19612
rect 36656 19610 36680 19612
rect 36736 19610 36760 19612
rect 36816 19610 36822 19612
rect 36576 19558 36578 19610
rect 36758 19558 36760 19610
rect 36514 19556 36520 19558
rect 36576 19556 36600 19558
rect 36656 19556 36680 19558
rect 36736 19556 36760 19558
rect 36816 19556 36822 19558
rect 36514 19547 36822 19556
rect 35854 19068 36162 19077
rect 35854 19066 35860 19068
rect 35916 19066 35940 19068
rect 35996 19066 36020 19068
rect 36076 19066 36100 19068
rect 36156 19066 36162 19068
rect 35916 19014 35918 19066
rect 36098 19014 36100 19066
rect 35854 19012 35860 19014
rect 35916 19012 35940 19014
rect 35996 19012 36020 19014
rect 36076 19012 36100 19014
rect 36156 19012 36162 19014
rect 35854 19003 36162 19012
rect 36514 18524 36822 18533
rect 36514 18522 36520 18524
rect 36576 18522 36600 18524
rect 36656 18522 36680 18524
rect 36736 18522 36760 18524
rect 36816 18522 36822 18524
rect 36576 18470 36578 18522
rect 36758 18470 36760 18522
rect 36514 18468 36520 18470
rect 36576 18468 36600 18470
rect 36656 18468 36680 18470
rect 36736 18468 36760 18470
rect 36816 18468 36822 18470
rect 36514 18459 36822 18468
rect 35854 17980 36162 17989
rect 35854 17978 35860 17980
rect 35916 17978 35940 17980
rect 35996 17978 36020 17980
rect 36076 17978 36100 17980
rect 36156 17978 36162 17980
rect 35916 17926 35918 17978
rect 36098 17926 36100 17978
rect 35854 17924 35860 17926
rect 35916 17924 35940 17926
rect 35996 17924 36020 17926
rect 36076 17924 36100 17926
rect 36156 17924 36162 17926
rect 35854 17915 36162 17924
rect 29276 17876 29328 17882
rect 29276 17818 29328 17824
rect 31116 17876 31168 17882
rect 31116 17818 31168 17824
rect 31668 17876 31720 17882
rect 31668 17818 31720 17824
rect 35440 17876 35492 17882
rect 35440 17818 35492 17824
rect 26804 16546 27384 16574
rect 31128 16574 31156 17818
rect 31680 16574 31708 17818
rect 36514 17436 36822 17445
rect 36514 17434 36520 17436
rect 36576 17434 36600 17436
rect 36656 17434 36680 17436
rect 36736 17434 36760 17436
rect 36816 17434 36822 17436
rect 36576 17382 36578 17434
rect 36758 17382 36760 17434
rect 36514 17380 36520 17382
rect 36576 17380 36600 17382
rect 36656 17380 36680 17382
rect 36736 17380 36760 17382
rect 36816 17380 36822 17382
rect 36514 17371 36822 17380
rect 35854 16892 36162 16901
rect 35854 16890 35860 16892
rect 35916 16890 35940 16892
rect 35996 16890 36020 16892
rect 36076 16890 36100 16892
rect 36156 16890 36162 16892
rect 35916 16838 35918 16890
rect 36098 16838 36100 16890
rect 35854 16836 35860 16838
rect 35916 16836 35940 16838
rect 35996 16836 36020 16838
rect 36076 16836 36100 16838
rect 36156 16836 36162 16838
rect 35854 16827 36162 16836
rect 31128 16546 31524 16574
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26332 11144 26384 11150
rect 26332 11086 26384 11092
rect 26700 11144 26752 11150
rect 26700 11086 26752 11092
rect 26056 10600 26108 10606
rect 26240 10600 26292 10606
rect 26056 10542 26108 10548
rect 26238 10568 26240 10577
rect 26292 10568 26294 10577
rect 26238 10503 26294 10512
rect 25964 10464 26016 10470
rect 25964 10406 26016 10412
rect 26056 10464 26108 10470
rect 26056 10406 26108 10412
rect 25872 9988 25924 9994
rect 25872 9930 25924 9936
rect 25594 9752 25650 9761
rect 25594 9687 25650 9696
rect 25976 9586 26004 10406
rect 26068 10062 26096 10406
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 26148 9920 26200 9926
rect 26148 9862 26200 9868
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 25056 8537 25084 8774
rect 25042 8528 25098 8537
rect 25042 8463 25098 8472
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 25056 7585 25084 7822
rect 25042 7576 25098 7585
rect 25042 7511 25098 7520
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24780 5222 24900 5250
rect 24596 4814 24716 4842
rect 24688 3534 24716 4814
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 24676 3528 24728 3534
rect 24504 3454 24624 3482
rect 24676 3470 24728 3476
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24398 2680 24454 2689
rect 24308 2644 24360 2650
rect 24398 2615 24454 2624
rect 24308 2586 24360 2592
rect 24412 2514 24440 2615
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 23860 1970 23888 2246
rect 23848 1964 23900 1970
rect 23848 1906 23900 1912
rect 23662 1456 23718 1465
rect 23662 1391 23718 1400
rect 23846 1184 23902 1193
rect 23846 1119 23902 1128
rect 23860 800 23888 1119
rect 24504 800 24532 3334
rect 24596 3176 24624 3454
rect 24596 3148 24716 3176
rect 24582 3088 24638 3097
rect 24582 3023 24584 3032
rect 24636 3023 24638 3032
rect 24584 2994 24636 3000
rect 24688 2922 24716 3148
rect 24676 2916 24728 2922
rect 24676 2858 24728 2864
rect 24780 2514 24808 4558
rect 24872 3641 24900 5222
rect 24858 3632 24914 3641
rect 24858 3567 24914 3576
rect 24964 3074 24992 7278
rect 25056 6934 25084 7278
rect 25044 6928 25096 6934
rect 25044 6870 25096 6876
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 25056 5137 25084 6054
rect 25042 5128 25098 5137
rect 25042 5063 25098 5072
rect 25042 3496 25098 3505
rect 25042 3431 25098 3440
rect 24872 3046 24992 3074
rect 25056 3058 25084 3431
rect 25148 3097 25176 8910
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25240 4622 25268 8774
rect 25332 6905 25360 9318
rect 25516 8401 25544 9454
rect 25688 9172 25740 9178
rect 25688 9114 25740 9120
rect 25700 8430 25728 9114
rect 25964 9104 26016 9110
rect 25964 9046 26016 9052
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25688 8424 25740 8430
rect 25502 8392 25558 8401
rect 25688 8366 25740 8372
rect 25502 8327 25558 8336
rect 25596 8356 25648 8362
rect 25596 8298 25648 8304
rect 25504 8016 25556 8022
rect 25504 7958 25556 7964
rect 25318 6896 25374 6905
rect 25318 6831 25374 6840
rect 25516 6798 25544 7958
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 25412 6316 25464 6322
rect 25412 6258 25464 6264
rect 25320 6112 25372 6118
rect 25320 6054 25372 6060
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25332 3777 25360 6054
rect 25424 5574 25452 6258
rect 25504 6180 25556 6186
rect 25504 6122 25556 6128
rect 25516 5710 25544 6122
rect 25504 5704 25556 5710
rect 25504 5646 25556 5652
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 25410 5264 25466 5273
rect 25410 5199 25466 5208
rect 25424 5166 25452 5199
rect 25412 5160 25464 5166
rect 25412 5102 25464 5108
rect 25412 5024 25464 5030
rect 25410 4992 25412 5001
rect 25464 4992 25544 5012
rect 25466 4984 25544 4992
rect 25410 4927 25466 4936
rect 25412 4752 25464 4758
rect 25412 4694 25464 4700
rect 25424 4486 25452 4694
rect 25412 4480 25464 4486
rect 25412 4422 25464 4428
rect 25318 3768 25374 3777
rect 25318 3703 25374 3712
rect 25424 3482 25452 4422
rect 25516 4185 25544 4984
rect 25502 4176 25558 4185
rect 25502 4111 25558 4120
rect 25608 3670 25636 8298
rect 25688 7812 25740 7818
rect 25688 7754 25740 7760
rect 25700 6322 25728 7754
rect 25792 6458 25820 8570
rect 25872 8560 25924 8566
rect 25872 8502 25924 8508
rect 25884 7954 25912 8502
rect 25872 7948 25924 7954
rect 25872 7890 25924 7896
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 25884 7002 25912 7142
rect 25872 6996 25924 7002
rect 25872 6938 25924 6944
rect 25872 6792 25924 6798
rect 25872 6734 25924 6740
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 25688 6316 25740 6322
rect 25688 6258 25740 6264
rect 25884 6254 25912 6734
rect 25780 6248 25832 6254
rect 25780 6190 25832 6196
rect 25872 6248 25924 6254
rect 25872 6190 25924 6196
rect 25686 5808 25742 5817
rect 25686 5743 25742 5752
rect 25700 5234 25728 5743
rect 25688 5228 25740 5234
rect 25688 5170 25740 5176
rect 25596 3664 25648 3670
rect 25596 3606 25648 3612
rect 25332 3454 25452 3482
rect 25228 3188 25280 3194
rect 25228 3130 25280 3136
rect 25134 3088 25190 3097
rect 25044 3052 25096 3058
rect 24872 2854 24900 3046
rect 25240 3058 25268 3130
rect 25134 3023 25190 3032
rect 25228 3052 25280 3058
rect 25044 2994 25096 3000
rect 25228 2994 25280 3000
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 25136 2848 25188 2854
rect 25228 2848 25280 2854
rect 25136 2790 25188 2796
rect 25226 2816 25228 2825
rect 25280 2816 25282 2825
rect 25148 2666 25176 2790
rect 25226 2751 25282 2760
rect 25332 2666 25360 3454
rect 25412 3392 25464 3398
rect 25410 3360 25412 3369
rect 25688 3392 25740 3398
rect 25464 3360 25466 3369
rect 25688 3334 25740 3340
rect 25410 3295 25466 3304
rect 25410 3088 25466 3097
rect 25410 3023 25466 3032
rect 25148 2638 25360 2666
rect 25318 2544 25374 2553
rect 24768 2508 24820 2514
rect 25318 2479 25374 2488
rect 24768 2450 24820 2456
rect 25332 2446 25360 2479
rect 24584 2440 24636 2446
rect 24582 2408 24584 2417
rect 25320 2440 25372 2446
rect 24636 2408 24638 2417
rect 25320 2382 25372 2388
rect 24582 2343 24638 2352
rect 25148 870 25268 898
rect 25148 800 25176 870
rect 23480 128 23532 134
rect 23480 70 23532 76
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25240 762 25268 870
rect 25424 762 25452 3023
rect 25700 1698 25728 3334
rect 25688 1692 25740 1698
rect 25688 1634 25740 1640
rect 25792 1630 25820 6190
rect 25976 5710 26004 9046
rect 26068 8430 26096 9862
rect 26056 8424 26108 8430
rect 26056 8366 26108 8372
rect 26068 7886 26096 8366
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26068 6458 26096 6734
rect 26056 6452 26108 6458
rect 26056 6394 26108 6400
rect 25964 5704 26016 5710
rect 25964 5646 26016 5652
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 25872 4208 25924 4214
rect 25872 4150 25924 4156
rect 25884 3126 25912 4150
rect 26068 4146 26096 5510
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 25964 4072 26016 4078
rect 25962 4040 25964 4049
rect 26016 4040 26018 4049
rect 25962 3975 26018 3984
rect 26160 3602 26188 9862
rect 26344 9674 26372 11086
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 26620 10470 26648 10542
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 26344 9646 26464 9674
rect 26238 8664 26294 8673
rect 26238 8599 26294 8608
rect 26252 6610 26280 8599
rect 26330 8528 26386 8537
rect 26330 8463 26386 8472
rect 26344 6730 26372 8463
rect 26436 8430 26464 9646
rect 26516 9648 26568 9654
rect 26516 9590 26568 9596
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26528 8090 26556 9590
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 26424 7404 26476 7410
rect 26424 7346 26476 7352
rect 26332 6724 26384 6730
rect 26332 6666 26384 6672
rect 26252 6582 26372 6610
rect 26238 6488 26294 6497
rect 26238 6423 26294 6432
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 26252 3482 26280 6423
rect 26344 5409 26372 6582
rect 26330 5400 26386 5409
rect 26330 5335 26386 5344
rect 26436 4282 26464 7346
rect 26514 6352 26570 6361
rect 26514 6287 26516 6296
rect 26568 6287 26570 6296
rect 26516 6258 26568 6264
rect 26620 4758 26648 9998
rect 26712 8294 26740 11086
rect 26700 8288 26752 8294
rect 26700 8230 26752 8236
rect 26712 7954 26740 8230
rect 26700 7948 26752 7954
rect 26700 7890 26752 7896
rect 26804 7478 26832 16546
rect 27896 12708 27948 12714
rect 27896 12650 27948 12656
rect 27710 12472 27766 12481
rect 27710 12407 27766 12416
rect 27068 11824 27120 11830
rect 27068 11766 27120 11772
rect 26976 11348 27028 11354
rect 26976 11290 27028 11296
rect 26884 10600 26936 10606
rect 26884 10542 26936 10548
rect 26896 9654 26924 10542
rect 26988 9761 27016 11290
rect 27080 11150 27108 11766
rect 27252 11688 27304 11694
rect 27252 11630 27304 11636
rect 27264 11150 27292 11630
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 27068 11144 27120 11150
rect 27068 11086 27120 11092
rect 27252 11144 27304 11150
rect 27252 11086 27304 11092
rect 27344 11144 27396 11150
rect 27344 11086 27396 11092
rect 26974 9752 27030 9761
rect 26974 9687 27030 9696
rect 26884 9648 26936 9654
rect 26884 9590 26936 9596
rect 26884 8560 26936 8566
rect 26882 8528 26884 8537
rect 27080 8537 27108 11086
rect 27160 11008 27212 11014
rect 27160 10950 27212 10956
rect 27172 10266 27200 10950
rect 27160 10260 27212 10266
rect 27160 10202 27212 10208
rect 27160 9512 27212 9518
rect 27160 9454 27212 9460
rect 26936 8528 26938 8537
rect 26882 8463 26938 8472
rect 27066 8528 27122 8537
rect 27066 8463 27122 8472
rect 26976 8424 27028 8430
rect 26976 8366 27028 8372
rect 26988 7721 27016 8366
rect 26974 7712 27030 7721
rect 26974 7647 27030 7656
rect 26792 7472 26844 7478
rect 26792 7414 26844 7420
rect 26988 7410 27016 7647
rect 26976 7404 27028 7410
rect 26976 7346 27028 7352
rect 27080 7290 27108 8463
rect 27172 8401 27200 9454
rect 27264 8838 27292 11086
rect 27356 10146 27384 11086
rect 27448 10266 27476 11290
rect 27528 10464 27580 10470
rect 27528 10406 27580 10412
rect 27436 10260 27488 10266
rect 27436 10202 27488 10208
rect 27356 10118 27476 10146
rect 27344 10056 27396 10062
rect 27344 9998 27396 10004
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27158 8392 27214 8401
rect 27158 8327 27214 8336
rect 27252 8356 27304 8362
rect 27252 8298 27304 8304
rect 27158 8120 27214 8129
rect 27158 8055 27214 8064
rect 27172 7750 27200 8055
rect 27160 7744 27212 7750
rect 27160 7686 27212 7692
rect 27172 7449 27200 7686
rect 27158 7440 27214 7449
rect 27158 7375 27214 7384
rect 26712 7262 27108 7290
rect 27160 7268 27212 7274
rect 26608 4752 26660 4758
rect 26608 4694 26660 4700
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 26424 4276 26476 4282
rect 26424 4218 26476 4224
rect 26424 4140 26476 4146
rect 26424 4082 26476 4088
rect 26436 3942 26464 4082
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26160 3454 26280 3482
rect 26160 3398 26188 3454
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 25872 3120 25924 3126
rect 25872 3062 25924 3068
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 26252 2281 26280 2450
rect 26238 2272 26294 2281
rect 26238 2207 26294 2216
rect 26344 1834 26372 3334
rect 26528 2650 26556 4558
rect 26712 4282 26740 7262
rect 27160 7210 27212 7216
rect 27172 7177 27200 7210
rect 27158 7168 27214 7177
rect 27158 7103 27214 7112
rect 26790 7032 26846 7041
rect 26790 6967 26846 6976
rect 26700 4276 26752 4282
rect 26700 4218 26752 4224
rect 26698 4040 26754 4049
rect 26698 3975 26700 3984
rect 26752 3975 26754 3984
rect 26700 3946 26752 3952
rect 26608 3528 26660 3534
rect 26608 3470 26660 3476
rect 26620 3194 26648 3470
rect 26804 3398 26832 6967
rect 26976 6860 27028 6866
rect 26896 6820 26976 6848
rect 26896 5166 26924 6820
rect 26976 6802 27028 6808
rect 27264 6458 27292 8298
rect 27252 6452 27304 6458
rect 27252 6394 27304 6400
rect 26976 5840 27028 5846
rect 26976 5782 27028 5788
rect 26988 5642 27016 5782
rect 26976 5636 27028 5642
rect 26976 5578 27028 5584
rect 27252 5568 27304 5574
rect 27252 5510 27304 5516
rect 27158 5264 27214 5273
rect 27158 5199 27214 5208
rect 26884 5160 26936 5166
rect 26884 5102 26936 5108
rect 26976 5160 27028 5166
rect 26976 5102 27028 5108
rect 26884 3460 26936 3466
rect 26884 3402 26936 3408
rect 26700 3392 26752 3398
rect 26698 3360 26700 3369
rect 26792 3392 26844 3398
rect 26752 3360 26754 3369
rect 26792 3334 26844 3340
rect 26698 3295 26754 3304
rect 26896 3194 26924 3402
rect 26608 3188 26660 3194
rect 26608 3130 26660 3136
rect 26884 3188 26936 3194
rect 26884 3130 26936 3136
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 26424 2508 26476 2514
rect 26424 2450 26476 2456
rect 26332 1828 26384 1834
rect 26332 1770 26384 1776
rect 25780 1624 25832 1630
rect 25780 1566 25832 1572
rect 25778 1048 25834 1057
rect 25778 983 25834 992
rect 25792 800 25820 983
rect 26436 800 26464 2450
rect 26988 2378 27016 5102
rect 27068 4480 27120 4486
rect 27068 4422 27120 4428
rect 27080 4078 27108 4422
rect 27068 4072 27120 4078
rect 27068 4014 27120 4020
rect 27066 3632 27122 3641
rect 27066 3567 27122 3576
rect 26976 2372 27028 2378
rect 26976 2314 27028 2320
rect 27080 800 27108 3567
rect 27172 2990 27200 5199
rect 27264 3058 27292 5510
rect 27356 3194 27384 9998
rect 27448 8945 27476 10118
rect 27540 9042 27568 10406
rect 27724 9654 27752 12407
rect 27908 10810 27936 12650
rect 30840 12096 30892 12102
rect 30840 12038 30892 12044
rect 28080 11824 28132 11830
rect 28080 11766 28132 11772
rect 30288 11824 30340 11830
rect 30288 11766 30340 11772
rect 27986 11384 28042 11393
rect 27986 11319 28042 11328
rect 28000 11286 28028 11319
rect 27988 11280 28040 11286
rect 27988 11222 28040 11228
rect 27804 10804 27856 10810
rect 27804 10746 27856 10752
rect 27896 10804 27948 10810
rect 27896 10746 27948 10752
rect 27816 10674 27844 10746
rect 27988 10736 28040 10742
rect 27988 10678 28040 10684
rect 27804 10668 27856 10674
rect 27804 10610 27856 10616
rect 27804 10056 27856 10062
rect 28000 10033 28028 10678
rect 27804 9998 27856 10004
rect 27986 10024 28042 10033
rect 27816 9722 27844 9998
rect 27986 9959 28042 9968
rect 27804 9716 27856 9722
rect 27804 9658 27856 9664
rect 27712 9648 27764 9654
rect 27712 9590 27764 9596
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 27712 8968 27764 8974
rect 27434 8936 27490 8945
rect 27712 8910 27764 8916
rect 27434 8871 27436 8880
rect 27488 8871 27490 8880
rect 27436 8842 27488 8848
rect 27724 8809 27752 8910
rect 27710 8800 27766 8809
rect 27710 8735 27766 8744
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 27710 8392 27766 8401
rect 27710 8327 27766 8336
rect 27526 8256 27582 8265
rect 27526 8191 27582 8200
rect 27540 8090 27568 8191
rect 27528 8084 27580 8090
rect 27528 8026 27580 8032
rect 27618 7984 27674 7993
rect 27540 7942 27618 7970
rect 27540 7886 27568 7942
rect 27618 7919 27674 7928
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27434 7712 27490 7721
rect 27434 7647 27490 7656
rect 27448 7478 27476 7647
rect 27526 7576 27582 7585
rect 27632 7546 27660 7822
rect 27526 7511 27582 7520
rect 27620 7540 27672 7546
rect 27540 7478 27568 7511
rect 27620 7482 27672 7488
rect 27436 7472 27488 7478
rect 27436 7414 27488 7420
rect 27528 7472 27580 7478
rect 27528 7414 27580 7420
rect 27448 7002 27476 7414
rect 27436 6996 27488 7002
rect 27436 6938 27488 6944
rect 27528 6248 27580 6254
rect 27448 6208 27528 6236
rect 27448 6118 27476 6208
rect 27528 6190 27580 6196
rect 27436 6112 27488 6118
rect 27436 6054 27488 6060
rect 27448 5273 27476 6054
rect 27528 5908 27580 5914
rect 27528 5850 27580 5856
rect 27434 5264 27490 5273
rect 27434 5199 27490 5208
rect 27540 5098 27568 5850
rect 27724 5658 27752 8327
rect 27816 7886 27844 8434
rect 28092 8362 28120 11766
rect 29644 11756 29696 11762
rect 29644 11698 29696 11704
rect 28908 11688 28960 11694
rect 28908 11630 28960 11636
rect 28170 11520 28226 11529
rect 28170 11455 28226 11464
rect 28184 11150 28212 11455
rect 28540 11212 28592 11218
rect 28540 11154 28592 11160
rect 28724 11212 28776 11218
rect 28724 11154 28776 11160
rect 28172 11144 28224 11150
rect 28172 11086 28224 11092
rect 28264 11144 28316 11150
rect 28264 11086 28316 11092
rect 28170 10976 28226 10985
rect 28170 10911 28226 10920
rect 28184 10810 28212 10911
rect 28172 10804 28224 10810
rect 28172 10746 28224 10752
rect 28172 8424 28224 8430
rect 28172 8366 28224 8372
rect 27896 8356 27948 8362
rect 27896 8298 27948 8304
rect 28080 8356 28132 8362
rect 28080 8298 28132 8304
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 27804 7200 27856 7206
rect 27804 7142 27856 7148
rect 27632 5630 27752 5658
rect 27528 5092 27580 5098
rect 27528 5034 27580 5040
rect 27632 4706 27660 5630
rect 27710 5536 27766 5545
rect 27710 5471 27766 5480
rect 27448 4678 27660 4706
rect 27448 3942 27476 4678
rect 27528 4616 27580 4622
rect 27528 4558 27580 4564
rect 27620 4616 27672 4622
rect 27620 4558 27672 4564
rect 27436 3936 27488 3942
rect 27436 3878 27488 3884
rect 27344 3188 27396 3194
rect 27344 3130 27396 3136
rect 27342 3088 27398 3097
rect 27252 3052 27304 3058
rect 27342 3023 27344 3032
rect 27252 2994 27304 3000
rect 27396 3023 27398 3032
rect 27344 2994 27396 3000
rect 27160 2984 27212 2990
rect 27160 2926 27212 2932
rect 27540 2106 27568 4558
rect 27632 3602 27660 4558
rect 27620 3596 27672 3602
rect 27620 3538 27672 3544
rect 27528 2100 27580 2106
rect 27528 2042 27580 2048
rect 27724 800 27752 5471
rect 27816 3126 27844 7142
rect 27908 6458 27936 8298
rect 27988 7744 28040 7750
rect 27988 7686 28040 7692
rect 28000 6633 28028 7686
rect 28092 7562 28120 8298
rect 28184 7857 28212 8366
rect 28276 8022 28304 11086
rect 28552 10266 28580 11154
rect 28632 10464 28684 10470
rect 28630 10432 28632 10441
rect 28684 10432 28686 10441
rect 28630 10367 28686 10376
rect 28540 10260 28592 10266
rect 28540 10202 28592 10208
rect 28632 9920 28684 9926
rect 28632 9862 28684 9868
rect 28540 9648 28592 9654
rect 28540 9590 28592 9596
rect 28448 9444 28500 9450
rect 28448 9386 28500 9392
rect 28356 9376 28408 9382
rect 28356 9318 28408 9324
rect 28264 8016 28316 8022
rect 28264 7958 28316 7964
rect 28170 7848 28226 7857
rect 28170 7783 28226 7792
rect 28092 7534 28304 7562
rect 28172 7404 28224 7410
rect 28172 7346 28224 7352
rect 28078 7304 28134 7313
rect 28078 7239 28134 7248
rect 27986 6624 28042 6633
rect 27986 6559 28042 6568
rect 27896 6452 27948 6458
rect 27896 6394 27948 6400
rect 27896 5568 27948 5574
rect 27896 5510 27948 5516
rect 27804 3120 27856 3126
rect 27804 3062 27856 3068
rect 27908 2446 27936 5510
rect 27986 5264 28042 5273
rect 27986 5199 28042 5208
rect 28000 4214 28028 5199
rect 28092 4486 28120 7239
rect 28184 6934 28212 7346
rect 28172 6928 28224 6934
rect 28172 6870 28224 6876
rect 28276 6798 28304 7534
rect 28264 6792 28316 6798
rect 28264 6734 28316 6740
rect 28264 6656 28316 6662
rect 28264 6598 28316 6604
rect 28172 6384 28224 6390
rect 28172 6326 28224 6332
rect 28184 5302 28212 6326
rect 28276 6322 28304 6598
rect 28264 6316 28316 6322
rect 28264 6258 28316 6264
rect 28262 5944 28318 5953
rect 28262 5879 28318 5888
rect 28172 5296 28224 5302
rect 28172 5238 28224 5244
rect 28276 4842 28304 5879
rect 28184 4814 28304 4842
rect 28080 4480 28132 4486
rect 28080 4422 28132 4428
rect 27988 4208 28040 4214
rect 27988 4150 28040 4156
rect 28078 3632 28134 3641
rect 28078 3567 28134 3576
rect 27988 3392 28040 3398
rect 27988 3334 28040 3340
rect 28000 3058 28028 3334
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 28092 2990 28120 3567
rect 28184 3194 28212 4814
rect 28368 4690 28396 9318
rect 28460 9042 28488 9386
rect 28448 9036 28500 9042
rect 28448 8978 28500 8984
rect 28448 8832 28500 8838
rect 28552 8820 28580 9590
rect 28644 9518 28672 9862
rect 28632 9512 28684 9518
rect 28632 9454 28684 9460
rect 28644 9081 28672 9454
rect 28630 9072 28686 9081
rect 28630 9007 28686 9016
rect 28500 8792 28580 8820
rect 28448 8774 28500 8780
rect 28460 6866 28488 8774
rect 28630 7984 28686 7993
rect 28630 7919 28686 7928
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28552 7274 28580 7822
rect 28540 7268 28592 7274
rect 28540 7210 28592 7216
rect 28644 6866 28672 7919
rect 28736 7410 28764 11154
rect 28814 10840 28870 10849
rect 28814 10775 28870 10784
rect 28828 10674 28856 10775
rect 28816 10668 28868 10674
rect 28816 10610 28868 10616
rect 28816 10464 28868 10470
rect 28816 10406 28868 10412
rect 28828 7954 28856 10406
rect 28816 7948 28868 7954
rect 28816 7890 28868 7896
rect 28724 7404 28776 7410
rect 28724 7346 28776 7352
rect 28448 6860 28500 6866
rect 28448 6802 28500 6808
rect 28632 6860 28684 6866
rect 28632 6802 28684 6808
rect 28540 6792 28592 6798
rect 28540 6734 28592 6740
rect 28446 6216 28502 6225
rect 28446 6151 28502 6160
rect 28264 4684 28316 4690
rect 28264 4626 28316 4632
rect 28356 4684 28408 4690
rect 28356 4626 28408 4632
rect 28276 4214 28304 4626
rect 28460 4486 28488 6151
rect 28448 4480 28500 4486
rect 28368 4428 28448 4434
rect 28368 4422 28500 4428
rect 28368 4406 28488 4422
rect 28264 4208 28316 4214
rect 28264 4150 28316 4156
rect 28276 3194 28304 4150
rect 28368 3738 28396 4406
rect 28446 4312 28502 4321
rect 28446 4247 28502 4256
rect 28460 4146 28488 4247
rect 28448 4140 28500 4146
rect 28448 4082 28500 4088
rect 28356 3732 28408 3738
rect 28356 3674 28408 3680
rect 28356 3596 28408 3602
rect 28356 3538 28408 3544
rect 28172 3188 28224 3194
rect 28172 3130 28224 3136
rect 28264 3188 28316 3194
rect 28264 3130 28316 3136
rect 28080 2984 28132 2990
rect 28080 2926 28132 2932
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 28080 2304 28132 2310
rect 28080 2246 28132 2252
rect 28092 1873 28120 2246
rect 28078 1864 28134 1873
rect 28078 1799 28134 1808
rect 28368 800 28396 3538
rect 28552 3466 28580 6734
rect 28644 6497 28672 6802
rect 28630 6488 28686 6497
rect 28920 6458 28948 11630
rect 29000 11620 29052 11626
rect 29000 11562 29052 11568
rect 29012 11354 29040 11562
rect 29276 11552 29328 11558
rect 29276 11494 29328 11500
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29184 11076 29236 11082
rect 29184 11018 29236 11024
rect 29000 10600 29052 10606
rect 29000 10542 29052 10548
rect 29012 9926 29040 10542
rect 29196 10441 29224 11018
rect 29182 10432 29238 10441
rect 29182 10367 29238 10376
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 29012 9625 29040 9862
rect 28998 9616 29054 9625
rect 28998 9551 29054 9560
rect 29000 9444 29052 9450
rect 29000 9386 29052 9392
rect 29092 9444 29144 9450
rect 29092 9386 29144 9392
rect 29012 8906 29040 9386
rect 29000 8900 29052 8906
rect 29000 8842 29052 8848
rect 29104 7954 29132 9386
rect 29184 9376 29236 9382
rect 29184 9318 29236 9324
rect 29196 8809 29224 9318
rect 29288 9042 29316 11494
rect 29656 11014 29684 11698
rect 29828 11144 29880 11150
rect 29828 11086 29880 11092
rect 29644 11008 29696 11014
rect 29644 10950 29696 10956
rect 29656 10810 29684 10950
rect 29644 10804 29696 10810
rect 29644 10746 29696 10752
rect 29736 10600 29788 10606
rect 29736 10542 29788 10548
rect 29460 10056 29512 10062
rect 29460 9998 29512 10004
rect 29276 9036 29328 9042
rect 29276 8978 29328 8984
rect 29368 8832 29420 8838
rect 29182 8800 29238 8809
rect 29368 8774 29420 8780
rect 29182 8735 29238 8744
rect 29092 7948 29144 7954
rect 29092 7890 29144 7896
rect 29092 7744 29144 7750
rect 29092 7686 29144 7692
rect 29000 6656 29052 6662
rect 29000 6598 29052 6604
rect 28630 6423 28686 6432
rect 28908 6452 28960 6458
rect 28908 6394 28960 6400
rect 28816 6248 28868 6254
rect 28816 6190 28868 6196
rect 28828 5370 28856 6190
rect 28816 5364 28868 5370
rect 28816 5306 28868 5312
rect 28724 5228 28776 5234
rect 28724 5170 28776 5176
rect 28736 3738 28764 5170
rect 29012 5166 29040 6598
rect 29104 5817 29132 7686
rect 29090 5808 29146 5817
rect 29090 5743 29146 5752
rect 29196 5702 29224 8735
rect 29104 5674 29224 5702
rect 29000 5160 29052 5166
rect 29000 5102 29052 5108
rect 28998 4992 29054 5001
rect 28998 4927 29054 4936
rect 28906 4856 28962 4865
rect 28906 4791 28962 4800
rect 28920 4690 28948 4791
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 28816 4548 28868 4554
rect 28816 4490 28868 4496
rect 28828 4282 28856 4490
rect 28816 4276 28868 4282
rect 28816 4218 28868 4224
rect 28724 3732 28776 3738
rect 28724 3674 28776 3680
rect 28540 3460 28592 3466
rect 28540 3402 28592 3408
rect 28552 3058 28580 3402
rect 28722 3224 28778 3233
rect 28722 3159 28778 3168
rect 28736 3126 28764 3159
rect 28724 3120 28776 3126
rect 28724 3062 28776 3068
rect 28540 3052 28592 3058
rect 28540 2994 28592 3000
rect 28814 2408 28870 2417
rect 28814 2343 28816 2352
rect 28868 2343 28870 2352
rect 28816 2314 28868 2320
rect 29012 800 29040 4927
rect 29104 4690 29132 5674
rect 29184 5568 29236 5574
rect 29184 5510 29236 5516
rect 29092 4684 29144 4690
rect 29092 4626 29144 4632
rect 29092 4072 29144 4078
rect 29092 4014 29144 4020
rect 29104 3534 29132 4014
rect 29196 4010 29224 5510
rect 29274 5400 29330 5409
rect 29274 5335 29330 5344
rect 29288 5234 29316 5335
rect 29276 5228 29328 5234
rect 29276 5170 29328 5176
rect 29380 5098 29408 8774
rect 29368 5092 29420 5098
rect 29368 5034 29420 5040
rect 29276 4684 29328 4690
rect 29276 4626 29328 4632
rect 29184 4004 29236 4010
rect 29184 3946 29236 3952
rect 29092 3528 29144 3534
rect 29092 3470 29144 3476
rect 29288 2990 29316 4626
rect 29472 4010 29500 9998
rect 29552 9988 29604 9994
rect 29552 9930 29604 9936
rect 29564 8022 29592 9930
rect 29644 9512 29696 9518
rect 29644 9454 29696 9460
rect 29656 9081 29684 9454
rect 29642 9072 29698 9081
rect 29642 9007 29698 9016
rect 29644 8968 29696 8974
rect 29644 8910 29696 8916
rect 29656 8634 29684 8910
rect 29644 8628 29696 8634
rect 29644 8570 29696 8576
rect 29644 8424 29696 8430
rect 29644 8366 29696 8372
rect 29552 8016 29604 8022
rect 29552 7958 29604 7964
rect 29552 7812 29604 7818
rect 29552 7754 29604 7760
rect 29564 7449 29592 7754
rect 29656 7478 29684 8366
rect 29644 7472 29696 7478
rect 29550 7440 29606 7449
rect 29644 7414 29696 7420
rect 29550 7375 29606 7384
rect 29642 5536 29698 5545
rect 29642 5471 29698 5480
rect 29552 5160 29604 5166
rect 29550 5128 29552 5137
rect 29604 5128 29606 5137
rect 29550 5063 29606 5072
rect 29656 4078 29684 5471
rect 29644 4072 29696 4078
rect 29644 4014 29696 4020
rect 29460 4004 29512 4010
rect 29460 3946 29512 3952
rect 29276 2984 29328 2990
rect 29276 2926 29328 2932
rect 29748 2774 29776 10542
rect 29840 7546 29868 11086
rect 30300 10674 30328 11766
rect 30380 11280 30432 11286
rect 30380 11222 30432 11228
rect 30288 10668 30340 10674
rect 30288 10610 30340 10616
rect 30196 10464 30248 10470
rect 30196 10406 30248 10412
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 29920 8424 29972 8430
rect 29920 8366 29972 8372
rect 29932 8090 29960 8366
rect 29920 8084 29972 8090
rect 29920 8026 29972 8032
rect 29920 7812 29972 7818
rect 29920 7754 29972 7760
rect 29828 7540 29880 7546
rect 29828 7482 29880 7488
rect 29932 6866 29960 7754
rect 29920 6860 29972 6866
rect 29920 6802 29972 6808
rect 29920 6656 29972 6662
rect 29920 6598 29972 6604
rect 29828 6248 29880 6254
rect 29828 6190 29880 6196
rect 29840 4826 29868 6190
rect 29828 4820 29880 4826
rect 29828 4762 29880 4768
rect 29932 2854 29960 6598
rect 30024 3126 30052 9862
rect 30208 9761 30236 10406
rect 30300 10266 30328 10610
rect 30288 10260 30340 10266
rect 30288 10202 30340 10208
rect 30194 9752 30250 9761
rect 30194 9687 30250 9696
rect 30196 8628 30248 8634
rect 30196 8570 30248 8576
rect 30208 8537 30236 8570
rect 30194 8528 30250 8537
rect 30194 8463 30250 8472
rect 30196 8016 30248 8022
rect 30196 7958 30248 7964
rect 30208 7750 30236 7958
rect 30300 7750 30328 10202
rect 30392 8090 30420 11222
rect 30472 9920 30524 9926
rect 30472 9862 30524 9868
rect 30484 9042 30512 9862
rect 30656 9648 30708 9654
rect 30656 9590 30708 9596
rect 30562 9480 30618 9489
rect 30562 9415 30618 9424
rect 30472 9036 30524 9042
rect 30472 8978 30524 8984
rect 30472 8900 30524 8906
rect 30472 8842 30524 8848
rect 30380 8084 30432 8090
rect 30380 8026 30432 8032
rect 30196 7744 30248 7750
rect 30196 7686 30248 7692
rect 30288 7744 30340 7750
rect 30288 7686 30340 7692
rect 30196 7540 30248 7546
rect 30196 7482 30248 7488
rect 30102 7304 30158 7313
rect 30208 7290 30236 7482
rect 30288 7472 30340 7478
rect 30340 7432 30420 7460
rect 30288 7414 30340 7420
rect 30208 7262 30328 7290
rect 30102 7239 30158 7248
rect 30116 6866 30144 7239
rect 30196 7200 30248 7206
rect 30196 7142 30248 7148
rect 30104 6860 30156 6866
rect 30104 6802 30156 6808
rect 30116 6769 30144 6802
rect 30102 6760 30158 6769
rect 30102 6695 30158 6704
rect 30102 6624 30158 6633
rect 30102 6559 30158 6568
rect 30116 6322 30144 6559
rect 30104 6316 30156 6322
rect 30104 6258 30156 6264
rect 30104 5704 30156 5710
rect 30104 5646 30156 5652
rect 30012 3120 30064 3126
rect 30012 3062 30064 3068
rect 29920 2848 29972 2854
rect 29920 2790 29972 2796
rect 29656 2746 29776 2774
rect 29656 800 29684 2746
rect 30116 2446 30144 5646
rect 30208 5574 30236 7142
rect 30300 6458 30328 7262
rect 30392 6458 30420 7432
rect 30484 6882 30512 8842
rect 30576 7002 30604 9415
rect 30668 8430 30696 9590
rect 30748 9376 30800 9382
rect 30748 9318 30800 9324
rect 30656 8424 30708 8430
rect 30656 8366 30708 8372
rect 30668 8129 30696 8366
rect 30654 8120 30710 8129
rect 30654 8055 30710 8064
rect 30656 7880 30708 7886
rect 30654 7848 30656 7857
rect 30708 7848 30710 7857
rect 30654 7783 30710 7792
rect 30654 7032 30710 7041
rect 30564 6996 30616 7002
rect 30654 6967 30710 6976
rect 30564 6938 30616 6944
rect 30484 6854 30604 6882
rect 30668 6866 30696 6967
rect 30576 6746 30604 6854
rect 30656 6860 30708 6866
rect 30656 6802 30708 6808
rect 30472 6724 30524 6730
rect 30576 6718 30696 6746
rect 30472 6666 30524 6672
rect 30288 6452 30340 6458
rect 30288 6394 30340 6400
rect 30380 6452 30432 6458
rect 30380 6394 30432 6400
rect 30196 5568 30248 5574
rect 30196 5510 30248 5516
rect 30392 5234 30420 6394
rect 30484 6322 30512 6666
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30472 6180 30524 6186
rect 30472 6122 30524 6128
rect 30380 5228 30432 5234
rect 30380 5170 30432 5176
rect 30196 5024 30248 5030
rect 30196 4966 30248 4972
rect 30208 3466 30236 4966
rect 30288 4480 30340 4486
rect 30288 4422 30340 4428
rect 30300 3738 30328 4422
rect 30288 3732 30340 3738
rect 30288 3674 30340 3680
rect 30392 3602 30420 5170
rect 30484 4622 30512 6122
rect 30562 5672 30618 5681
rect 30562 5607 30618 5616
rect 30576 5030 30604 5607
rect 30668 5574 30696 6718
rect 30656 5568 30708 5574
rect 30656 5510 30708 5516
rect 30564 5024 30616 5030
rect 30564 4966 30616 4972
rect 30472 4616 30524 4622
rect 30472 4558 30524 4564
rect 30668 4468 30696 5510
rect 30484 4440 30696 4468
rect 30380 3596 30432 3602
rect 30380 3538 30432 3544
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 30196 3460 30248 3466
rect 30196 3402 30248 3408
rect 30300 3074 30328 3470
rect 30380 3460 30432 3466
rect 30380 3402 30432 3408
rect 30392 3176 30420 3402
rect 30484 3398 30512 4440
rect 30656 4276 30708 4282
rect 30656 4218 30708 4224
rect 30564 3460 30616 3466
rect 30564 3402 30616 3408
rect 30472 3392 30524 3398
rect 30472 3334 30524 3340
rect 30472 3188 30524 3194
rect 30392 3148 30472 3176
rect 30472 3130 30524 3136
rect 30300 3046 30512 3074
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30288 2508 30340 2514
rect 30288 2450 30340 2456
rect 30104 2440 30156 2446
rect 30104 2382 30156 2388
rect 30300 800 30328 2450
rect 30392 2446 30420 2790
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 30484 1970 30512 3046
rect 30576 2854 30604 3402
rect 30668 3398 30696 4218
rect 30760 3534 30788 9318
rect 30852 8022 30880 12038
rect 31300 10804 31352 10810
rect 31300 10746 31352 10752
rect 31208 10736 31260 10742
rect 31206 10704 31208 10713
rect 31260 10704 31262 10713
rect 31206 10639 31262 10648
rect 31206 10160 31262 10169
rect 31206 10095 31208 10104
rect 31260 10095 31262 10104
rect 31208 10066 31260 10072
rect 31312 9674 31340 10746
rect 31496 10606 31524 16546
rect 31588 16546 31708 16574
rect 31484 10600 31536 10606
rect 31484 10542 31536 10548
rect 31036 9646 31340 9674
rect 31588 9654 31616 16546
rect 36514 16348 36822 16357
rect 36514 16346 36520 16348
rect 36576 16346 36600 16348
rect 36656 16346 36680 16348
rect 36736 16346 36760 16348
rect 36816 16346 36822 16348
rect 36576 16294 36578 16346
rect 36758 16294 36760 16346
rect 36514 16292 36520 16294
rect 36576 16292 36600 16294
rect 36656 16292 36680 16294
rect 36736 16292 36760 16294
rect 36816 16292 36822 16294
rect 36514 16283 36822 16292
rect 35854 15804 36162 15813
rect 35854 15802 35860 15804
rect 35916 15802 35940 15804
rect 35996 15802 36020 15804
rect 36076 15802 36100 15804
rect 36156 15802 36162 15804
rect 35916 15750 35918 15802
rect 36098 15750 36100 15802
rect 35854 15748 35860 15750
rect 35916 15748 35940 15750
rect 35996 15748 36020 15750
rect 36076 15748 36100 15750
rect 36156 15748 36162 15750
rect 35854 15739 36162 15748
rect 36514 15260 36822 15269
rect 36514 15258 36520 15260
rect 36576 15258 36600 15260
rect 36656 15258 36680 15260
rect 36736 15258 36760 15260
rect 36816 15258 36822 15260
rect 36576 15206 36578 15258
rect 36758 15206 36760 15258
rect 36514 15204 36520 15206
rect 36576 15204 36600 15206
rect 36656 15204 36680 15206
rect 36736 15204 36760 15206
rect 36816 15204 36822 15206
rect 36514 15195 36822 15204
rect 35854 14716 36162 14725
rect 35854 14714 35860 14716
rect 35916 14714 35940 14716
rect 35996 14714 36020 14716
rect 36076 14714 36100 14716
rect 36156 14714 36162 14716
rect 35916 14662 35918 14714
rect 36098 14662 36100 14714
rect 35854 14660 35860 14662
rect 35916 14660 35940 14662
rect 35996 14660 36020 14662
rect 36076 14660 36100 14662
rect 36156 14660 36162 14662
rect 35854 14651 36162 14660
rect 39132 14521 39160 37198
rect 40880 36922 40908 37198
rect 42720 37194 42748 39200
rect 43352 37256 43404 37262
rect 43352 37198 43404 37204
rect 42708 37188 42760 37194
rect 42708 37130 42760 37136
rect 40868 36916 40920 36922
rect 40868 36858 40920 36864
rect 43364 32434 43392 37198
rect 44560 36666 44588 39200
rect 46400 37194 46428 39200
rect 48240 37346 48268 39200
rect 48148 37318 48268 37346
rect 46480 37256 46532 37262
rect 46480 37198 46532 37204
rect 46388 37188 46440 37194
rect 46388 37130 46440 37136
rect 44732 36712 44784 36718
rect 44560 36660 44732 36666
rect 44560 36654 44784 36660
rect 44560 36638 44772 36654
rect 43352 32428 43404 32434
rect 43352 32370 43404 32376
rect 46492 24138 46520 37198
rect 48148 37194 48176 37318
rect 48228 37256 48280 37262
rect 48228 37198 48280 37204
rect 48136 37188 48188 37194
rect 48136 37130 48188 37136
rect 48240 36922 48268 37198
rect 48228 36916 48280 36922
rect 48228 36858 48280 36864
rect 50080 36718 50108 39200
rect 51920 37618 51948 39200
rect 51920 37590 52132 37618
rect 52104 37262 52132 37590
rect 51908 37256 51960 37262
rect 51908 37198 51960 37204
rect 52092 37256 52144 37262
rect 52092 37198 52144 37204
rect 51920 36922 51948 37198
rect 53760 37194 53788 39200
rect 55600 37346 55628 39200
rect 55600 37318 55720 37346
rect 53840 37256 53892 37262
rect 53840 37198 53892 37204
rect 55588 37256 55640 37262
rect 55588 37198 55640 37204
rect 53748 37188 53800 37194
rect 53748 37130 53800 37136
rect 51908 36916 51960 36922
rect 51908 36858 51960 36864
rect 50160 36780 50212 36786
rect 50160 36722 50212 36728
rect 50068 36712 50120 36718
rect 50068 36654 50120 36660
rect 50172 29646 50200 36722
rect 50160 29640 50212 29646
rect 50160 29582 50212 29588
rect 53852 26926 53880 37198
rect 55600 36922 55628 37198
rect 55692 37194 55720 37318
rect 57440 37194 57468 39200
rect 58808 37256 58860 37262
rect 58808 37198 58860 37204
rect 55680 37188 55732 37194
rect 55680 37130 55732 37136
rect 57428 37188 57480 37194
rect 57428 37130 57480 37136
rect 55588 36916 55640 36922
rect 55588 36858 55640 36864
rect 53840 26920 53892 26926
rect 53840 26862 53892 26868
rect 46480 24132 46532 24138
rect 46480 24074 46532 24080
rect 39118 14512 39174 14521
rect 58820 14482 58848 37198
rect 59280 36854 59308 39200
rect 66574 37564 66882 37573
rect 66574 37562 66580 37564
rect 66636 37562 66660 37564
rect 66716 37562 66740 37564
rect 66796 37562 66820 37564
rect 66876 37562 66882 37564
rect 66636 37510 66638 37562
rect 66818 37510 66820 37562
rect 66574 37508 66580 37510
rect 66636 37508 66660 37510
rect 66716 37508 66740 37510
rect 66796 37508 66820 37510
rect 66876 37508 66882 37510
rect 66574 37499 66882 37508
rect 67234 37020 67542 37029
rect 67234 37018 67240 37020
rect 67296 37018 67320 37020
rect 67376 37018 67400 37020
rect 67456 37018 67480 37020
rect 67536 37018 67542 37020
rect 67296 36966 67298 37018
rect 67478 36966 67480 37018
rect 67234 36964 67240 36966
rect 67296 36964 67320 36966
rect 67376 36964 67400 36966
rect 67456 36964 67480 36966
rect 67536 36964 67542 36966
rect 67234 36955 67542 36964
rect 59268 36848 59320 36854
rect 59268 36790 59320 36796
rect 66574 36476 66882 36485
rect 66574 36474 66580 36476
rect 66636 36474 66660 36476
rect 66716 36474 66740 36476
rect 66796 36474 66820 36476
rect 66876 36474 66882 36476
rect 66636 36422 66638 36474
rect 66818 36422 66820 36474
rect 66574 36420 66580 36422
rect 66636 36420 66660 36422
rect 66716 36420 66740 36422
rect 66796 36420 66820 36422
rect 66876 36420 66882 36422
rect 66574 36411 66882 36420
rect 67234 35932 67542 35941
rect 67234 35930 67240 35932
rect 67296 35930 67320 35932
rect 67376 35930 67400 35932
rect 67456 35930 67480 35932
rect 67536 35930 67542 35932
rect 67296 35878 67298 35930
rect 67478 35878 67480 35930
rect 67234 35876 67240 35878
rect 67296 35876 67320 35878
rect 67376 35876 67400 35878
rect 67456 35876 67480 35878
rect 67536 35876 67542 35878
rect 67234 35867 67542 35876
rect 66574 35388 66882 35397
rect 66574 35386 66580 35388
rect 66636 35386 66660 35388
rect 66716 35386 66740 35388
rect 66796 35386 66820 35388
rect 66876 35386 66882 35388
rect 66636 35334 66638 35386
rect 66818 35334 66820 35386
rect 66574 35332 66580 35334
rect 66636 35332 66660 35334
rect 66716 35332 66740 35334
rect 66796 35332 66820 35334
rect 66876 35332 66882 35334
rect 66574 35323 66882 35332
rect 67234 34844 67542 34853
rect 67234 34842 67240 34844
rect 67296 34842 67320 34844
rect 67376 34842 67400 34844
rect 67456 34842 67480 34844
rect 67536 34842 67542 34844
rect 67296 34790 67298 34842
rect 67478 34790 67480 34842
rect 67234 34788 67240 34790
rect 67296 34788 67320 34790
rect 67376 34788 67400 34790
rect 67456 34788 67480 34790
rect 67536 34788 67542 34790
rect 67234 34779 67542 34788
rect 66574 34300 66882 34309
rect 66574 34298 66580 34300
rect 66636 34298 66660 34300
rect 66716 34298 66740 34300
rect 66796 34298 66820 34300
rect 66876 34298 66882 34300
rect 66636 34246 66638 34298
rect 66818 34246 66820 34298
rect 66574 34244 66580 34246
rect 66636 34244 66660 34246
rect 66716 34244 66740 34246
rect 66796 34244 66820 34246
rect 66876 34244 66882 34246
rect 66574 34235 66882 34244
rect 67234 33756 67542 33765
rect 67234 33754 67240 33756
rect 67296 33754 67320 33756
rect 67376 33754 67400 33756
rect 67456 33754 67480 33756
rect 67536 33754 67542 33756
rect 67296 33702 67298 33754
rect 67478 33702 67480 33754
rect 67234 33700 67240 33702
rect 67296 33700 67320 33702
rect 67376 33700 67400 33702
rect 67456 33700 67480 33702
rect 67536 33700 67542 33702
rect 67234 33691 67542 33700
rect 66574 33212 66882 33221
rect 66574 33210 66580 33212
rect 66636 33210 66660 33212
rect 66716 33210 66740 33212
rect 66796 33210 66820 33212
rect 66876 33210 66882 33212
rect 66636 33158 66638 33210
rect 66818 33158 66820 33210
rect 66574 33156 66580 33158
rect 66636 33156 66660 33158
rect 66716 33156 66740 33158
rect 66796 33156 66820 33158
rect 66876 33156 66882 33158
rect 66574 33147 66882 33156
rect 67234 32668 67542 32677
rect 67234 32666 67240 32668
rect 67296 32666 67320 32668
rect 67376 32666 67400 32668
rect 67456 32666 67480 32668
rect 67536 32666 67542 32668
rect 67296 32614 67298 32666
rect 67478 32614 67480 32666
rect 67234 32612 67240 32614
rect 67296 32612 67320 32614
rect 67376 32612 67400 32614
rect 67456 32612 67480 32614
rect 67536 32612 67542 32614
rect 67234 32603 67542 32612
rect 66574 32124 66882 32133
rect 66574 32122 66580 32124
rect 66636 32122 66660 32124
rect 66716 32122 66740 32124
rect 66796 32122 66820 32124
rect 66876 32122 66882 32124
rect 66636 32070 66638 32122
rect 66818 32070 66820 32122
rect 66574 32068 66580 32070
rect 66636 32068 66660 32070
rect 66716 32068 66740 32070
rect 66796 32068 66820 32070
rect 66876 32068 66882 32070
rect 66574 32059 66882 32068
rect 67234 31580 67542 31589
rect 67234 31578 67240 31580
rect 67296 31578 67320 31580
rect 67376 31578 67400 31580
rect 67456 31578 67480 31580
rect 67536 31578 67542 31580
rect 67296 31526 67298 31578
rect 67478 31526 67480 31578
rect 67234 31524 67240 31526
rect 67296 31524 67320 31526
rect 67376 31524 67400 31526
rect 67456 31524 67480 31526
rect 67536 31524 67542 31526
rect 67234 31515 67542 31524
rect 66574 31036 66882 31045
rect 66574 31034 66580 31036
rect 66636 31034 66660 31036
rect 66716 31034 66740 31036
rect 66796 31034 66820 31036
rect 66876 31034 66882 31036
rect 66636 30982 66638 31034
rect 66818 30982 66820 31034
rect 66574 30980 66580 30982
rect 66636 30980 66660 30982
rect 66716 30980 66740 30982
rect 66796 30980 66820 30982
rect 66876 30980 66882 30982
rect 66574 30971 66882 30980
rect 67234 30492 67542 30501
rect 67234 30490 67240 30492
rect 67296 30490 67320 30492
rect 67376 30490 67400 30492
rect 67456 30490 67480 30492
rect 67536 30490 67542 30492
rect 67296 30438 67298 30490
rect 67478 30438 67480 30490
rect 67234 30436 67240 30438
rect 67296 30436 67320 30438
rect 67376 30436 67400 30438
rect 67456 30436 67480 30438
rect 67536 30436 67542 30438
rect 67234 30427 67542 30436
rect 66574 29948 66882 29957
rect 66574 29946 66580 29948
rect 66636 29946 66660 29948
rect 66716 29946 66740 29948
rect 66796 29946 66820 29948
rect 66876 29946 66882 29948
rect 66636 29894 66638 29946
rect 66818 29894 66820 29946
rect 66574 29892 66580 29894
rect 66636 29892 66660 29894
rect 66716 29892 66740 29894
rect 66796 29892 66820 29894
rect 66876 29892 66882 29894
rect 66574 29883 66882 29892
rect 67234 29404 67542 29413
rect 67234 29402 67240 29404
rect 67296 29402 67320 29404
rect 67376 29402 67400 29404
rect 67456 29402 67480 29404
rect 67536 29402 67542 29404
rect 67296 29350 67298 29402
rect 67478 29350 67480 29402
rect 67234 29348 67240 29350
rect 67296 29348 67320 29350
rect 67376 29348 67400 29350
rect 67456 29348 67480 29350
rect 67536 29348 67542 29350
rect 67234 29339 67542 29348
rect 66574 28860 66882 28869
rect 66574 28858 66580 28860
rect 66636 28858 66660 28860
rect 66716 28858 66740 28860
rect 66796 28858 66820 28860
rect 66876 28858 66882 28860
rect 66636 28806 66638 28858
rect 66818 28806 66820 28858
rect 66574 28804 66580 28806
rect 66636 28804 66660 28806
rect 66716 28804 66740 28806
rect 66796 28804 66820 28806
rect 66876 28804 66882 28806
rect 66574 28795 66882 28804
rect 67234 28316 67542 28325
rect 67234 28314 67240 28316
rect 67296 28314 67320 28316
rect 67376 28314 67400 28316
rect 67456 28314 67480 28316
rect 67536 28314 67542 28316
rect 67296 28262 67298 28314
rect 67478 28262 67480 28314
rect 67234 28260 67240 28262
rect 67296 28260 67320 28262
rect 67376 28260 67400 28262
rect 67456 28260 67480 28262
rect 67536 28260 67542 28262
rect 67234 28251 67542 28260
rect 66574 27772 66882 27781
rect 66574 27770 66580 27772
rect 66636 27770 66660 27772
rect 66716 27770 66740 27772
rect 66796 27770 66820 27772
rect 66876 27770 66882 27772
rect 66636 27718 66638 27770
rect 66818 27718 66820 27770
rect 66574 27716 66580 27718
rect 66636 27716 66660 27718
rect 66716 27716 66740 27718
rect 66796 27716 66820 27718
rect 66876 27716 66882 27718
rect 66574 27707 66882 27716
rect 67234 27228 67542 27237
rect 67234 27226 67240 27228
rect 67296 27226 67320 27228
rect 67376 27226 67400 27228
rect 67456 27226 67480 27228
rect 67536 27226 67542 27228
rect 67296 27174 67298 27226
rect 67478 27174 67480 27226
rect 67234 27172 67240 27174
rect 67296 27172 67320 27174
rect 67376 27172 67400 27174
rect 67456 27172 67480 27174
rect 67536 27172 67542 27174
rect 67234 27163 67542 27172
rect 66574 26684 66882 26693
rect 66574 26682 66580 26684
rect 66636 26682 66660 26684
rect 66716 26682 66740 26684
rect 66796 26682 66820 26684
rect 66876 26682 66882 26684
rect 66636 26630 66638 26682
rect 66818 26630 66820 26682
rect 66574 26628 66580 26630
rect 66636 26628 66660 26630
rect 66716 26628 66740 26630
rect 66796 26628 66820 26630
rect 66876 26628 66882 26630
rect 66574 26619 66882 26628
rect 67234 26140 67542 26149
rect 67234 26138 67240 26140
rect 67296 26138 67320 26140
rect 67376 26138 67400 26140
rect 67456 26138 67480 26140
rect 67536 26138 67542 26140
rect 67296 26086 67298 26138
rect 67478 26086 67480 26138
rect 67234 26084 67240 26086
rect 67296 26084 67320 26086
rect 67376 26084 67400 26086
rect 67456 26084 67480 26086
rect 67536 26084 67542 26086
rect 67234 26075 67542 26084
rect 66574 25596 66882 25605
rect 66574 25594 66580 25596
rect 66636 25594 66660 25596
rect 66716 25594 66740 25596
rect 66796 25594 66820 25596
rect 66876 25594 66882 25596
rect 66636 25542 66638 25594
rect 66818 25542 66820 25594
rect 66574 25540 66580 25542
rect 66636 25540 66660 25542
rect 66716 25540 66740 25542
rect 66796 25540 66820 25542
rect 66876 25540 66882 25542
rect 66574 25531 66882 25540
rect 67234 25052 67542 25061
rect 67234 25050 67240 25052
rect 67296 25050 67320 25052
rect 67376 25050 67400 25052
rect 67456 25050 67480 25052
rect 67536 25050 67542 25052
rect 67296 24998 67298 25050
rect 67478 24998 67480 25050
rect 67234 24996 67240 24998
rect 67296 24996 67320 24998
rect 67376 24996 67400 24998
rect 67456 24996 67480 24998
rect 67536 24996 67542 24998
rect 67234 24987 67542 24996
rect 66574 24508 66882 24517
rect 66574 24506 66580 24508
rect 66636 24506 66660 24508
rect 66716 24506 66740 24508
rect 66796 24506 66820 24508
rect 66876 24506 66882 24508
rect 66636 24454 66638 24506
rect 66818 24454 66820 24506
rect 66574 24452 66580 24454
rect 66636 24452 66660 24454
rect 66716 24452 66740 24454
rect 66796 24452 66820 24454
rect 66876 24452 66882 24454
rect 66574 24443 66882 24452
rect 67234 23964 67542 23973
rect 67234 23962 67240 23964
rect 67296 23962 67320 23964
rect 67376 23962 67400 23964
rect 67456 23962 67480 23964
rect 67536 23962 67542 23964
rect 67296 23910 67298 23962
rect 67478 23910 67480 23962
rect 67234 23908 67240 23910
rect 67296 23908 67320 23910
rect 67376 23908 67400 23910
rect 67456 23908 67480 23910
rect 67536 23908 67542 23910
rect 67234 23899 67542 23908
rect 66574 23420 66882 23429
rect 66574 23418 66580 23420
rect 66636 23418 66660 23420
rect 66716 23418 66740 23420
rect 66796 23418 66820 23420
rect 66876 23418 66882 23420
rect 66636 23366 66638 23418
rect 66818 23366 66820 23418
rect 66574 23364 66580 23366
rect 66636 23364 66660 23366
rect 66716 23364 66740 23366
rect 66796 23364 66820 23366
rect 66876 23364 66882 23366
rect 66574 23355 66882 23364
rect 67234 22876 67542 22885
rect 67234 22874 67240 22876
rect 67296 22874 67320 22876
rect 67376 22874 67400 22876
rect 67456 22874 67480 22876
rect 67536 22874 67542 22876
rect 67296 22822 67298 22874
rect 67478 22822 67480 22874
rect 67234 22820 67240 22822
rect 67296 22820 67320 22822
rect 67376 22820 67400 22822
rect 67456 22820 67480 22822
rect 67536 22820 67542 22822
rect 67234 22811 67542 22820
rect 66574 22332 66882 22341
rect 66574 22330 66580 22332
rect 66636 22330 66660 22332
rect 66716 22330 66740 22332
rect 66796 22330 66820 22332
rect 66876 22330 66882 22332
rect 66636 22278 66638 22330
rect 66818 22278 66820 22330
rect 66574 22276 66580 22278
rect 66636 22276 66660 22278
rect 66716 22276 66740 22278
rect 66796 22276 66820 22278
rect 66876 22276 66882 22278
rect 66574 22267 66882 22276
rect 67234 21788 67542 21797
rect 67234 21786 67240 21788
rect 67296 21786 67320 21788
rect 67376 21786 67400 21788
rect 67456 21786 67480 21788
rect 67536 21786 67542 21788
rect 67296 21734 67298 21786
rect 67478 21734 67480 21786
rect 67234 21732 67240 21734
rect 67296 21732 67320 21734
rect 67376 21732 67400 21734
rect 67456 21732 67480 21734
rect 67536 21732 67542 21734
rect 67234 21723 67542 21732
rect 66574 21244 66882 21253
rect 66574 21242 66580 21244
rect 66636 21242 66660 21244
rect 66716 21242 66740 21244
rect 66796 21242 66820 21244
rect 66876 21242 66882 21244
rect 66636 21190 66638 21242
rect 66818 21190 66820 21242
rect 66574 21188 66580 21190
rect 66636 21188 66660 21190
rect 66716 21188 66740 21190
rect 66796 21188 66820 21190
rect 66876 21188 66882 21190
rect 66574 21179 66882 21188
rect 67234 20700 67542 20709
rect 67234 20698 67240 20700
rect 67296 20698 67320 20700
rect 67376 20698 67400 20700
rect 67456 20698 67480 20700
rect 67536 20698 67542 20700
rect 67296 20646 67298 20698
rect 67478 20646 67480 20698
rect 67234 20644 67240 20646
rect 67296 20644 67320 20646
rect 67376 20644 67400 20646
rect 67456 20644 67480 20646
rect 67536 20644 67542 20646
rect 67234 20635 67542 20644
rect 66574 20156 66882 20165
rect 66574 20154 66580 20156
rect 66636 20154 66660 20156
rect 66716 20154 66740 20156
rect 66796 20154 66820 20156
rect 66876 20154 66882 20156
rect 66636 20102 66638 20154
rect 66818 20102 66820 20154
rect 66574 20100 66580 20102
rect 66636 20100 66660 20102
rect 66716 20100 66740 20102
rect 66796 20100 66820 20102
rect 66876 20100 66882 20102
rect 66574 20091 66882 20100
rect 67234 19612 67542 19621
rect 67234 19610 67240 19612
rect 67296 19610 67320 19612
rect 67376 19610 67400 19612
rect 67456 19610 67480 19612
rect 67536 19610 67542 19612
rect 67296 19558 67298 19610
rect 67478 19558 67480 19610
rect 67234 19556 67240 19558
rect 67296 19556 67320 19558
rect 67376 19556 67400 19558
rect 67456 19556 67480 19558
rect 67536 19556 67542 19558
rect 67234 19547 67542 19556
rect 66574 19068 66882 19077
rect 66574 19066 66580 19068
rect 66636 19066 66660 19068
rect 66716 19066 66740 19068
rect 66796 19066 66820 19068
rect 66876 19066 66882 19068
rect 66636 19014 66638 19066
rect 66818 19014 66820 19066
rect 66574 19012 66580 19014
rect 66636 19012 66660 19014
rect 66716 19012 66740 19014
rect 66796 19012 66820 19014
rect 66876 19012 66882 19014
rect 66574 19003 66882 19012
rect 67234 18524 67542 18533
rect 67234 18522 67240 18524
rect 67296 18522 67320 18524
rect 67376 18522 67400 18524
rect 67456 18522 67480 18524
rect 67536 18522 67542 18524
rect 67296 18470 67298 18522
rect 67478 18470 67480 18522
rect 67234 18468 67240 18470
rect 67296 18468 67320 18470
rect 67376 18468 67400 18470
rect 67456 18468 67480 18470
rect 67536 18468 67542 18470
rect 67234 18459 67542 18468
rect 66574 17980 66882 17989
rect 66574 17978 66580 17980
rect 66636 17978 66660 17980
rect 66716 17978 66740 17980
rect 66796 17978 66820 17980
rect 66876 17978 66882 17980
rect 66636 17926 66638 17978
rect 66818 17926 66820 17978
rect 66574 17924 66580 17926
rect 66636 17924 66660 17926
rect 66716 17924 66740 17926
rect 66796 17924 66820 17926
rect 66876 17924 66882 17926
rect 66574 17915 66882 17924
rect 67234 17436 67542 17445
rect 67234 17434 67240 17436
rect 67296 17434 67320 17436
rect 67376 17434 67400 17436
rect 67456 17434 67480 17436
rect 67536 17434 67542 17436
rect 67296 17382 67298 17434
rect 67478 17382 67480 17434
rect 67234 17380 67240 17382
rect 67296 17380 67320 17382
rect 67376 17380 67400 17382
rect 67456 17380 67480 17382
rect 67536 17380 67542 17382
rect 67234 17371 67542 17380
rect 66574 16892 66882 16901
rect 66574 16890 66580 16892
rect 66636 16890 66660 16892
rect 66716 16890 66740 16892
rect 66796 16890 66820 16892
rect 66876 16890 66882 16892
rect 66636 16838 66638 16890
rect 66818 16838 66820 16890
rect 66574 16836 66580 16838
rect 66636 16836 66660 16838
rect 66716 16836 66740 16838
rect 66796 16836 66820 16838
rect 66876 16836 66882 16838
rect 66574 16827 66882 16836
rect 67234 16348 67542 16357
rect 67234 16346 67240 16348
rect 67296 16346 67320 16348
rect 67376 16346 67400 16348
rect 67456 16346 67480 16348
rect 67536 16346 67542 16348
rect 67296 16294 67298 16346
rect 67478 16294 67480 16346
rect 67234 16292 67240 16294
rect 67296 16292 67320 16294
rect 67376 16292 67400 16294
rect 67456 16292 67480 16294
rect 67536 16292 67542 16294
rect 67234 16283 67542 16292
rect 66574 15804 66882 15813
rect 66574 15802 66580 15804
rect 66636 15802 66660 15804
rect 66716 15802 66740 15804
rect 66796 15802 66820 15804
rect 66876 15802 66882 15804
rect 66636 15750 66638 15802
rect 66818 15750 66820 15802
rect 66574 15748 66580 15750
rect 66636 15748 66660 15750
rect 66716 15748 66740 15750
rect 66796 15748 66820 15750
rect 66876 15748 66882 15750
rect 66574 15739 66882 15748
rect 67234 15260 67542 15269
rect 67234 15258 67240 15260
rect 67296 15258 67320 15260
rect 67376 15258 67400 15260
rect 67456 15258 67480 15260
rect 67536 15258 67542 15260
rect 67296 15206 67298 15258
rect 67478 15206 67480 15258
rect 67234 15204 67240 15206
rect 67296 15204 67320 15206
rect 67376 15204 67400 15206
rect 67456 15204 67480 15206
rect 67536 15204 67542 15206
rect 67234 15195 67542 15204
rect 66574 14716 66882 14725
rect 66574 14714 66580 14716
rect 66636 14714 66660 14716
rect 66716 14714 66740 14716
rect 66796 14714 66820 14716
rect 66876 14714 66882 14716
rect 66636 14662 66638 14714
rect 66818 14662 66820 14714
rect 66574 14660 66580 14662
rect 66636 14660 66660 14662
rect 66716 14660 66740 14662
rect 66796 14660 66820 14662
rect 66876 14660 66882 14662
rect 66574 14651 66882 14660
rect 39118 14447 39174 14456
rect 58808 14476 58860 14482
rect 58808 14418 58860 14424
rect 36514 14172 36822 14181
rect 36514 14170 36520 14172
rect 36576 14170 36600 14172
rect 36656 14170 36680 14172
rect 36736 14170 36760 14172
rect 36816 14170 36822 14172
rect 36576 14118 36578 14170
rect 36758 14118 36760 14170
rect 36514 14116 36520 14118
rect 36576 14116 36600 14118
rect 36656 14116 36680 14118
rect 36736 14116 36760 14118
rect 36816 14116 36822 14118
rect 36514 14107 36822 14116
rect 67234 14172 67542 14181
rect 67234 14170 67240 14172
rect 67296 14170 67320 14172
rect 67376 14170 67400 14172
rect 67456 14170 67480 14172
rect 67536 14170 67542 14172
rect 67296 14118 67298 14170
rect 67478 14118 67480 14170
rect 67234 14116 67240 14118
rect 67296 14116 67320 14118
rect 67376 14116 67400 14118
rect 67456 14116 67480 14118
rect 67536 14116 67542 14118
rect 67234 14107 67542 14116
rect 35854 13628 36162 13637
rect 35854 13626 35860 13628
rect 35916 13626 35940 13628
rect 35996 13626 36020 13628
rect 36076 13626 36100 13628
rect 36156 13626 36162 13628
rect 35916 13574 35918 13626
rect 36098 13574 36100 13626
rect 35854 13572 35860 13574
rect 35916 13572 35940 13574
rect 35996 13572 36020 13574
rect 36076 13572 36100 13574
rect 36156 13572 36162 13574
rect 35854 13563 36162 13572
rect 66574 13628 66882 13637
rect 66574 13626 66580 13628
rect 66636 13626 66660 13628
rect 66716 13626 66740 13628
rect 66796 13626 66820 13628
rect 66876 13626 66882 13628
rect 66636 13574 66638 13626
rect 66818 13574 66820 13626
rect 66574 13572 66580 13574
rect 66636 13572 66660 13574
rect 66716 13572 66740 13574
rect 66796 13572 66820 13574
rect 66876 13572 66882 13574
rect 66574 13563 66882 13572
rect 36514 13084 36822 13093
rect 36514 13082 36520 13084
rect 36576 13082 36600 13084
rect 36656 13082 36680 13084
rect 36736 13082 36760 13084
rect 36816 13082 36822 13084
rect 36576 13030 36578 13082
rect 36758 13030 36760 13082
rect 36514 13028 36520 13030
rect 36576 13028 36600 13030
rect 36656 13028 36680 13030
rect 36736 13028 36760 13030
rect 36816 13028 36822 13030
rect 36514 13019 36822 13028
rect 67234 13084 67542 13093
rect 67234 13082 67240 13084
rect 67296 13082 67320 13084
rect 67376 13082 67400 13084
rect 67456 13082 67480 13084
rect 67536 13082 67542 13084
rect 67296 13030 67298 13082
rect 67478 13030 67480 13082
rect 67234 13028 67240 13030
rect 67296 13028 67320 13030
rect 67376 13028 67400 13030
rect 67456 13028 67480 13030
rect 67536 13028 67542 13030
rect 67234 13019 67542 13028
rect 38016 12640 38068 12646
rect 38016 12582 38068 12588
rect 35854 12540 36162 12549
rect 35854 12538 35860 12540
rect 35916 12538 35940 12540
rect 35996 12538 36020 12540
rect 36076 12538 36100 12540
rect 36156 12538 36162 12540
rect 35916 12486 35918 12538
rect 36098 12486 36100 12538
rect 35854 12484 35860 12486
rect 35916 12484 35940 12486
rect 35996 12484 36020 12486
rect 36076 12484 36100 12486
rect 36156 12484 36162 12486
rect 35854 12475 36162 12484
rect 36514 11996 36822 12005
rect 36514 11994 36520 11996
rect 36576 11994 36600 11996
rect 36656 11994 36680 11996
rect 36736 11994 36760 11996
rect 36816 11994 36822 11996
rect 36576 11942 36578 11994
rect 36758 11942 36760 11994
rect 36514 11940 36520 11942
rect 36576 11940 36600 11942
rect 36656 11940 36680 11942
rect 36736 11940 36760 11942
rect 36816 11940 36822 11942
rect 36514 11931 36822 11940
rect 36360 11892 36412 11898
rect 36360 11834 36412 11840
rect 35854 11452 36162 11461
rect 35854 11450 35860 11452
rect 35916 11450 35940 11452
rect 35996 11450 36020 11452
rect 36076 11450 36100 11452
rect 36156 11450 36162 11452
rect 35916 11398 35918 11450
rect 36098 11398 36100 11450
rect 35854 11396 35860 11398
rect 35916 11396 35940 11398
rect 35996 11396 36020 11398
rect 36076 11396 36100 11398
rect 36156 11396 36162 11398
rect 35854 11387 36162 11396
rect 32128 11076 32180 11082
rect 32128 11018 32180 11024
rect 31668 10532 31720 10538
rect 31668 10474 31720 10480
rect 31576 9648 31628 9654
rect 30932 9512 30984 9518
rect 30932 9454 30984 9460
rect 30840 8016 30892 8022
rect 30840 7958 30892 7964
rect 30840 7744 30892 7750
rect 30840 7686 30892 7692
rect 30852 6304 30880 7686
rect 30944 6497 30972 9454
rect 31036 7002 31064 9646
rect 31576 9590 31628 9596
rect 31300 9512 31352 9518
rect 31300 9454 31352 9460
rect 31576 9512 31628 9518
rect 31680 9500 31708 10474
rect 31850 10160 31906 10169
rect 31850 10095 31906 10104
rect 31864 10062 31892 10095
rect 31852 10056 31904 10062
rect 31852 9998 31904 10004
rect 31850 9616 31906 9625
rect 31850 9551 31906 9560
rect 31864 9500 31892 9551
rect 31680 9472 31892 9500
rect 31576 9454 31628 9460
rect 31116 8900 31168 8906
rect 31116 8842 31168 8848
rect 31128 8362 31156 8842
rect 31116 8356 31168 8362
rect 31116 8298 31168 8304
rect 31208 8288 31260 8294
rect 31208 8230 31260 8236
rect 31220 7970 31248 8230
rect 31128 7942 31248 7970
rect 31128 7410 31156 7942
rect 31208 7880 31260 7886
rect 31208 7822 31260 7828
rect 31116 7404 31168 7410
rect 31116 7346 31168 7352
rect 31024 6996 31076 7002
rect 31024 6938 31076 6944
rect 31114 6896 31170 6905
rect 31114 6831 31170 6840
rect 31128 6798 31156 6831
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 31220 6662 31248 7822
rect 31208 6656 31260 6662
rect 31208 6598 31260 6604
rect 30930 6488 30986 6497
rect 30930 6423 30986 6432
rect 30852 6276 31064 6304
rect 30930 6216 30986 6225
rect 30930 6151 30986 6160
rect 30840 6112 30892 6118
rect 30840 6054 30892 6060
rect 30852 5778 30880 6054
rect 30840 5772 30892 5778
rect 30840 5714 30892 5720
rect 30838 4856 30894 4865
rect 30838 4791 30894 4800
rect 30852 4690 30880 4791
rect 30840 4684 30892 4690
rect 30840 4626 30892 4632
rect 30838 4312 30894 4321
rect 30838 4247 30894 4256
rect 30748 3528 30800 3534
rect 30748 3470 30800 3476
rect 30656 3392 30708 3398
rect 30656 3334 30708 3340
rect 30852 2854 30880 4247
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 30840 2848 30892 2854
rect 30840 2790 30892 2796
rect 30472 1964 30524 1970
rect 30472 1906 30524 1912
rect 30944 800 30972 6151
rect 31036 3108 31064 6276
rect 31206 6216 31262 6225
rect 31206 6151 31262 6160
rect 31220 5778 31248 6151
rect 31208 5772 31260 5778
rect 31208 5714 31260 5720
rect 31206 5400 31262 5409
rect 31206 5335 31262 5344
rect 31220 4622 31248 5335
rect 31312 4826 31340 9454
rect 31392 9376 31444 9382
rect 31392 9318 31444 9324
rect 31404 8401 31432 9318
rect 31390 8392 31446 8401
rect 31390 8327 31446 8336
rect 31390 8120 31446 8129
rect 31390 8055 31446 8064
rect 31404 7886 31432 8055
rect 31482 7984 31538 7993
rect 31482 7919 31538 7928
rect 31392 7880 31444 7886
rect 31392 7822 31444 7828
rect 31392 7744 31444 7750
rect 31392 7686 31444 7692
rect 31404 7478 31432 7686
rect 31392 7472 31444 7478
rect 31392 7414 31444 7420
rect 31404 6934 31432 7414
rect 31392 6928 31444 6934
rect 31392 6870 31444 6876
rect 31496 6390 31524 7919
rect 31484 6384 31536 6390
rect 31484 6326 31536 6332
rect 31496 5710 31524 6326
rect 31484 5704 31536 5710
rect 31484 5646 31536 5652
rect 31588 5273 31616 9454
rect 31864 8974 31892 9472
rect 32036 9512 32088 9518
rect 32036 9454 32088 9460
rect 31944 9104 31996 9110
rect 31944 9046 31996 9052
rect 31852 8968 31904 8974
rect 31852 8910 31904 8916
rect 31668 8900 31720 8906
rect 31668 8842 31720 8848
rect 31680 8294 31708 8842
rect 31760 8832 31812 8838
rect 31760 8774 31812 8780
rect 31772 8401 31800 8774
rect 31758 8392 31814 8401
rect 31758 8327 31814 8336
rect 31668 8288 31720 8294
rect 31668 8230 31720 8236
rect 31680 7993 31708 8230
rect 31666 7984 31722 7993
rect 31666 7919 31722 7928
rect 31760 7880 31812 7886
rect 31758 7848 31760 7857
rect 31812 7848 31814 7857
rect 31758 7783 31814 7792
rect 31666 7712 31722 7721
rect 31666 7647 31722 7656
rect 31680 7546 31708 7647
rect 31668 7540 31720 7546
rect 31668 7482 31720 7488
rect 31668 7404 31720 7410
rect 31668 7346 31720 7352
rect 31680 6866 31708 7346
rect 31772 6934 31800 7783
rect 31864 7041 31892 8910
rect 31956 8838 31984 9046
rect 31944 8832 31996 8838
rect 31944 8774 31996 8780
rect 31944 8492 31996 8498
rect 31944 8434 31996 8440
rect 31956 7449 31984 8434
rect 31942 7440 31998 7449
rect 31942 7375 31998 7384
rect 31850 7032 31906 7041
rect 31850 6967 31906 6976
rect 31760 6928 31812 6934
rect 31760 6870 31812 6876
rect 31668 6860 31720 6866
rect 31668 6802 31720 6808
rect 31680 6225 31708 6802
rect 31956 6798 31984 7375
rect 31852 6792 31904 6798
rect 31852 6734 31904 6740
rect 31944 6792 31996 6798
rect 31944 6734 31996 6740
rect 31864 6390 31892 6734
rect 31944 6656 31996 6662
rect 31944 6598 31996 6604
rect 31852 6384 31904 6390
rect 31852 6326 31904 6332
rect 31956 6322 31984 6598
rect 31944 6316 31996 6322
rect 31944 6258 31996 6264
rect 31666 6216 31722 6225
rect 31666 6151 31722 6160
rect 31666 5808 31722 5817
rect 31666 5743 31722 5752
rect 31680 5710 31708 5743
rect 31668 5704 31720 5710
rect 31944 5704 31996 5710
rect 31668 5646 31720 5652
rect 31772 5664 31944 5692
rect 31574 5264 31630 5273
rect 31574 5199 31630 5208
rect 31300 4820 31352 4826
rect 31300 4762 31352 4768
rect 31576 4820 31628 4826
rect 31576 4762 31628 4768
rect 31208 4616 31260 4622
rect 31208 4558 31260 4564
rect 31588 4554 31616 4762
rect 31668 4752 31720 4758
rect 31668 4694 31720 4700
rect 31576 4548 31628 4554
rect 31576 4490 31628 4496
rect 31116 4276 31168 4282
rect 31116 4218 31168 4224
rect 31128 4146 31156 4218
rect 31116 4140 31168 4146
rect 31116 4082 31168 4088
rect 31680 4010 31708 4694
rect 31576 4004 31628 4010
rect 31576 3946 31628 3952
rect 31668 4004 31720 4010
rect 31668 3946 31720 3952
rect 31300 3596 31352 3602
rect 31300 3538 31352 3544
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 31220 3126 31248 3470
rect 31116 3120 31168 3126
rect 31036 3080 31116 3108
rect 31116 3062 31168 3068
rect 31208 3120 31260 3126
rect 31208 3062 31260 3068
rect 31312 2990 31340 3538
rect 31300 2984 31352 2990
rect 31300 2926 31352 2932
rect 31392 2304 31444 2310
rect 31392 2246 31444 2252
rect 31404 1766 31432 2246
rect 31588 2038 31616 3946
rect 31772 3233 31800 5664
rect 31944 5646 31996 5652
rect 31850 5536 31906 5545
rect 31850 5471 31906 5480
rect 31864 5370 31892 5471
rect 31852 5364 31904 5370
rect 31852 5306 31904 5312
rect 31852 5024 31904 5030
rect 31852 4966 31904 4972
rect 31864 4690 31892 4966
rect 31852 4684 31904 4690
rect 31852 4626 31904 4632
rect 32048 3670 32076 9454
rect 32140 6390 32168 11018
rect 34244 10736 34296 10742
rect 34244 10678 34296 10684
rect 33876 10668 33928 10674
rect 33876 10610 33928 10616
rect 33140 10600 33192 10606
rect 33140 10542 33192 10548
rect 33324 10600 33376 10606
rect 33324 10542 33376 10548
rect 33600 10600 33652 10606
rect 33600 10542 33652 10548
rect 32312 10464 32364 10470
rect 32312 10406 32364 10412
rect 32496 10464 32548 10470
rect 32496 10406 32548 10412
rect 32220 9512 32272 9518
rect 32220 9454 32272 9460
rect 32232 8673 32260 9454
rect 32218 8664 32274 8673
rect 32218 8599 32274 8608
rect 32220 8424 32272 8430
rect 32220 8366 32272 8372
rect 32232 7546 32260 8366
rect 32324 7857 32352 10406
rect 32404 9988 32456 9994
rect 32404 9930 32456 9936
rect 32416 8974 32444 9930
rect 32404 8968 32456 8974
rect 32404 8910 32456 8916
rect 32404 8832 32456 8838
rect 32404 8774 32456 8780
rect 32416 8634 32444 8774
rect 32404 8628 32456 8634
rect 32404 8570 32456 8576
rect 32404 8424 32456 8430
rect 32404 8366 32456 8372
rect 32416 8265 32444 8366
rect 32402 8256 32458 8265
rect 32402 8191 32458 8200
rect 32310 7848 32366 7857
rect 32310 7783 32366 7792
rect 32404 7812 32456 7818
rect 32404 7754 32456 7760
rect 32312 7744 32364 7750
rect 32310 7712 32312 7721
rect 32364 7712 32366 7721
rect 32310 7647 32366 7656
rect 32220 7540 32272 7546
rect 32220 7482 32272 7488
rect 32312 7404 32364 7410
rect 32312 7346 32364 7352
rect 32218 7304 32274 7313
rect 32218 7239 32220 7248
rect 32272 7239 32274 7248
rect 32220 7210 32272 7216
rect 32128 6384 32180 6390
rect 32128 6326 32180 6332
rect 32232 6322 32260 7210
rect 32324 7041 32352 7346
rect 32416 7206 32444 7754
rect 32508 7410 32536 10406
rect 32956 10124 33008 10130
rect 32956 10066 33008 10072
rect 32588 10056 32640 10062
rect 32588 9998 32640 10004
rect 32864 10056 32916 10062
rect 32864 9998 32916 10004
rect 32496 7404 32548 7410
rect 32496 7346 32548 7352
rect 32404 7200 32456 7206
rect 32404 7142 32456 7148
rect 32310 7032 32366 7041
rect 32310 6967 32366 6976
rect 32220 6316 32272 6322
rect 32220 6258 32272 6264
rect 32220 6180 32272 6186
rect 32220 6122 32272 6128
rect 32126 6080 32182 6089
rect 32126 6015 32182 6024
rect 32140 5681 32168 6015
rect 32232 5953 32260 6122
rect 32218 5944 32274 5953
rect 32218 5879 32274 5888
rect 32126 5672 32182 5681
rect 32232 5642 32260 5879
rect 32126 5607 32182 5616
rect 32220 5636 32272 5642
rect 32220 5578 32272 5584
rect 32218 5264 32274 5273
rect 32324 5234 32352 6967
rect 32416 6497 32444 7142
rect 32402 6488 32458 6497
rect 32402 6423 32458 6432
rect 32416 5370 32444 6423
rect 32404 5364 32456 5370
rect 32456 5324 32536 5352
rect 32404 5306 32456 5312
rect 32218 5199 32274 5208
rect 32312 5228 32364 5234
rect 32126 4856 32182 4865
rect 32126 4791 32182 4800
rect 32140 4486 32168 4791
rect 32232 4690 32260 5199
rect 32312 5170 32364 5176
rect 32402 4992 32458 5001
rect 32402 4927 32458 4936
rect 32220 4684 32272 4690
rect 32220 4626 32272 4632
rect 32128 4480 32180 4486
rect 32128 4422 32180 4428
rect 32232 4282 32260 4626
rect 32220 4276 32272 4282
rect 32220 4218 32272 4224
rect 31852 3664 31904 3670
rect 31852 3606 31904 3612
rect 32036 3664 32088 3670
rect 32036 3606 32088 3612
rect 31864 3466 31892 3606
rect 31852 3460 31904 3466
rect 31852 3402 31904 3408
rect 31758 3224 31814 3233
rect 31758 3159 31814 3168
rect 32232 2990 32260 4218
rect 32416 3466 32444 4927
rect 32508 4282 32536 5324
rect 32496 4276 32548 4282
rect 32496 4218 32548 4224
rect 32496 4072 32548 4078
rect 32600 4060 32628 9998
rect 32680 9920 32732 9926
rect 32680 9862 32732 9868
rect 32692 4146 32720 9862
rect 32876 9654 32904 9998
rect 32864 9648 32916 9654
rect 32864 9590 32916 9596
rect 32772 9376 32824 9382
rect 32772 9318 32824 9324
rect 32784 4826 32812 9318
rect 32864 9172 32916 9178
rect 32864 9114 32916 9120
rect 32876 7546 32904 9114
rect 32864 7540 32916 7546
rect 32864 7482 32916 7488
rect 32864 7336 32916 7342
rect 32864 7278 32916 7284
rect 32876 7002 32904 7278
rect 32864 6996 32916 7002
rect 32864 6938 32916 6944
rect 32968 5250 32996 10066
rect 33046 9616 33102 9625
rect 33046 9551 33048 9560
rect 33100 9551 33102 9560
rect 33048 9522 33100 9528
rect 33152 9178 33180 10542
rect 33336 9722 33364 10542
rect 33416 9920 33468 9926
rect 33416 9862 33468 9868
rect 33324 9716 33376 9722
rect 33324 9658 33376 9664
rect 33232 9580 33284 9586
rect 33232 9522 33284 9528
rect 33244 9489 33272 9522
rect 33230 9480 33286 9489
rect 33230 9415 33286 9424
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 33140 8968 33192 8974
rect 33336 8922 33364 9658
rect 33140 8910 33192 8916
rect 33046 8800 33102 8809
rect 33046 8735 33102 8744
rect 33060 8498 33088 8735
rect 33152 8673 33180 8910
rect 33244 8894 33364 8922
rect 33138 8664 33194 8673
rect 33138 8599 33194 8608
rect 33140 8560 33192 8566
rect 33140 8502 33192 8508
rect 33048 8492 33100 8498
rect 33048 8434 33100 8440
rect 33152 8129 33180 8502
rect 33138 8120 33194 8129
rect 33138 8055 33194 8064
rect 33048 7540 33100 7546
rect 33048 7482 33100 7488
rect 33060 6225 33088 7482
rect 33140 7472 33192 7478
rect 33140 7414 33192 7420
rect 33152 6798 33180 7414
rect 33244 7410 33272 8894
rect 33324 8832 33376 8838
rect 33324 8774 33376 8780
rect 33336 8401 33364 8774
rect 33322 8392 33378 8401
rect 33322 8327 33378 8336
rect 33324 8288 33376 8294
rect 33324 8230 33376 8236
rect 33232 7404 33284 7410
rect 33232 7346 33284 7352
rect 33232 6860 33284 6866
rect 33232 6802 33284 6808
rect 33140 6792 33192 6798
rect 33140 6734 33192 6740
rect 33046 6216 33102 6225
rect 33046 6151 33102 6160
rect 32876 5222 32996 5250
rect 33060 5250 33088 6151
rect 33152 5370 33180 6734
rect 33244 6390 33272 6802
rect 33336 6633 33364 8230
rect 33322 6624 33378 6633
rect 33322 6559 33378 6568
rect 33232 6384 33284 6390
rect 33232 6326 33284 6332
rect 33140 5364 33192 5370
rect 33140 5306 33192 5312
rect 33060 5222 33180 5250
rect 32772 4820 32824 4826
rect 32772 4762 32824 4768
rect 32680 4140 32732 4146
rect 32680 4082 32732 4088
rect 32548 4032 32628 4060
rect 32784 4026 32812 4762
rect 32496 4014 32548 4020
rect 32692 3998 32812 4026
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 32692 3194 32720 3998
rect 32772 3936 32824 3942
rect 32772 3878 32824 3884
rect 32784 3602 32812 3878
rect 32772 3596 32824 3602
rect 32772 3538 32824 3544
rect 32876 3505 32904 5222
rect 32956 5160 33008 5166
rect 32956 5102 33008 5108
rect 32968 4690 32996 5102
rect 32956 4684 33008 4690
rect 32956 4626 33008 4632
rect 32956 4276 33008 4282
rect 32956 4218 33008 4224
rect 32862 3496 32918 3505
rect 32968 3466 32996 4218
rect 33048 4140 33100 4146
rect 33048 4082 33100 4088
rect 33060 3913 33088 4082
rect 33046 3904 33102 3913
rect 33046 3839 33102 3848
rect 32862 3431 32918 3440
rect 32956 3460 33008 3466
rect 32956 3402 33008 3408
rect 32680 3188 32732 3194
rect 32680 3130 32732 3136
rect 32968 3126 32996 3402
rect 33152 3126 33180 5222
rect 33232 5024 33284 5030
rect 33232 4966 33284 4972
rect 33244 4146 33272 4966
rect 33322 4584 33378 4593
rect 33322 4519 33378 4528
rect 33232 4140 33284 4146
rect 33232 4082 33284 4088
rect 33336 3738 33364 4519
rect 33324 3732 33376 3738
rect 33324 3674 33376 3680
rect 33336 3194 33364 3674
rect 33324 3188 33376 3194
rect 33324 3130 33376 3136
rect 32956 3120 33008 3126
rect 32956 3062 33008 3068
rect 33140 3120 33192 3126
rect 33140 3062 33192 3068
rect 32220 2984 32272 2990
rect 32220 2926 32272 2932
rect 33046 2952 33102 2961
rect 33046 2887 33048 2896
rect 33100 2887 33102 2896
rect 33048 2858 33100 2864
rect 32220 2508 32272 2514
rect 32220 2450 32272 2456
rect 31576 2032 31628 2038
rect 31576 1974 31628 1980
rect 31392 1760 31444 1766
rect 31392 1702 31444 1708
rect 31496 870 31616 898
rect 25240 734 25452 762
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31496 338 31524 870
rect 31588 800 31616 870
rect 32232 800 32260 2450
rect 32772 2440 32824 2446
rect 32772 2382 32824 2388
rect 33324 2440 33376 2446
rect 33428 2428 33456 9862
rect 33508 9580 33560 9586
rect 33508 9522 33560 9528
rect 33520 9178 33548 9522
rect 33508 9172 33560 9178
rect 33508 9114 33560 9120
rect 33508 8900 33560 8906
rect 33508 8842 33560 8848
rect 33520 8498 33548 8842
rect 33508 8492 33560 8498
rect 33508 8434 33560 8440
rect 33508 7948 33560 7954
rect 33508 7890 33560 7896
rect 33520 7410 33548 7890
rect 33508 7404 33560 7410
rect 33508 7346 33560 7352
rect 33508 6792 33560 6798
rect 33508 6734 33560 6740
rect 33520 6662 33548 6734
rect 33508 6656 33560 6662
rect 33508 6598 33560 6604
rect 33508 5840 33560 5846
rect 33508 5782 33560 5788
rect 33520 5302 33548 5782
rect 33508 5296 33560 5302
rect 33508 5238 33560 5244
rect 33506 4448 33562 4457
rect 33506 4383 33562 4392
rect 33520 3194 33548 4383
rect 33508 3188 33560 3194
rect 33508 3130 33560 3136
rect 33612 2774 33640 10542
rect 33690 9344 33746 9353
rect 33690 9279 33746 9288
rect 33704 5710 33732 9279
rect 33888 8838 33916 10610
rect 34152 9376 34204 9382
rect 34152 9318 34204 9324
rect 34060 9036 34112 9042
rect 33980 8996 34060 9024
rect 33876 8832 33928 8838
rect 33876 8774 33928 8780
rect 33888 8498 33916 8774
rect 33784 8492 33836 8498
rect 33784 8434 33836 8440
rect 33876 8492 33928 8498
rect 33876 8434 33928 8440
rect 33796 7585 33824 8434
rect 33888 8362 33916 8434
rect 33876 8356 33928 8362
rect 33876 8298 33928 8304
rect 33874 8120 33930 8129
rect 33874 8055 33930 8064
rect 33888 7954 33916 8055
rect 33876 7948 33928 7954
rect 33876 7890 33928 7896
rect 33782 7576 33838 7585
rect 33782 7511 33838 7520
rect 33782 6488 33838 6497
rect 33782 6423 33838 6432
rect 33796 6390 33824 6423
rect 33784 6384 33836 6390
rect 33784 6326 33836 6332
rect 33876 6112 33928 6118
rect 33876 6054 33928 6060
rect 33784 5908 33836 5914
rect 33784 5850 33836 5856
rect 33692 5704 33744 5710
rect 33692 5646 33744 5652
rect 33692 5568 33744 5574
rect 33692 5510 33744 5516
rect 33704 5370 33732 5510
rect 33692 5364 33744 5370
rect 33692 5306 33744 5312
rect 33796 4826 33824 5850
rect 33888 5166 33916 6054
rect 33980 5681 34008 8996
rect 34060 8978 34112 8984
rect 34164 8566 34192 9318
rect 34152 8560 34204 8566
rect 34152 8502 34204 8508
rect 34152 8356 34204 8362
rect 34152 8298 34204 8304
rect 34164 7954 34192 8298
rect 34152 7948 34204 7954
rect 34152 7890 34204 7896
rect 34060 7404 34112 7410
rect 34060 7346 34112 7352
rect 34072 6662 34100 7346
rect 34060 6656 34112 6662
rect 34060 6598 34112 6604
rect 34164 6458 34192 7890
rect 34256 7732 34284 10678
rect 34888 10668 34940 10674
rect 34888 10610 34940 10616
rect 35164 10668 35216 10674
rect 35164 10610 35216 10616
rect 34796 10464 34848 10470
rect 34796 10406 34848 10412
rect 34336 10260 34388 10266
rect 34336 10202 34388 10208
rect 34348 7886 34376 10202
rect 34808 10130 34836 10406
rect 34796 10124 34848 10130
rect 34796 10066 34848 10072
rect 34520 8968 34572 8974
rect 34520 8910 34572 8916
rect 34532 8838 34560 8910
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34428 8492 34480 8498
rect 34428 8434 34480 8440
rect 34336 7880 34388 7886
rect 34336 7822 34388 7828
rect 34440 7818 34468 8434
rect 34428 7812 34480 7818
rect 34428 7754 34480 7760
rect 34336 7744 34388 7750
rect 34256 7704 34336 7732
rect 34336 7686 34388 7692
rect 34440 7562 34468 7754
rect 34256 7534 34468 7562
rect 34256 7206 34284 7534
rect 34336 7336 34388 7342
rect 34336 7278 34388 7284
rect 34428 7336 34480 7342
rect 34428 7278 34480 7284
rect 34244 7200 34296 7206
rect 34244 7142 34296 7148
rect 34256 6730 34284 7142
rect 34244 6724 34296 6730
rect 34244 6666 34296 6672
rect 34348 6633 34376 7278
rect 34440 6866 34468 7278
rect 34428 6860 34480 6866
rect 34428 6802 34480 6808
rect 34428 6724 34480 6730
rect 34428 6666 34480 6672
rect 34334 6624 34390 6633
rect 34334 6559 34390 6568
rect 34152 6452 34204 6458
rect 34152 6394 34204 6400
rect 34244 6452 34296 6458
rect 34244 6394 34296 6400
rect 34164 5846 34192 6394
rect 34152 5840 34204 5846
rect 34152 5782 34204 5788
rect 33966 5672 34022 5681
rect 33966 5607 34022 5616
rect 34150 5672 34206 5681
rect 34150 5607 34206 5616
rect 33968 5568 34020 5574
rect 33968 5510 34020 5516
rect 33876 5160 33928 5166
rect 33876 5102 33928 5108
rect 33784 4820 33836 4826
rect 33784 4762 33836 4768
rect 33784 4480 33836 4486
rect 33784 4422 33836 4428
rect 33796 3505 33824 4422
rect 33980 4078 34008 5510
rect 34060 5228 34112 5234
rect 34060 5170 34112 5176
rect 34072 4282 34100 5170
rect 34060 4276 34112 4282
rect 34060 4218 34112 4224
rect 33968 4072 34020 4078
rect 33968 4014 34020 4020
rect 34058 3632 34114 3641
rect 34058 3567 34114 3576
rect 33782 3496 33838 3505
rect 33782 3431 33838 3440
rect 33782 3360 33838 3369
rect 33782 3295 33838 3304
rect 33796 3058 33824 3295
rect 33874 3224 33930 3233
rect 34072 3194 34100 3567
rect 33874 3159 33930 3168
rect 34060 3188 34112 3194
rect 33888 3058 33916 3159
rect 34060 3130 34112 3136
rect 33784 3052 33836 3058
rect 33784 2994 33836 3000
rect 33876 3052 33928 3058
rect 33876 2994 33928 3000
rect 33376 2400 33456 2428
rect 33520 2746 33640 2774
rect 33324 2382 33376 2388
rect 32784 1834 32812 2382
rect 32772 1828 32824 1834
rect 32772 1770 32824 1776
rect 32784 870 32904 898
rect 31484 332 31536 338
rect 31484 274 31536 280
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32784 270 32812 870
rect 32876 800 32904 870
rect 33520 800 33548 2746
rect 34164 2582 34192 5607
rect 34256 5409 34284 6394
rect 34348 5778 34376 6559
rect 34336 5772 34388 5778
rect 34336 5714 34388 5720
rect 34336 5636 34388 5642
rect 34336 5578 34388 5584
rect 34242 5400 34298 5409
rect 34242 5335 34298 5344
rect 34244 5092 34296 5098
rect 34244 5034 34296 5040
rect 34256 3738 34284 5034
rect 34244 3732 34296 3738
rect 34244 3674 34296 3680
rect 34348 3641 34376 5578
rect 34334 3632 34390 3641
rect 34334 3567 34390 3576
rect 34440 3534 34468 6666
rect 34532 4078 34560 8774
rect 34796 8560 34848 8566
rect 34796 8502 34848 8508
rect 34612 8424 34664 8430
rect 34612 8366 34664 8372
rect 34624 7546 34652 8366
rect 34702 8256 34758 8265
rect 34702 8191 34758 8200
rect 34612 7540 34664 7546
rect 34612 7482 34664 7488
rect 34612 6928 34664 6934
rect 34612 6870 34664 6876
rect 34624 6730 34652 6870
rect 34716 6866 34744 8191
rect 34808 7970 34836 8502
rect 34900 8090 34928 10610
rect 34980 9512 35032 9518
rect 34980 9454 35032 9460
rect 34888 8084 34940 8090
rect 34888 8026 34940 8032
rect 34808 7942 34928 7970
rect 34900 7886 34928 7942
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 34888 7880 34940 7886
rect 34888 7822 34940 7828
rect 34704 6860 34756 6866
rect 34704 6802 34756 6808
rect 34612 6724 34664 6730
rect 34612 6666 34664 6672
rect 34624 6390 34652 6666
rect 34612 6384 34664 6390
rect 34612 6326 34664 6332
rect 34704 5568 34756 5574
rect 34704 5510 34756 5516
rect 34610 5264 34666 5273
rect 34610 5199 34612 5208
rect 34664 5199 34666 5208
rect 34612 5170 34664 5176
rect 34612 4616 34664 4622
rect 34612 4558 34664 4564
rect 34624 4214 34652 4558
rect 34612 4208 34664 4214
rect 34612 4150 34664 4156
rect 34520 4072 34572 4078
rect 34520 4014 34572 4020
rect 34428 3528 34480 3534
rect 34716 3482 34744 5510
rect 34808 3738 34836 7822
rect 34886 6896 34942 6905
rect 34886 6831 34942 6840
rect 34900 6798 34928 6831
rect 34888 6792 34940 6798
rect 34888 6734 34940 6740
rect 34992 5658 35020 9454
rect 35072 9444 35124 9450
rect 35072 9386 35124 9392
rect 35084 8974 35112 9386
rect 35072 8968 35124 8974
rect 35072 8910 35124 8916
rect 35072 8832 35124 8838
rect 35072 8774 35124 8780
rect 35084 8566 35112 8774
rect 35072 8560 35124 8566
rect 35072 8502 35124 8508
rect 35072 8424 35124 8430
rect 35072 8366 35124 8372
rect 35084 5794 35112 8366
rect 35176 7002 35204 10610
rect 35440 10464 35492 10470
rect 35440 10406 35492 10412
rect 35348 9444 35400 9450
rect 35348 9386 35400 9392
rect 35256 9376 35308 9382
rect 35256 9318 35308 9324
rect 35268 8537 35296 9318
rect 35254 8528 35310 8537
rect 35254 8463 35310 8472
rect 35164 6996 35216 7002
rect 35164 6938 35216 6944
rect 35256 6928 35308 6934
rect 35256 6870 35308 6876
rect 35164 6792 35216 6798
rect 35162 6760 35164 6769
rect 35216 6760 35218 6769
rect 35162 6695 35218 6704
rect 35164 6656 35216 6662
rect 35164 6598 35216 6604
rect 35176 6225 35204 6598
rect 35162 6216 35218 6225
rect 35162 6151 35218 6160
rect 35268 5914 35296 6870
rect 35256 5908 35308 5914
rect 35256 5850 35308 5856
rect 35084 5766 35296 5794
rect 34992 5630 35112 5658
rect 34980 5568 35032 5574
rect 34980 5510 35032 5516
rect 34888 5092 34940 5098
rect 34888 5034 34940 5040
rect 34900 4690 34928 5034
rect 34992 4758 35020 5510
rect 34980 4752 35032 4758
rect 34980 4694 35032 4700
rect 34888 4684 34940 4690
rect 34888 4626 34940 4632
rect 34888 4072 34940 4078
rect 34888 4014 34940 4020
rect 34796 3732 34848 3738
rect 34796 3674 34848 3680
rect 34428 3470 34480 3476
rect 34532 3454 34744 3482
rect 34532 3176 34560 3454
rect 34612 3392 34664 3398
rect 34612 3334 34664 3340
rect 34624 3194 34652 3334
rect 34440 3148 34560 3176
rect 34612 3188 34664 3194
rect 34440 2922 34468 3148
rect 34612 3130 34664 3136
rect 34612 2984 34664 2990
rect 34612 2926 34664 2932
rect 34428 2916 34480 2922
rect 34428 2858 34480 2864
rect 34624 2650 34652 2926
rect 34900 2854 34928 4014
rect 35084 3466 35112 5630
rect 35164 5228 35216 5234
rect 35164 5170 35216 5176
rect 35176 5030 35204 5170
rect 35164 5024 35216 5030
rect 35164 4966 35216 4972
rect 35268 4321 35296 5766
rect 35254 4312 35310 4321
rect 35254 4247 35310 4256
rect 35164 4072 35216 4078
rect 35164 4014 35216 4020
rect 35176 3602 35204 4014
rect 35256 4004 35308 4010
rect 35256 3946 35308 3952
rect 35164 3596 35216 3602
rect 35164 3538 35216 3544
rect 34980 3460 35032 3466
rect 34980 3402 35032 3408
rect 35072 3460 35124 3466
rect 35072 3402 35124 3408
rect 34888 2848 34940 2854
rect 34888 2790 34940 2796
rect 34612 2644 34664 2650
rect 34612 2586 34664 2592
rect 34152 2576 34204 2582
rect 34152 2518 34204 2524
rect 34152 2372 34204 2378
rect 34152 2314 34204 2320
rect 34164 800 34192 2314
rect 34992 2310 35020 3402
rect 35176 3369 35204 3538
rect 35162 3360 35218 3369
rect 35162 3295 35218 3304
rect 35072 2848 35124 2854
rect 35072 2790 35124 2796
rect 34980 2304 35032 2310
rect 34980 2246 35032 2252
rect 34808 870 34928 898
rect 34808 800 34836 870
rect 32772 264 32824 270
rect 32772 206 32824 212
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 34900 762 34928 870
rect 35084 762 35112 2790
rect 35268 2446 35296 3946
rect 35360 2774 35388 9386
rect 35452 9042 35480 10406
rect 35854 10364 36162 10373
rect 35854 10362 35860 10364
rect 35916 10362 35940 10364
rect 35996 10362 36020 10364
rect 36076 10362 36100 10364
rect 36156 10362 36162 10364
rect 35916 10310 35918 10362
rect 36098 10310 36100 10362
rect 35854 10308 35860 10310
rect 35916 10308 35940 10310
rect 35996 10308 36020 10310
rect 36076 10308 36100 10310
rect 36156 10308 36162 10310
rect 35854 10299 36162 10308
rect 35624 10056 35676 10062
rect 35624 9998 35676 10004
rect 35636 9178 35664 9998
rect 36268 9920 36320 9926
rect 36268 9862 36320 9868
rect 36280 9586 36308 9862
rect 36372 9674 36400 11834
rect 36514 10908 36822 10917
rect 36514 10906 36520 10908
rect 36576 10906 36600 10908
rect 36656 10906 36680 10908
rect 36736 10906 36760 10908
rect 36816 10906 36822 10908
rect 36576 10854 36578 10906
rect 36758 10854 36760 10906
rect 36514 10852 36520 10854
rect 36576 10852 36600 10854
rect 36656 10852 36680 10854
rect 36736 10852 36760 10854
rect 36816 10852 36822 10854
rect 36514 10843 36822 10852
rect 37188 10192 37240 10198
rect 37188 10134 37240 10140
rect 36912 10056 36964 10062
rect 36912 9998 36964 10004
rect 36514 9820 36822 9829
rect 36514 9818 36520 9820
rect 36576 9818 36600 9820
rect 36656 9818 36680 9820
rect 36736 9818 36760 9820
rect 36816 9818 36822 9820
rect 36576 9766 36578 9818
rect 36758 9766 36760 9818
rect 36514 9764 36520 9766
rect 36576 9764 36600 9766
rect 36656 9764 36680 9766
rect 36736 9764 36760 9766
rect 36816 9764 36822 9766
rect 36514 9755 36822 9764
rect 36372 9646 36492 9674
rect 36268 9580 36320 9586
rect 36268 9522 36320 9528
rect 36360 9512 36412 9518
rect 35714 9480 35770 9489
rect 36360 9454 36412 9460
rect 35714 9415 35770 9424
rect 35624 9172 35676 9178
rect 35624 9114 35676 9120
rect 35440 9036 35492 9042
rect 35440 8978 35492 8984
rect 35728 8922 35756 9415
rect 35854 9276 36162 9285
rect 35854 9274 35860 9276
rect 35916 9274 35940 9276
rect 35996 9274 36020 9276
rect 36076 9274 36100 9276
rect 36156 9274 36162 9276
rect 35916 9222 35918 9274
rect 36098 9222 36100 9274
rect 35854 9220 35860 9222
rect 35916 9220 35940 9222
rect 35996 9220 36020 9222
rect 36076 9220 36100 9222
rect 36156 9220 36162 9222
rect 35854 9211 36162 9220
rect 36084 9104 36136 9110
rect 36084 9046 36136 9052
rect 35728 8894 35848 8922
rect 35716 8832 35768 8838
rect 35716 8774 35768 8780
rect 35728 8430 35756 8774
rect 35820 8430 35848 8894
rect 36096 8498 36124 9046
rect 36372 9024 36400 9454
rect 36464 9110 36492 9646
rect 36452 9104 36504 9110
rect 36452 9046 36504 9052
rect 36188 8996 36400 9024
rect 36188 8650 36216 8996
rect 36268 8900 36320 8906
rect 36320 8860 36400 8888
rect 36268 8842 36320 8848
rect 36188 8622 36308 8650
rect 36084 8492 36136 8498
rect 36084 8434 36136 8440
rect 35716 8424 35768 8430
rect 35716 8366 35768 8372
rect 35808 8424 35860 8430
rect 35808 8366 35860 8372
rect 35820 8276 35848 8366
rect 35728 8248 35848 8276
rect 35624 7744 35676 7750
rect 35624 7686 35676 7692
rect 35532 7268 35584 7274
rect 35532 7210 35584 7216
rect 35440 6928 35492 6934
rect 35440 6870 35492 6876
rect 35452 6322 35480 6870
rect 35440 6316 35492 6322
rect 35440 6258 35492 6264
rect 35440 6112 35492 6118
rect 35440 6054 35492 6060
rect 35452 5166 35480 6054
rect 35544 5710 35572 7210
rect 35532 5704 35584 5710
rect 35532 5646 35584 5652
rect 35440 5160 35492 5166
rect 35440 5102 35492 5108
rect 35440 4480 35492 4486
rect 35440 4422 35492 4428
rect 35452 3602 35480 4422
rect 35532 3936 35584 3942
rect 35532 3878 35584 3884
rect 35440 3596 35492 3602
rect 35440 3538 35492 3544
rect 35544 2854 35572 3878
rect 35636 3126 35664 7686
rect 35728 7410 35756 8248
rect 35854 8188 36162 8197
rect 35854 8186 35860 8188
rect 35916 8186 35940 8188
rect 35996 8186 36020 8188
rect 36076 8186 36100 8188
rect 36156 8186 36162 8188
rect 35916 8134 35918 8186
rect 36098 8134 36100 8186
rect 35854 8132 35860 8134
rect 35916 8132 35940 8134
rect 35996 8132 36020 8134
rect 36076 8132 36100 8134
rect 36156 8132 36162 8134
rect 35854 8123 36162 8132
rect 35992 7812 36044 7818
rect 35992 7754 36044 7760
rect 36004 7585 36032 7754
rect 36280 7721 36308 8622
rect 36266 7712 36322 7721
rect 36266 7647 36322 7656
rect 35990 7576 36046 7585
rect 35990 7511 36046 7520
rect 36268 7540 36320 7546
rect 36268 7482 36320 7488
rect 35716 7404 35768 7410
rect 35716 7346 35768 7352
rect 35716 7200 35768 7206
rect 35716 7142 35768 7148
rect 35728 6254 35756 7142
rect 35854 7100 36162 7109
rect 35854 7098 35860 7100
rect 35916 7098 35940 7100
rect 35996 7098 36020 7100
rect 36076 7098 36100 7100
rect 36156 7098 36162 7100
rect 35916 7046 35918 7098
rect 36098 7046 36100 7098
rect 35854 7044 35860 7046
rect 35916 7044 35940 7046
rect 35996 7044 36020 7046
rect 36076 7044 36100 7046
rect 36156 7044 36162 7046
rect 35854 7035 36162 7044
rect 35808 6792 35860 6798
rect 35806 6760 35808 6769
rect 35860 6760 35862 6769
rect 36280 6746 36308 7482
rect 36372 7002 36400 8860
rect 36514 8732 36822 8741
rect 36514 8730 36520 8732
rect 36576 8730 36600 8732
rect 36656 8730 36680 8732
rect 36736 8730 36760 8732
rect 36816 8730 36822 8732
rect 36576 8678 36578 8730
rect 36758 8678 36760 8730
rect 36514 8676 36520 8678
rect 36576 8676 36600 8678
rect 36656 8676 36680 8678
rect 36736 8676 36760 8678
rect 36816 8676 36822 8678
rect 36514 8667 36822 8676
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 36740 7750 36768 8434
rect 36728 7744 36780 7750
rect 36728 7686 36780 7692
rect 36514 7644 36822 7653
rect 36514 7642 36520 7644
rect 36576 7642 36600 7644
rect 36656 7642 36680 7644
rect 36736 7642 36760 7644
rect 36816 7642 36822 7644
rect 36576 7590 36578 7642
rect 36758 7590 36760 7642
rect 36514 7588 36520 7590
rect 36576 7588 36600 7590
rect 36656 7588 36680 7590
rect 36736 7588 36760 7590
rect 36816 7588 36822 7590
rect 36514 7579 36822 7588
rect 36360 6996 36412 7002
rect 36360 6938 36412 6944
rect 35806 6695 35862 6704
rect 35992 6724 36044 6730
rect 35992 6666 36044 6672
rect 36188 6718 36308 6746
rect 36360 6724 36412 6730
rect 35900 6656 35952 6662
rect 35898 6624 35900 6633
rect 35952 6624 35954 6633
rect 35898 6559 35954 6568
rect 36004 6458 36032 6666
rect 35992 6452 36044 6458
rect 35992 6394 36044 6400
rect 36188 6322 36216 6718
rect 36360 6666 36412 6672
rect 36372 6458 36400 6666
rect 36514 6556 36822 6565
rect 36514 6554 36520 6556
rect 36576 6554 36600 6556
rect 36656 6554 36680 6556
rect 36736 6554 36760 6556
rect 36816 6554 36822 6556
rect 36576 6502 36578 6554
rect 36758 6502 36760 6554
rect 36514 6500 36520 6502
rect 36576 6500 36600 6502
rect 36656 6500 36680 6502
rect 36736 6500 36760 6502
rect 36816 6500 36822 6502
rect 36514 6491 36822 6500
rect 36360 6452 36412 6458
rect 36360 6394 36412 6400
rect 36924 6338 36952 9998
rect 37096 9444 37148 9450
rect 37096 9386 37148 9392
rect 37004 9376 37056 9382
rect 37004 9318 37056 9324
rect 36176 6316 36228 6322
rect 36176 6258 36228 6264
rect 36268 6316 36320 6322
rect 36268 6258 36320 6264
rect 36372 6310 36952 6338
rect 35716 6248 35768 6254
rect 35716 6190 35768 6196
rect 35714 6080 35770 6089
rect 35714 6015 35770 6024
rect 35728 5914 35756 6015
rect 35854 6012 36162 6021
rect 35854 6010 35860 6012
rect 35916 6010 35940 6012
rect 35996 6010 36020 6012
rect 36076 6010 36100 6012
rect 36156 6010 36162 6012
rect 35916 5958 35918 6010
rect 36098 5958 36100 6010
rect 35854 5956 35860 5958
rect 35916 5956 35940 5958
rect 35996 5956 36020 5958
rect 36076 5956 36100 5958
rect 36156 5956 36162 5958
rect 35854 5947 36162 5956
rect 35716 5908 35768 5914
rect 35716 5850 35768 5856
rect 35992 5908 36044 5914
rect 35992 5850 36044 5856
rect 36004 5710 36032 5850
rect 36280 5846 36308 6258
rect 36268 5840 36320 5846
rect 36268 5782 36320 5788
rect 35992 5704 36044 5710
rect 35992 5646 36044 5652
rect 36176 5704 36228 5710
rect 36176 5646 36228 5652
rect 36084 5228 36136 5234
rect 36188 5216 36216 5646
rect 36268 5636 36320 5642
rect 36268 5578 36320 5584
rect 36136 5188 36216 5216
rect 36084 5170 36136 5176
rect 35854 4924 36162 4933
rect 35854 4922 35860 4924
rect 35916 4922 35940 4924
rect 35996 4922 36020 4924
rect 36076 4922 36100 4924
rect 36156 4922 36162 4924
rect 35916 4870 35918 4922
rect 36098 4870 36100 4922
rect 35854 4868 35860 4870
rect 35916 4868 35940 4870
rect 35996 4868 36020 4870
rect 36076 4868 36100 4870
rect 36156 4868 36162 4870
rect 35854 4859 36162 4868
rect 36280 4826 36308 5578
rect 36084 4820 36136 4826
rect 36268 4820 36320 4826
rect 36136 4780 36216 4808
rect 36084 4762 36136 4768
rect 36084 4548 36136 4554
rect 36084 4490 36136 4496
rect 35714 4176 35770 4185
rect 36096 4146 36124 4490
rect 36188 4146 36216 4780
rect 36268 4762 36320 4768
rect 35714 4111 35770 4120
rect 36084 4140 36136 4146
rect 35728 3738 35756 4111
rect 36084 4082 36136 4088
rect 36176 4140 36228 4146
rect 36176 4082 36228 4088
rect 36188 3890 36216 4082
rect 36188 3862 36308 3890
rect 35854 3836 36162 3845
rect 35854 3834 35860 3836
rect 35916 3834 35940 3836
rect 35996 3834 36020 3836
rect 36076 3834 36100 3836
rect 36156 3834 36162 3836
rect 35916 3782 35918 3834
rect 36098 3782 36100 3834
rect 35854 3780 35860 3782
rect 35916 3780 35940 3782
rect 35996 3780 36020 3782
rect 36076 3780 36100 3782
rect 36156 3780 36162 3782
rect 35854 3771 36162 3780
rect 36280 3754 36308 3862
rect 35716 3732 35768 3738
rect 35716 3674 35768 3680
rect 36188 3726 36308 3754
rect 35716 3460 35768 3466
rect 35716 3402 35768 3408
rect 35624 3120 35676 3126
rect 35624 3062 35676 3068
rect 35532 2848 35584 2854
rect 35532 2790 35584 2796
rect 35360 2746 35480 2774
rect 35256 2440 35308 2446
rect 35256 2382 35308 2388
rect 35452 800 35480 2746
rect 35624 2440 35676 2446
rect 35624 2382 35676 2388
rect 35636 1970 35664 2382
rect 35624 1964 35676 1970
rect 35624 1906 35676 1912
rect 35728 1630 35756 3402
rect 35808 3188 35860 3194
rect 35860 3148 36032 3176
rect 35808 3130 35860 3136
rect 36004 3058 36032 3148
rect 35992 3052 36044 3058
rect 35992 2994 36044 3000
rect 36188 2854 36216 3726
rect 36268 3052 36320 3058
rect 36268 2994 36320 3000
rect 36176 2848 36228 2854
rect 36280 2825 36308 2994
rect 36176 2790 36228 2796
rect 36266 2816 36322 2825
rect 35854 2748 36162 2757
rect 36266 2751 36322 2760
rect 35854 2746 35860 2748
rect 35916 2746 35940 2748
rect 35996 2746 36020 2748
rect 36076 2746 36100 2748
rect 36156 2746 36162 2748
rect 35916 2694 35918 2746
rect 36098 2694 36100 2746
rect 35854 2692 35860 2694
rect 35916 2692 35940 2694
rect 35996 2692 36020 2694
rect 36076 2692 36100 2694
rect 36156 2692 36162 2694
rect 35854 2683 36162 2692
rect 35808 2576 35860 2582
rect 35808 2518 35860 2524
rect 35820 1902 35848 2518
rect 35992 2440 36044 2446
rect 35992 2382 36044 2388
rect 36004 2106 36032 2382
rect 35992 2100 36044 2106
rect 35992 2042 36044 2048
rect 35808 1896 35860 1902
rect 35808 1838 35860 1844
rect 35716 1624 35768 1630
rect 35716 1566 35768 1572
rect 36082 1456 36138 1465
rect 36082 1391 36138 1400
rect 36096 800 36124 1391
rect 34900 734 35112 762
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36372 762 36400 6310
rect 36912 6112 36964 6118
rect 36912 6054 36964 6060
rect 36450 5944 36506 5953
rect 36450 5879 36452 5888
rect 36504 5879 36506 5888
rect 36452 5850 36504 5856
rect 36514 5468 36822 5477
rect 36514 5466 36520 5468
rect 36576 5466 36600 5468
rect 36656 5466 36680 5468
rect 36736 5466 36760 5468
rect 36816 5466 36822 5468
rect 36576 5414 36578 5466
rect 36758 5414 36760 5466
rect 36514 5412 36520 5414
rect 36576 5412 36600 5414
rect 36656 5412 36680 5414
rect 36736 5412 36760 5414
rect 36816 5412 36822 5414
rect 36514 5403 36822 5412
rect 36820 5364 36872 5370
rect 36820 5306 36872 5312
rect 36544 5296 36596 5302
rect 36544 5238 36596 5244
rect 36452 5160 36504 5166
rect 36452 5102 36504 5108
rect 36464 4826 36492 5102
rect 36556 5098 36584 5238
rect 36544 5092 36596 5098
rect 36544 5034 36596 5040
rect 36832 5001 36860 5306
rect 36818 4992 36874 5001
rect 36818 4927 36874 4936
rect 36452 4820 36504 4826
rect 36452 4762 36504 4768
rect 36924 4690 36952 6054
rect 36912 4684 36964 4690
rect 36912 4626 36964 4632
rect 36514 4380 36822 4389
rect 36514 4378 36520 4380
rect 36576 4378 36600 4380
rect 36656 4378 36680 4380
rect 36736 4378 36760 4380
rect 36816 4378 36822 4380
rect 36576 4326 36578 4378
rect 36758 4326 36760 4378
rect 36514 4324 36520 4326
rect 36576 4324 36600 4326
rect 36656 4324 36680 4326
rect 36736 4324 36760 4326
rect 36816 4324 36822 4326
rect 36514 4315 36822 4324
rect 36820 4140 36872 4146
rect 36820 4082 36872 4088
rect 36452 3936 36504 3942
rect 36452 3878 36504 3884
rect 36464 3738 36492 3878
rect 36452 3732 36504 3738
rect 36452 3674 36504 3680
rect 36832 3602 36860 4082
rect 36820 3596 36872 3602
rect 36820 3538 36872 3544
rect 36636 3528 36688 3534
rect 37016 3482 37044 9318
rect 36688 3476 37044 3482
rect 36636 3470 37044 3476
rect 36648 3454 37044 3470
rect 37108 3398 37136 9386
rect 37200 8537 37228 10134
rect 37924 9512 37976 9518
rect 37924 9454 37976 9460
rect 37464 8968 37516 8974
rect 37370 8936 37426 8945
rect 37464 8910 37516 8916
rect 37370 8871 37372 8880
rect 37424 8871 37426 8880
rect 37372 8842 37424 8848
rect 37186 8528 37242 8537
rect 37186 8463 37242 8472
rect 37188 8424 37240 8430
rect 37188 8366 37240 8372
rect 37200 7970 37228 8366
rect 37200 7942 37320 7970
rect 37292 7698 37320 7942
rect 37476 7834 37504 8910
rect 37648 8356 37700 8362
rect 37648 8298 37700 8304
rect 37556 8288 37608 8294
rect 37556 8230 37608 8236
rect 37568 8090 37596 8230
rect 37556 8084 37608 8090
rect 37556 8026 37608 8032
rect 37200 7670 37320 7698
rect 37384 7806 37504 7834
rect 37200 3942 37228 7670
rect 37280 7200 37332 7206
rect 37280 7142 37332 7148
rect 37292 6254 37320 7142
rect 37280 6248 37332 6254
rect 37280 6190 37332 6196
rect 37280 5772 37332 5778
rect 37280 5714 37332 5720
rect 37292 5681 37320 5714
rect 37278 5672 37334 5681
rect 37278 5607 37334 5616
rect 37280 4072 37332 4078
rect 37280 4014 37332 4020
rect 37188 3936 37240 3942
rect 37188 3878 37240 3884
rect 37096 3392 37148 3398
rect 37096 3334 37148 3340
rect 36514 3292 36822 3301
rect 36514 3290 36520 3292
rect 36576 3290 36600 3292
rect 36656 3290 36680 3292
rect 36736 3290 36760 3292
rect 36816 3290 36822 3292
rect 36576 3238 36578 3290
rect 36758 3238 36760 3290
rect 36514 3236 36520 3238
rect 36576 3236 36600 3238
rect 36656 3236 36680 3238
rect 36736 3236 36760 3238
rect 36816 3236 36822 3238
rect 36514 3227 36822 3236
rect 36910 2952 36966 2961
rect 36910 2887 36966 2896
rect 36514 2204 36822 2213
rect 36514 2202 36520 2204
rect 36576 2202 36600 2204
rect 36656 2202 36680 2204
rect 36736 2202 36760 2204
rect 36816 2202 36822 2204
rect 36576 2150 36578 2202
rect 36758 2150 36760 2202
rect 36514 2148 36520 2150
rect 36576 2148 36600 2150
rect 36656 2148 36680 2150
rect 36736 2148 36760 2150
rect 36816 2148 36822 2150
rect 36514 2139 36822 2148
rect 36924 1698 36952 2887
rect 36912 1692 36964 1698
rect 36912 1634 36964 1640
rect 37292 1465 37320 4014
rect 37278 1456 37334 1465
rect 37278 1391 37334 1400
rect 36648 870 36768 898
rect 36648 762 36676 870
rect 36740 800 36768 870
rect 37384 800 37412 7806
rect 37464 7744 37516 7750
rect 37464 7686 37516 7692
rect 37476 7410 37504 7686
rect 37464 7404 37516 7410
rect 37464 7346 37516 7352
rect 37464 7268 37516 7274
rect 37464 7210 37516 7216
rect 37476 4826 37504 7210
rect 37556 6180 37608 6186
rect 37556 6122 37608 6128
rect 37568 5914 37596 6122
rect 37556 5908 37608 5914
rect 37556 5850 37608 5856
rect 37556 5228 37608 5234
rect 37556 5170 37608 5176
rect 37568 5001 37596 5170
rect 37554 4992 37610 5001
rect 37554 4927 37610 4936
rect 37464 4820 37516 4826
rect 37464 4762 37516 4768
rect 37556 4480 37608 4486
rect 37556 4422 37608 4428
rect 37568 3126 37596 4422
rect 37660 3126 37688 8298
rect 37830 6488 37886 6497
rect 37830 6423 37886 6432
rect 37844 6322 37872 6423
rect 37832 6316 37884 6322
rect 37832 6258 37884 6264
rect 37830 6216 37886 6225
rect 37830 6151 37886 6160
rect 37844 5710 37872 6151
rect 37832 5704 37884 5710
rect 37832 5646 37884 5652
rect 37832 5568 37884 5574
rect 37832 5510 37884 5516
rect 37740 5296 37792 5302
rect 37740 5238 37792 5244
rect 37752 5098 37780 5238
rect 37740 5092 37792 5098
rect 37740 5034 37792 5040
rect 37738 4720 37794 4729
rect 37738 4655 37794 4664
rect 37752 4622 37780 4655
rect 37844 4622 37872 5510
rect 37936 5137 37964 9454
rect 37922 5128 37978 5137
rect 37922 5063 37978 5072
rect 37924 5024 37976 5030
rect 37924 4966 37976 4972
rect 37936 4826 37964 4966
rect 37924 4820 37976 4826
rect 37924 4762 37976 4768
rect 37740 4616 37792 4622
rect 37740 4558 37792 4564
rect 37832 4616 37884 4622
rect 37832 4558 37884 4564
rect 37844 3194 37872 4558
rect 37922 3632 37978 3641
rect 37922 3567 37978 3576
rect 37936 3466 37964 3567
rect 37924 3460 37976 3466
rect 37924 3402 37976 3408
rect 37832 3188 37884 3194
rect 37832 3130 37884 3136
rect 37556 3120 37608 3126
rect 37556 3062 37608 3068
rect 37648 3120 37700 3126
rect 37648 3062 37700 3068
rect 37568 2825 37596 3062
rect 37554 2816 37610 2825
rect 37554 2751 37610 2760
rect 38028 2446 38056 12582
rect 66574 12540 66882 12549
rect 66574 12538 66580 12540
rect 66636 12538 66660 12540
rect 66716 12538 66740 12540
rect 66796 12538 66820 12540
rect 66876 12538 66882 12540
rect 66636 12486 66638 12538
rect 66818 12486 66820 12538
rect 66574 12484 66580 12486
rect 66636 12484 66660 12486
rect 66716 12484 66740 12486
rect 66796 12484 66820 12486
rect 66876 12484 66882 12486
rect 66574 12475 66882 12484
rect 67234 11996 67542 12005
rect 67234 11994 67240 11996
rect 67296 11994 67320 11996
rect 67376 11994 67400 11996
rect 67456 11994 67480 11996
rect 67536 11994 67542 11996
rect 67296 11942 67298 11994
rect 67478 11942 67480 11994
rect 67234 11940 67240 11942
rect 67296 11940 67320 11942
rect 67376 11940 67400 11942
rect 67456 11940 67480 11942
rect 67536 11940 67542 11942
rect 67234 11931 67542 11940
rect 38844 11620 38896 11626
rect 38844 11562 38896 11568
rect 38752 9920 38804 9926
rect 38752 9862 38804 9868
rect 38764 9586 38792 9862
rect 38752 9580 38804 9586
rect 38752 9522 38804 9528
rect 38200 9376 38252 9382
rect 38200 9318 38252 9324
rect 38212 7993 38240 9318
rect 38292 9036 38344 9042
rect 38292 8978 38344 8984
rect 38198 7984 38254 7993
rect 38198 7919 38254 7928
rect 38200 7880 38252 7886
rect 38200 7822 38252 7828
rect 38212 6866 38240 7822
rect 38200 6860 38252 6866
rect 38200 6802 38252 6808
rect 38106 6760 38162 6769
rect 38106 6695 38162 6704
rect 38120 4808 38148 6695
rect 38212 6322 38240 6802
rect 38200 6316 38252 6322
rect 38200 6258 38252 6264
rect 38212 5574 38240 6258
rect 38200 5568 38252 5574
rect 38200 5510 38252 5516
rect 38120 4780 38240 4808
rect 38212 4146 38240 4780
rect 38200 4140 38252 4146
rect 38200 4082 38252 4088
rect 38108 4072 38160 4078
rect 38108 4014 38160 4020
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 38120 1442 38148 4014
rect 38304 1873 38332 8978
rect 38660 8832 38712 8838
rect 38660 8774 38712 8780
rect 38672 8401 38700 8774
rect 38658 8392 38714 8401
rect 38658 8327 38714 8336
rect 38384 7812 38436 7818
rect 38384 7754 38436 7760
rect 38396 6730 38424 7754
rect 38568 7404 38620 7410
rect 38568 7346 38620 7352
rect 38384 6724 38436 6730
rect 38384 6666 38436 6672
rect 38396 6390 38424 6666
rect 38580 6633 38608 7346
rect 38566 6624 38622 6633
rect 38566 6559 38622 6568
rect 38474 6488 38530 6497
rect 38614 6452 38666 6458
rect 38530 6432 38614 6440
rect 38474 6423 38614 6432
rect 38488 6412 38614 6423
rect 38614 6394 38666 6400
rect 38384 6384 38436 6390
rect 38384 6326 38436 6332
rect 38568 6248 38620 6254
rect 38474 6216 38530 6225
rect 38568 6190 38620 6196
rect 38474 6151 38530 6160
rect 38384 4548 38436 4554
rect 38384 4490 38436 4496
rect 38396 2990 38424 4490
rect 38488 3194 38516 6151
rect 38580 5953 38608 6190
rect 38566 5944 38622 5953
rect 38566 5879 38622 5888
rect 38660 5908 38712 5914
rect 38660 5850 38712 5856
rect 38568 5704 38620 5710
rect 38568 5646 38620 5652
rect 38580 4146 38608 5646
rect 38672 5166 38700 5850
rect 38660 5160 38712 5166
rect 38660 5102 38712 5108
rect 38568 4140 38620 4146
rect 38568 4082 38620 4088
rect 38660 4140 38712 4146
rect 38660 4082 38712 4088
rect 38672 3602 38700 4082
rect 38660 3596 38712 3602
rect 38660 3538 38712 3544
rect 38658 3496 38714 3505
rect 38658 3431 38714 3440
rect 38476 3188 38528 3194
rect 38476 3130 38528 3136
rect 38384 2984 38436 2990
rect 38384 2926 38436 2932
rect 38290 1864 38346 1873
rect 38290 1799 38346 1808
rect 38028 1414 38148 1442
rect 38028 800 38056 1414
rect 38672 800 38700 3431
rect 38752 3392 38804 3398
rect 38752 3334 38804 3340
rect 38764 2378 38792 3334
rect 38856 2446 38884 11562
rect 66574 11452 66882 11461
rect 66574 11450 66580 11452
rect 66636 11450 66660 11452
rect 66716 11450 66740 11452
rect 66796 11450 66820 11452
rect 66876 11450 66882 11452
rect 66636 11398 66638 11450
rect 66818 11398 66820 11450
rect 66574 11396 66580 11398
rect 66636 11396 66660 11398
rect 66716 11396 66740 11398
rect 66796 11396 66820 11398
rect 66876 11396 66882 11398
rect 66574 11387 66882 11396
rect 67234 10908 67542 10917
rect 67234 10906 67240 10908
rect 67296 10906 67320 10908
rect 67376 10906 67400 10908
rect 67456 10906 67480 10908
rect 67536 10906 67542 10908
rect 67296 10854 67298 10906
rect 67478 10854 67480 10906
rect 67234 10852 67240 10854
rect 67296 10852 67320 10854
rect 67376 10852 67400 10854
rect 67456 10852 67480 10854
rect 67536 10852 67542 10854
rect 67234 10843 67542 10852
rect 66574 10364 66882 10373
rect 66574 10362 66580 10364
rect 66636 10362 66660 10364
rect 66716 10362 66740 10364
rect 66796 10362 66820 10364
rect 66876 10362 66882 10364
rect 66636 10310 66638 10362
rect 66818 10310 66820 10362
rect 66574 10308 66580 10310
rect 66636 10308 66660 10310
rect 66716 10308 66740 10310
rect 66796 10308 66820 10310
rect 66876 10308 66882 10310
rect 66574 10299 66882 10308
rect 67234 9820 67542 9829
rect 67234 9818 67240 9820
rect 67296 9818 67320 9820
rect 67376 9818 67400 9820
rect 67456 9818 67480 9820
rect 67536 9818 67542 9820
rect 67296 9766 67298 9818
rect 67478 9766 67480 9818
rect 67234 9764 67240 9766
rect 67296 9764 67320 9766
rect 67376 9764 67400 9766
rect 67456 9764 67480 9766
rect 67536 9764 67542 9766
rect 67234 9755 67542 9764
rect 66574 9276 66882 9285
rect 66574 9274 66580 9276
rect 66636 9274 66660 9276
rect 66716 9274 66740 9276
rect 66796 9274 66820 9276
rect 66876 9274 66882 9276
rect 66636 9222 66638 9274
rect 66818 9222 66820 9274
rect 66574 9220 66580 9222
rect 66636 9220 66660 9222
rect 66716 9220 66740 9222
rect 66796 9220 66820 9222
rect 66876 9220 66882 9222
rect 66574 9211 66882 9220
rect 67234 8732 67542 8741
rect 67234 8730 67240 8732
rect 67296 8730 67320 8732
rect 67376 8730 67400 8732
rect 67456 8730 67480 8732
rect 67536 8730 67542 8732
rect 67296 8678 67298 8730
rect 67478 8678 67480 8730
rect 67234 8676 67240 8678
rect 67296 8676 67320 8678
rect 67376 8676 67400 8678
rect 67456 8676 67480 8678
rect 67536 8676 67542 8678
rect 67234 8667 67542 8676
rect 39304 8424 39356 8430
rect 39304 8366 39356 8372
rect 39212 7744 39264 7750
rect 39212 7686 39264 7692
rect 39120 6656 39172 6662
rect 39120 6598 39172 6604
rect 38936 6384 38988 6390
rect 38934 6352 38936 6361
rect 38988 6352 38990 6361
rect 38934 6287 38990 6296
rect 39132 5778 39160 6598
rect 39120 5772 39172 5778
rect 39120 5714 39172 5720
rect 39028 5568 39080 5574
rect 39028 5510 39080 5516
rect 39040 5166 39068 5510
rect 39028 5160 39080 5166
rect 39028 5102 39080 5108
rect 38936 3936 38988 3942
rect 38936 3878 38988 3884
rect 38948 3670 38976 3878
rect 38936 3664 38988 3670
rect 38936 3606 38988 3612
rect 38844 2440 38896 2446
rect 38844 2382 38896 2388
rect 38936 2440 38988 2446
rect 38936 2382 38988 2388
rect 38752 2372 38804 2378
rect 38752 2314 38804 2320
rect 38948 2038 38976 2382
rect 38936 2032 38988 2038
rect 38936 1974 38988 1980
rect 39224 1834 39252 7686
rect 39212 1828 39264 1834
rect 39212 1770 39264 1776
rect 39316 800 39344 8366
rect 41420 8356 41472 8362
rect 41420 8298 41472 8304
rect 40408 7948 40460 7954
rect 40408 7890 40460 7896
rect 40132 7744 40184 7750
rect 40132 7686 40184 7692
rect 39394 6896 39450 6905
rect 39394 6831 39396 6840
rect 39448 6831 39450 6840
rect 39396 6802 39448 6808
rect 39408 5710 39436 6802
rect 39580 6724 39632 6730
rect 39580 6666 39632 6672
rect 39486 6352 39542 6361
rect 39486 6287 39542 6296
rect 39396 5704 39448 5710
rect 39396 5646 39448 5652
rect 39500 4554 39528 6287
rect 39592 5914 39620 6666
rect 39856 6112 39908 6118
rect 39856 6054 39908 6060
rect 39580 5908 39632 5914
rect 39580 5850 39632 5856
rect 39868 5370 39896 6054
rect 39764 5364 39816 5370
rect 39764 5306 39816 5312
rect 39856 5364 39908 5370
rect 39856 5306 39908 5312
rect 39488 4548 39540 4554
rect 39488 4490 39540 4496
rect 39776 3602 39804 5306
rect 39868 4690 39896 5306
rect 40144 5302 40172 7686
rect 40224 6860 40276 6866
rect 40224 6802 40276 6808
rect 40236 6254 40264 6802
rect 40224 6248 40276 6254
rect 40224 6190 40276 6196
rect 40236 5817 40264 6190
rect 40222 5808 40278 5817
rect 40222 5743 40278 5752
rect 40132 5296 40184 5302
rect 40132 5238 40184 5244
rect 39948 5024 40000 5030
rect 39948 4966 40000 4972
rect 39960 4690 39988 4966
rect 39856 4684 39908 4690
rect 39856 4626 39908 4632
rect 39948 4684 40000 4690
rect 39948 4626 40000 4632
rect 40040 4548 40092 4554
rect 40040 4490 40092 4496
rect 40132 4548 40184 4554
rect 40132 4490 40184 4496
rect 40052 4214 40080 4490
rect 39948 4208 40000 4214
rect 39948 4150 40000 4156
rect 40040 4208 40092 4214
rect 40040 4150 40092 4156
rect 39764 3596 39816 3602
rect 39764 3538 39816 3544
rect 39960 3398 39988 4150
rect 39948 3392 40000 3398
rect 39948 3334 40000 3340
rect 40052 3058 40080 4150
rect 40040 3052 40092 3058
rect 40040 2994 40092 3000
rect 40144 2774 40172 4490
rect 40316 3732 40368 3738
rect 40316 3674 40368 3680
rect 40328 3534 40356 3674
rect 40316 3528 40368 3534
rect 40316 3470 40368 3476
rect 40328 2990 40356 3470
rect 40316 2984 40368 2990
rect 40316 2926 40368 2932
rect 40052 2746 40172 2774
rect 40420 2774 40448 7890
rect 40868 7812 40920 7818
rect 40868 7754 40920 7760
rect 40500 7744 40552 7750
rect 40500 7686 40552 7692
rect 40512 6390 40540 7686
rect 40684 7200 40736 7206
rect 40684 7142 40736 7148
rect 40592 6656 40644 6662
rect 40592 6598 40644 6604
rect 40604 6458 40632 6598
rect 40592 6452 40644 6458
rect 40592 6394 40644 6400
rect 40500 6384 40552 6390
rect 40500 6326 40552 6332
rect 40500 5568 40552 5574
rect 40500 5510 40552 5516
rect 40512 5234 40540 5510
rect 40500 5228 40552 5234
rect 40500 5170 40552 5176
rect 40420 2746 40540 2774
rect 40052 2514 40080 2746
rect 39856 2508 39908 2514
rect 39856 2450 39908 2456
rect 40040 2508 40092 2514
rect 40040 2450 40092 2456
rect 39868 1170 39896 2450
rect 40512 1902 40540 2746
rect 40696 1970 40724 7142
rect 40880 6458 40908 7754
rect 41432 7410 41460 8298
rect 66574 8188 66882 8197
rect 66574 8186 66580 8188
rect 66636 8186 66660 8188
rect 66716 8186 66740 8188
rect 66796 8186 66820 8188
rect 66876 8186 66882 8188
rect 66636 8134 66638 8186
rect 66818 8134 66820 8186
rect 66574 8132 66580 8134
rect 66636 8132 66660 8134
rect 66716 8132 66740 8134
rect 66796 8132 66820 8134
rect 66876 8132 66882 8134
rect 66574 8123 66882 8132
rect 41604 7880 41656 7886
rect 41604 7822 41656 7828
rect 41420 7404 41472 7410
rect 41420 7346 41472 7352
rect 41420 6656 41472 6662
rect 41420 6598 41472 6604
rect 41512 6656 41564 6662
rect 41512 6598 41564 6604
rect 40868 6452 40920 6458
rect 40868 6394 40920 6400
rect 40880 5642 40908 6394
rect 41432 6322 41460 6598
rect 41420 6316 41472 6322
rect 41420 6258 41472 6264
rect 41328 6248 41380 6254
rect 41328 6190 41380 6196
rect 41144 6112 41196 6118
rect 41144 6054 41196 6060
rect 41156 5778 41184 6054
rect 41144 5772 41196 5778
rect 41144 5714 41196 5720
rect 40868 5636 40920 5642
rect 40868 5578 40920 5584
rect 41340 4758 41368 6190
rect 41420 5840 41472 5846
rect 41420 5782 41472 5788
rect 41328 4752 41380 4758
rect 41328 4694 41380 4700
rect 40960 4548 41012 4554
rect 40960 4490 41012 4496
rect 40972 4282 41000 4490
rect 40960 4276 41012 4282
rect 40960 4218 41012 4224
rect 41328 4276 41380 4282
rect 41328 4218 41380 4224
rect 40972 3058 41000 4218
rect 41144 3392 41196 3398
rect 41144 3334 41196 3340
rect 41236 3392 41288 3398
rect 41236 3334 41288 3340
rect 41156 3194 41184 3334
rect 41144 3188 41196 3194
rect 41144 3130 41196 3136
rect 40960 3052 41012 3058
rect 40960 2994 41012 3000
rect 41156 2514 41184 3130
rect 41144 2508 41196 2514
rect 41144 2450 41196 2456
rect 40684 1964 40736 1970
rect 40684 1906 40736 1912
rect 40500 1896 40552 1902
rect 40500 1838 40552 1844
rect 41248 1766 41276 3334
rect 41236 1760 41288 1766
rect 41236 1702 41288 1708
rect 41340 1170 41368 4218
rect 41432 2922 41460 5782
rect 41420 2916 41472 2922
rect 41420 2858 41472 2864
rect 41524 2774 41552 6598
rect 41616 5914 41644 7822
rect 67234 7644 67542 7653
rect 67234 7642 67240 7644
rect 67296 7642 67320 7644
rect 67376 7642 67400 7644
rect 67456 7642 67480 7644
rect 67536 7642 67542 7644
rect 67296 7590 67298 7642
rect 67478 7590 67480 7642
rect 67234 7588 67240 7590
rect 67296 7588 67320 7590
rect 67376 7588 67400 7590
rect 67456 7588 67480 7590
rect 67536 7588 67542 7590
rect 67234 7579 67542 7588
rect 66574 7100 66882 7109
rect 66574 7098 66580 7100
rect 66636 7098 66660 7100
rect 66716 7098 66740 7100
rect 66796 7098 66820 7100
rect 66876 7098 66882 7100
rect 66636 7046 66638 7098
rect 66818 7046 66820 7098
rect 66574 7044 66580 7046
rect 66636 7044 66660 7046
rect 66716 7044 66740 7046
rect 66796 7044 66820 7046
rect 66876 7044 66882 7046
rect 66574 7035 66882 7044
rect 44088 6792 44140 6798
rect 44088 6734 44140 6740
rect 43352 6724 43404 6730
rect 43352 6666 43404 6672
rect 41788 6656 41840 6662
rect 41788 6598 41840 6604
rect 41604 5908 41656 5914
rect 41604 5850 41656 5856
rect 41800 5710 41828 6598
rect 42524 6384 42576 6390
rect 42524 6326 42576 6332
rect 41972 6248 42024 6254
rect 41972 6190 42024 6196
rect 41788 5704 41840 5710
rect 41788 5646 41840 5652
rect 41696 5568 41748 5574
rect 41696 5510 41748 5516
rect 41604 5364 41656 5370
rect 41604 5306 41656 5312
rect 41616 5166 41644 5306
rect 41604 5160 41656 5166
rect 41604 5102 41656 5108
rect 41604 4208 41656 4214
rect 41604 4150 41656 4156
rect 41616 4078 41644 4150
rect 41708 4078 41736 5510
rect 41788 4616 41840 4622
rect 41788 4558 41840 4564
rect 41604 4072 41656 4078
rect 41604 4014 41656 4020
rect 41696 4072 41748 4078
rect 41696 4014 41748 4020
rect 41696 3460 41748 3466
rect 41696 3402 41748 3408
rect 41708 3194 41736 3402
rect 41696 3188 41748 3194
rect 41696 3130 41748 3136
rect 41524 2746 41644 2774
rect 41616 2650 41644 2746
rect 41604 2644 41656 2650
rect 41604 2586 41656 2592
rect 41800 2417 41828 4558
rect 41984 2582 42012 6190
rect 42064 5704 42116 5710
rect 42064 5646 42116 5652
rect 42076 5370 42104 5646
rect 42536 5370 42564 6326
rect 43076 6316 43128 6322
rect 43076 6258 43128 6264
rect 42616 6112 42668 6118
rect 42616 6054 42668 6060
rect 42800 6112 42852 6118
rect 42800 6054 42852 6060
rect 42628 5778 42656 6054
rect 42616 5772 42668 5778
rect 42616 5714 42668 5720
rect 42064 5364 42116 5370
rect 42064 5306 42116 5312
rect 42524 5364 42576 5370
rect 42524 5306 42576 5312
rect 42156 5296 42208 5302
rect 42156 5238 42208 5244
rect 42064 5160 42116 5166
rect 42064 5102 42116 5108
rect 42076 3534 42104 5102
rect 42064 3528 42116 3534
rect 42064 3470 42116 3476
rect 42168 2990 42196 5238
rect 42616 4616 42668 4622
rect 42616 4558 42668 4564
rect 42248 4480 42300 4486
rect 42248 4422 42300 4428
rect 42260 4214 42288 4422
rect 42628 4214 42656 4558
rect 42248 4208 42300 4214
rect 42248 4150 42300 4156
rect 42616 4208 42668 4214
rect 42616 4150 42668 4156
rect 42812 4078 42840 6054
rect 42984 5704 43036 5710
rect 42984 5646 43036 5652
rect 42892 5092 42944 5098
rect 42892 5034 42944 5040
rect 42800 4072 42852 4078
rect 42800 4014 42852 4020
rect 42248 4004 42300 4010
rect 42248 3946 42300 3952
rect 42260 3602 42288 3946
rect 42904 3942 42932 5034
rect 42892 3936 42944 3942
rect 42892 3878 42944 3884
rect 42996 3618 43024 5646
rect 43088 5234 43116 6258
rect 43168 5704 43220 5710
rect 43168 5646 43220 5652
rect 43076 5228 43128 5234
rect 43076 5170 43128 5176
rect 43076 5024 43128 5030
rect 43076 4966 43128 4972
rect 43088 4758 43116 4966
rect 43076 4752 43128 4758
rect 43076 4694 43128 4700
rect 43076 4616 43128 4622
rect 43076 4558 43128 4564
rect 43088 4078 43116 4558
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 42248 3596 42300 3602
rect 42248 3538 42300 3544
rect 42812 3590 43024 3618
rect 42260 3176 42288 3538
rect 42812 3466 42840 3590
rect 42800 3460 42852 3466
rect 42800 3402 42852 3408
rect 42984 3460 43036 3466
rect 42984 3402 43036 3408
rect 42340 3188 42392 3194
rect 42260 3148 42340 3176
rect 42340 3130 42392 3136
rect 42996 3126 43024 3402
rect 42984 3120 43036 3126
rect 42982 3088 42984 3097
rect 43036 3088 43038 3097
rect 42982 3023 43038 3032
rect 42156 2984 42208 2990
rect 42156 2926 42208 2932
rect 42800 2848 42852 2854
rect 42720 2796 42800 2802
rect 42720 2790 42852 2796
rect 42720 2774 42840 2790
rect 41972 2576 42024 2582
rect 41972 2518 42024 2524
rect 41880 2508 41932 2514
rect 41880 2450 41932 2456
rect 41786 2408 41842 2417
rect 41786 2343 41842 2352
rect 39868 1142 39988 1170
rect 39960 800 39988 1142
rect 40592 1148 40644 1154
rect 40592 1090 40644 1096
rect 41248 1142 41368 1170
rect 40604 800 40632 1090
rect 41248 800 41276 1142
rect 41892 800 41920 2450
rect 42720 2378 42748 2774
rect 42708 2372 42760 2378
rect 42708 2314 42760 2320
rect 42524 1352 42576 1358
rect 42524 1294 42576 1300
rect 42536 800 42564 1294
rect 43180 800 43208 5646
rect 43364 4690 43392 6666
rect 43536 5228 43588 5234
rect 43536 5170 43588 5176
rect 43352 4684 43404 4690
rect 43352 4626 43404 4632
rect 43260 4480 43312 4486
rect 43260 4422 43312 4428
rect 43352 4480 43404 4486
rect 43352 4422 43404 4428
rect 43272 4010 43300 4422
rect 43260 4004 43312 4010
rect 43260 3946 43312 3952
rect 43364 3058 43392 4422
rect 43548 3942 43576 5170
rect 44100 4690 44128 6734
rect 67234 6556 67542 6565
rect 67234 6554 67240 6556
rect 67296 6554 67320 6556
rect 67376 6554 67400 6556
rect 67456 6554 67480 6556
rect 67536 6554 67542 6556
rect 67296 6502 67298 6554
rect 67478 6502 67480 6554
rect 67234 6500 67240 6502
rect 67296 6500 67320 6502
rect 67376 6500 67400 6502
rect 67456 6500 67480 6502
rect 67536 6500 67542 6502
rect 67234 6491 67542 6500
rect 66574 6012 66882 6021
rect 66574 6010 66580 6012
rect 66636 6010 66660 6012
rect 66716 6010 66740 6012
rect 66796 6010 66820 6012
rect 66876 6010 66882 6012
rect 66636 5958 66638 6010
rect 66818 5958 66820 6010
rect 66574 5956 66580 5958
rect 66636 5956 66660 5958
rect 66716 5956 66740 5958
rect 66796 5956 66820 5958
rect 66876 5956 66882 5958
rect 66574 5947 66882 5956
rect 45928 5704 45980 5710
rect 45928 5646 45980 5652
rect 48780 5704 48832 5710
rect 48780 5646 48832 5652
rect 44272 5568 44324 5574
rect 44272 5510 44324 5516
rect 44284 5234 44312 5510
rect 44914 5264 44970 5273
rect 44272 5228 44324 5234
rect 44914 5199 44970 5208
rect 44272 5170 44324 5176
rect 44640 5160 44692 5166
rect 44640 5102 44692 5108
rect 44732 5160 44784 5166
rect 44732 5102 44784 5108
rect 44088 4684 44140 4690
rect 44088 4626 44140 4632
rect 44180 4616 44232 4622
rect 44180 4558 44232 4564
rect 44192 4282 44220 4558
rect 44180 4276 44232 4282
rect 44180 4218 44232 4224
rect 43812 4072 43864 4078
rect 43812 4014 43864 4020
rect 43536 3936 43588 3942
rect 43536 3878 43588 3884
rect 43824 3126 43852 4014
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 44284 3398 44312 3538
rect 44272 3392 44324 3398
rect 44272 3334 44324 3340
rect 43812 3120 43864 3126
rect 43812 3062 43864 3068
rect 43352 3052 43404 3058
rect 43352 2994 43404 3000
rect 43536 2848 43588 2854
rect 43536 2790 43588 2796
rect 43548 2650 43576 2790
rect 43536 2644 43588 2650
rect 43536 2586 43588 2592
rect 44284 2514 44312 3334
rect 44652 2582 44680 5102
rect 44744 2650 44772 5102
rect 44928 4078 44956 5199
rect 45836 5024 45888 5030
rect 45836 4966 45888 4972
rect 45192 4684 45244 4690
rect 45192 4626 45244 4632
rect 44824 4072 44876 4078
rect 44824 4014 44876 4020
rect 44916 4072 44968 4078
rect 44916 4014 44968 4020
rect 44836 3194 44864 4014
rect 44916 3392 44968 3398
rect 44916 3334 44968 3340
rect 44824 3188 44876 3194
rect 44824 3130 44876 3136
rect 44732 2644 44784 2650
rect 44732 2586 44784 2592
rect 44640 2576 44692 2582
rect 44640 2518 44692 2524
rect 44272 2508 44324 2514
rect 44272 2450 44324 2456
rect 44836 2446 44864 3130
rect 44928 2990 44956 3334
rect 45100 3120 45152 3126
rect 45100 3062 45152 3068
rect 44916 2984 44968 2990
rect 44916 2926 44968 2932
rect 44824 2440 44876 2446
rect 44824 2382 44876 2388
rect 43812 2372 43864 2378
rect 43812 2314 43864 2320
rect 43824 800 43852 2314
rect 44456 2032 44508 2038
rect 44456 1974 44508 1980
rect 44468 800 44496 1974
rect 45112 800 45140 3062
rect 45204 1154 45232 4626
rect 45468 4548 45520 4554
rect 45468 4490 45520 4496
rect 45652 4548 45704 4554
rect 45652 4490 45704 4496
rect 45376 4208 45428 4214
rect 45376 4150 45428 4156
rect 45388 3194 45416 4150
rect 45376 3188 45428 3194
rect 45376 3130 45428 3136
rect 45480 2922 45508 4490
rect 45560 4480 45612 4486
rect 45560 4422 45612 4428
rect 45572 3602 45600 4422
rect 45560 3596 45612 3602
rect 45560 3538 45612 3544
rect 45664 3058 45692 4490
rect 45744 3596 45796 3602
rect 45744 3538 45796 3544
rect 45652 3052 45704 3058
rect 45652 2994 45704 3000
rect 45468 2916 45520 2922
rect 45468 2858 45520 2864
rect 45192 1148 45244 1154
rect 45192 1090 45244 1096
rect 45756 800 45784 3538
rect 45848 3058 45876 4966
rect 45940 3194 45968 5646
rect 46940 5568 46992 5574
rect 46940 5510 46992 5516
rect 46952 5234 46980 5510
rect 46940 5228 46992 5234
rect 46940 5170 46992 5176
rect 46296 5024 46348 5030
rect 46296 4966 46348 4972
rect 46112 3936 46164 3942
rect 46112 3878 46164 3884
rect 45928 3188 45980 3194
rect 45928 3130 45980 3136
rect 46124 3058 46152 3878
rect 46308 3534 46336 4966
rect 47032 4820 47084 4826
rect 47032 4762 47084 4768
rect 46940 4072 46992 4078
rect 46940 4014 46992 4020
rect 46388 3936 46440 3942
rect 46388 3878 46440 3884
rect 46400 3670 46428 3878
rect 46952 3738 46980 4014
rect 46940 3732 46992 3738
rect 46940 3674 46992 3680
rect 46388 3664 46440 3670
rect 46388 3606 46440 3612
rect 46296 3528 46348 3534
rect 46296 3470 46348 3476
rect 46480 3528 46532 3534
rect 46480 3470 46532 3476
rect 46664 3528 46716 3534
rect 46664 3470 46716 3476
rect 46940 3528 46992 3534
rect 46940 3470 46992 3476
rect 45836 3052 45888 3058
rect 45836 2994 45888 3000
rect 46112 3052 46164 3058
rect 46112 2994 46164 3000
rect 46492 2990 46520 3470
rect 45928 2984 45980 2990
rect 45928 2926 45980 2932
rect 46480 2984 46532 2990
rect 46480 2926 46532 2932
rect 45836 2644 45888 2650
rect 45836 2586 45888 2592
rect 45848 2446 45876 2586
rect 45940 2446 45968 2926
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 45928 2440 45980 2446
rect 45928 2382 45980 2388
rect 46400 870 46520 898
rect 46400 800 46428 870
rect 36372 734 36676 762
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 46492 762 46520 870
rect 46676 762 46704 3470
rect 46848 3460 46900 3466
rect 46848 3402 46900 3408
rect 46860 2650 46888 3402
rect 46952 3126 46980 3470
rect 46940 3120 46992 3126
rect 46940 3062 46992 3068
rect 46848 2644 46900 2650
rect 46848 2586 46900 2592
rect 47044 2514 47072 4762
rect 47216 4684 47268 4690
rect 47216 4626 47268 4632
rect 47228 4078 47256 4626
rect 48044 4616 48096 4622
rect 48044 4558 48096 4564
rect 47124 4072 47176 4078
rect 47124 4014 47176 4020
rect 47216 4072 47268 4078
rect 47216 4014 47268 4020
rect 47032 2508 47084 2514
rect 47032 2450 47084 2456
rect 47136 1358 47164 4014
rect 47492 3936 47544 3942
rect 47492 3878 47544 3884
rect 47504 3058 47532 3878
rect 48056 3194 48084 4558
rect 48320 4480 48372 4486
rect 48320 4422 48372 4428
rect 48044 3188 48096 3194
rect 48044 3130 48096 3136
rect 47492 3052 47544 3058
rect 47492 2994 47544 3000
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47400 2304 47452 2310
rect 47400 2246 47452 2252
rect 47412 2106 47440 2246
rect 47400 2100 47452 2106
rect 47400 2042 47452 2048
rect 47124 1352 47176 1358
rect 47124 1294 47176 1300
rect 47688 800 47716 2926
rect 48332 2446 48360 4422
rect 48596 4072 48648 4078
rect 48596 4014 48648 4020
rect 48608 3398 48636 4014
rect 48792 3738 48820 5646
rect 49792 5636 49844 5642
rect 49792 5578 49844 5584
rect 48872 4616 48924 4622
rect 48872 4558 48924 4564
rect 48884 4010 48912 4558
rect 48872 4004 48924 4010
rect 48872 3946 48924 3952
rect 49240 3936 49292 3942
rect 49240 3878 49292 3884
rect 48780 3732 48832 3738
rect 48780 3674 48832 3680
rect 48596 3392 48648 3398
rect 48596 3334 48648 3340
rect 49252 3058 49280 3878
rect 49804 3534 49832 5578
rect 67234 5468 67542 5477
rect 67234 5466 67240 5468
rect 67296 5466 67320 5468
rect 67376 5466 67400 5468
rect 67456 5466 67480 5468
rect 67536 5466 67542 5468
rect 67296 5414 67298 5466
rect 67478 5414 67480 5466
rect 67234 5412 67240 5414
rect 67296 5412 67320 5414
rect 67376 5412 67400 5414
rect 67456 5412 67480 5414
rect 67536 5412 67542 5414
rect 67234 5403 67542 5412
rect 76932 5160 76984 5166
rect 76932 5102 76984 5108
rect 76656 5024 76708 5030
rect 76656 4966 76708 4972
rect 66574 4924 66882 4933
rect 66574 4922 66580 4924
rect 66636 4922 66660 4924
rect 66716 4922 66740 4924
rect 66796 4922 66820 4924
rect 66876 4922 66882 4924
rect 66636 4870 66638 4922
rect 66818 4870 66820 4922
rect 66574 4868 66580 4870
rect 66636 4868 66660 4870
rect 66716 4868 66740 4870
rect 66796 4868 66820 4870
rect 66876 4868 66882 4870
rect 66574 4859 66882 4868
rect 51078 4720 51134 4729
rect 51078 4655 51134 4664
rect 49976 4548 50028 4554
rect 49976 4490 50028 4496
rect 49884 3936 49936 3942
rect 49884 3878 49936 3884
rect 49792 3528 49844 3534
rect 49792 3470 49844 3476
rect 49240 3052 49292 3058
rect 49240 2994 49292 3000
rect 49792 3052 49844 3058
rect 49792 2994 49844 3000
rect 49608 2576 49660 2582
rect 49608 2518 49660 2524
rect 48320 2440 48372 2446
rect 48320 2382 48372 2388
rect 49620 800 49648 2518
rect 49804 2514 49832 2994
rect 49792 2508 49844 2514
rect 49792 2450 49844 2456
rect 49896 2446 49924 3878
rect 49988 2650 50016 4490
rect 50528 4480 50580 4486
rect 50528 4422 50580 4428
rect 50540 4146 50568 4422
rect 50528 4140 50580 4146
rect 50528 4082 50580 4088
rect 50068 4072 50120 4078
rect 50068 4014 50120 4020
rect 50080 3194 50108 4014
rect 51092 3942 51120 4655
rect 67234 4380 67542 4389
rect 67234 4378 67240 4380
rect 67296 4378 67320 4380
rect 67376 4378 67400 4380
rect 67456 4378 67480 4380
rect 67536 4378 67542 4380
rect 67296 4326 67298 4378
rect 67478 4326 67480 4378
rect 67234 4324 67240 4326
rect 67296 4324 67320 4326
rect 67376 4324 67400 4326
rect 67456 4324 67480 4326
rect 67536 4324 67542 4326
rect 67234 4315 67542 4324
rect 52644 4208 52696 4214
rect 52642 4176 52644 4185
rect 52696 4176 52698 4185
rect 52642 4111 52698 4120
rect 74632 4140 74684 4146
rect 74632 4082 74684 4088
rect 65432 4072 65484 4078
rect 65432 4014 65484 4020
rect 67916 4072 67968 4078
rect 67916 4014 67968 4020
rect 71688 4072 71740 4078
rect 71688 4014 71740 4020
rect 74080 4072 74132 4078
rect 74080 4014 74132 4020
rect 51080 3936 51132 3942
rect 51080 3878 51132 3884
rect 52368 3936 52420 3942
rect 52368 3878 52420 3884
rect 50620 3392 50672 3398
rect 50620 3334 50672 3340
rect 50068 3188 50120 3194
rect 50068 3130 50120 3136
rect 50632 3058 50660 3334
rect 51092 3058 51120 3878
rect 51264 3528 51316 3534
rect 51264 3470 51316 3476
rect 51276 3194 51304 3470
rect 51448 3392 51500 3398
rect 51448 3334 51500 3340
rect 51264 3188 51316 3194
rect 51264 3130 51316 3136
rect 51460 3058 51488 3334
rect 52380 3058 52408 3878
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 53656 3528 53708 3534
rect 53656 3470 53708 3476
rect 57336 3528 57388 3534
rect 57336 3470 57388 3476
rect 58072 3528 58124 3534
rect 58072 3470 58124 3476
rect 60924 3528 60976 3534
rect 60924 3470 60976 3476
rect 62120 3528 62172 3534
rect 62120 3470 62172 3476
rect 64696 3528 64748 3534
rect 64696 3470 64748 3476
rect 52472 3194 52500 3470
rect 53012 3392 53064 3398
rect 53012 3334 53064 3340
rect 52460 3188 52512 3194
rect 52460 3130 52512 3136
rect 50620 3052 50672 3058
rect 50620 2994 50672 3000
rect 51080 3052 51132 3058
rect 51080 2994 51132 3000
rect 51448 3052 51500 3058
rect 51448 2994 51500 3000
rect 52092 3052 52144 3058
rect 52092 2994 52144 3000
rect 52368 3052 52420 3058
rect 52368 2994 52420 3000
rect 51540 2984 51592 2990
rect 51540 2926 51592 2932
rect 49976 2644 50028 2650
rect 49976 2586 50028 2592
rect 49884 2440 49936 2446
rect 49884 2382 49936 2388
rect 50528 2440 50580 2446
rect 50528 2382 50580 2388
rect 50540 2038 50568 2382
rect 50528 2032 50580 2038
rect 50528 1974 50580 1980
rect 51552 800 51580 2926
rect 52104 2514 52132 2994
rect 52092 2508 52144 2514
rect 52092 2450 52144 2456
rect 53024 2446 53052 3334
rect 53668 3194 53696 3470
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 53656 3188 53708 3194
rect 53656 3130 53708 3136
rect 56060 3058 56088 3334
rect 57348 3194 57376 3470
rect 57428 3392 57480 3398
rect 57428 3334 57480 3340
rect 57336 3188 57388 3194
rect 57336 3130 57388 3136
rect 57440 3058 57468 3334
rect 58084 3194 58112 3470
rect 58624 3392 58676 3398
rect 58624 3334 58676 3340
rect 58072 3188 58124 3194
rect 58072 3130 58124 3136
rect 54024 3052 54076 3058
rect 54024 2994 54076 3000
rect 56048 3052 56100 3058
rect 56048 2994 56100 3000
rect 57428 3052 57480 3058
rect 57428 2994 57480 3000
rect 53472 2984 53524 2990
rect 53472 2926 53524 2932
rect 53012 2440 53064 2446
rect 53012 2382 53064 2388
rect 53484 800 53512 2926
rect 54036 2514 54064 2994
rect 55312 2848 55364 2854
rect 55312 2790 55364 2796
rect 54024 2508 54076 2514
rect 54024 2450 54076 2456
rect 55324 2446 55352 2790
rect 58636 2446 58664 3334
rect 60936 3194 60964 3470
rect 61108 3392 61160 3398
rect 61108 3334 61160 3340
rect 60924 3188 60976 3194
rect 60924 3130 60976 3136
rect 61120 3058 61148 3334
rect 62132 3194 62160 3470
rect 62764 3392 62816 3398
rect 62764 3334 62816 3340
rect 62120 3188 62172 3194
rect 62120 3130 62172 3136
rect 61108 3052 61160 3058
rect 61108 2994 61160 3000
rect 61752 3052 61804 3058
rect 61752 2994 61804 3000
rect 61200 2984 61252 2990
rect 61200 2926 61252 2932
rect 59268 2848 59320 2854
rect 59268 2790 59320 2796
rect 55312 2440 55364 2446
rect 55312 2382 55364 2388
rect 55404 2440 55456 2446
rect 55404 2382 55456 2388
rect 58624 2440 58676 2446
rect 58624 2382 58676 2388
rect 55416 800 55444 2382
rect 57336 2372 57388 2378
rect 57336 2314 57388 2320
rect 57348 800 57376 2314
rect 59280 800 59308 2790
rect 61212 800 61240 2926
rect 61764 2514 61792 2994
rect 61752 2508 61804 2514
rect 61752 2450 61804 2456
rect 62776 2446 62804 3334
rect 64708 3194 64736 3470
rect 64880 3392 64932 3398
rect 64880 3334 64932 3340
rect 64696 3188 64748 3194
rect 64696 3130 64748 3136
rect 64892 3058 64920 3334
rect 65444 3194 65472 4014
rect 66260 3936 66312 3942
rect 66260 3878 66312 3884
rect 65432 3188 65484 3194
rect 65432 3130 65484 3136
rect 64880 3052 64932 3058
rect 64880 2994 64932 3000
rect 65524 3052 65576 3058
rect 65524 2994 65576 3000
rect 65064 2984 65116 2990
rect 65064 2926 65116 2932
rect 62764 2440 62816 2446
rect 62764 2382 62816 2388
rect 63132 2440 63184 2446
rect 63132 2382 63184 2388
rect 63144 800 63172 2382
rect 65076 800 65104 2926
rect 65536 2514 65564 2994
rect 65524 2508 65576 2514
rect 65524 2450 65576 2456
rect 66272 2446 66300 3878
rect 66574 3836 66882 3845
rect 66574 3834 66580 3836
rect 66636 3834 66660 3836
rect 66716 3834 66740 3836
rect 66796 3834 66820 3836
rect 66876 3834 66882 3836
rect 66636 3782 66638 3834
rect 66818 3782 66820 3834
rect 66574 3780 66580 3782
rect 66636 3780 66660 3782
rect 66716 3780 66740 3782
rect 66796 3780 66820 3782
rect 66876 3780 66882 3782
rect 66574 3771 66882 3780
rect 67928 3738 67956 4014
rect 68284 3936 68336 3942
rect 68284 3878 68336 3884
rect 67916 3732 67968 3738
rect 67916 3674 67968 3680
rect 67088 3528 67140 3534
rect 67088 3470 67140 3476
rect 67100 3194 67128 3470
rect 67234 3292 67542 3301
rect 67234 3290 67240 3292
rect 67296 3290 67320 3292
rect 67376 3290 67400 3292
rect 67456 3290 67480 3292
rect 67536 3290 67542 3292
rect 67296 3238 67298 3290
rect 67478 3238 67480 3290
rect 67234 3236 67240 3238
rect 67296 3236 67320 3238
rect 67376 3236 67400 3238
rect 67456 3236 67480 3238
rect 67536 3236 67542 3238
rect 67234 3227 67542 3236
rect 67088 3188 67140 3194
rect 67088 3130 67140 3136
rect 67640 3052 67692 3058
rect 67640 2994 67692 3000
rect 66996 2916 67048 2922
rect 66996 2858 67048 2864
rect 66574 2748 66882 2757
rect 66574 2746 66580 2748
rect 66636 2746 66660 2748
rect 66716 2746 66740 2748
rect 66796 2746 66820 2748
rect 66876 2746 66882 2748
rect 66636 2694 66638 2746
rect 66818 2694 66820 2746
rect 66574 2692 66580 2694
rect 66636 2692 66660 2694
rect 66716 2692 66740 2694
rect 66796 2692 66820 2694
rect 66876 2692 66882 2694
rect 66574 2683 66882 2692
rect 66260 2440 66312 2446
rect 66260 2382 66312 2388
rect 67008 800 67036 2858
rect 67652 2514 67680 2994
rect 67640 2508 67692 2514
rect 67640 2450 67692 2456
rect 68296 2446 68324 3878
rect 71700 3738 71728 4014
rect 72424 3936 72476 3942
rect 72424 3878 72476 3884
rect 71688 3732 71740 3738
rect 71688 3674 71740 3680
rect 72436 3602 72464 3878
rect 74092 3777 74120 4014
rect 74078 3768 74134 3777
rect 74078 3703 74134 3712
rect 72424 3596 72476 3602
rect 72424 3538 72476 3544
rect 69112 3528 69164 3534
rect 69112 3470 69164 3476
rect 72240 3528 72292 3534
rect 72240 3470 72292 3476
rect 69124 3194 69152 3470
rect 71504 3392 71556 3398
rect 71504 3334 71556 3340
rect 69112 3188 69164 3194
rect 69112 3130 69164 3136
rect 70308 3120 70360 3126
rect 70308 3062 70360 3068
rect 69480 3052 69532 3058
rect 69480 2994 69532 3000
rect 68928 2984 68980 2990
rect 68928 2926 68980 2932
rect 68284 2440 68336 2446
rect 68284 2382 68336 2388
rect 67234 2204 67542 2213
rect 67234 2202 67240 2204
rect 67296 2202 67320 2204
rect 67376 2202 67400 2204
rect 67456 2202 67480 2204
rect 67536 2202 67542 2204
rect 67296 2150 67298 2202
rect 67478 2150 67480 2202
rect 67234 2148 67240 2150
rect 67296 2148 67320 2150
rect 67376 2148 67400 2150
rect 67456 2148 67480 2150
rect 67536 2148 67542 2150
rect 67234 2139 67542 2148
rect 68940 800 68968 2926
rect 69492 2514 69520 2994
rect 70320 2514 70348 3062
rect 71516 3058 71544 3334
rect 71504 3052 71556 3058
rect 71504 2994 71556 3000
rect 70860 2984 70912 2990
rect 70860 2926 70912 2932
rect 70492 2848 70544 2854
rect 70492 2790 70544 2796
rect 69480 2508 69532 2514
rect 69480 2450 69532 2456
rect 70308 2508 70360 2514
rect 70308 2450 70360 2456
rect 70504 2446 70532 2790
rect 70492 2440 70544 2446
rect 70492 2382 70544 2388
rect 70872 800 70900 2926
rect 72252 2650 72280 3470
rect 73068 3392 73120 3398
rect 73068 3334 73120 3340
rect 72608 3052 72660 3058
rect 72608 2994 72660 3000
rect 72240 2644 72292 2650
rect 72240 2586 72292 2592
rect 72620 2514 72648 2994
rect 72608 2508 72660 2514
rect 72608 2450 72660 2456
rect 72792 2508 72844 2514
rect 72792 2450 72844 2456
rect 72804 800 72832 2450
rect 73080 2446 73108 3334
rect 74092 3058 74120 3703
rect 74448 3528 74500 3534
rect 74448 3470 74500 3476
rect 74460 3194 74488 3470
rect 74540 3392 74592 3398
rect 74540 3334 74592 3340
rect 74448 3188 74500 3194
rect 74448 3130 74500 3136
rect 74552 3058 74580 3334
rect 74080 3052 74132 3058
rect 74080 2994 74132 3000
rect 74540 3052 74592 3058
rect 74540 2994 74592 3000
rect 74644 2650 74672 4082
rect 76564 4072 76616 4078
rect 76564 4014 76616 4020
rect 75460 3460 75512 3466
rect 75460 3402 75512 3408
rect 74724 2984 74776 2990
rect 74724 2926 74776 2932
rect 74632 2644 74684 2650
rect 74632 2586 74684 2592
rect 73068 2440 73120 2446
rect 73068 2382 73120 2388
rect 74736 800 74764 2926
rect 75472 2514 75500 3402
rect 76196 2848 76248 2854
rect 76196 2790 76248 2796
rect 75460 2508 75512 2514
rect 75460 2450 75512 2456
rect 76208 2446 76236 2790
rect 76196 2440 76248 2446
rect 76196 2382 76248 2388
rect 76576 2122 76604 4014
rect 76668 3534 76696 4966
rect 76944 4826 76972 5102
rect 76932 4820 76984 4826
rect 76932 4762 76984 4768
rect 77576 4616 77628 4622
rect 77576 4558 77628 4564
rect 77024 4072 77076 4078
rect 77024 4014 77076 4020
rect 77036 3602 77064 4014
rect 77588 3738 77616 4558
rect 77576 3732 77628 3738
rect 77576 3674 77628 3680
rect 77024 3596 77076 3602
rect 77024 3538 77076 3544
rect 76656 3528 76708 3534
rect 76656 3470 76708 3476
rect 76656 3052 76708 3058
rect 76656 2994 76708 3000
rect 76668 2650 76696 2994
rect 76656 2644 76708 2650
rect 76656 2586 76708 2592
rect 76576 2094 76696 2122
rect 76668 800 76696 2094
rect 46492 734 46704 762
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 77298 0 77354 800
<< via2 >>
rect 5140 37562 5196 37564
rect 5220 37562 5276 37564
rect 5300 37562 5356 37564
rect 5380 37562 5436 37564
rect 5140 37510 5186 37562
rect 5186 37510 5196 37562
rect 5220 37510 5250 37562
rect 5250 37510 5262 37562
rect 5262 37510 5276 37562
rect 5300 37510 5314 37562
rect 5314 37510 5326 37562
rect 5326 37510 5356 37562
rect 5380 37510 5390 37562
rect 5390 37510 5436 37562
rect 5140 37508 5196 37510
rect 5220 37508 5276 37510
rect 5300 37508 5356 37510
rect 5380 37508 5436 37510
rect 5800 37018 5856 37020
rect 5880 37018 5936 37020
rect 5960 37018 6016 37020
rect 6040 37018 6096 37020
rect 5800 36966 5846 37018
rect 5846 36966 5856 37018
rect 5880 36966 5910 37018
rect 5910 36966 5922 37018
rect 5922 36966 5936 37018
rect 5960 36966 5974 37018
rect 5974 36966 5986 37018
rect 5986 36966 6016 37018
rect 6040 36966 6050 37018
rect 6050 36966 6096 37018
rect 5800 36964 5856 36966
rect 5880 36964 5936 36966
rect 5960 36964 6016 36966
rect 6040 36964 6096 36966
rect 7010 36488 7066 36544
rect 5140 36474 5196 36476
rect 5220 36474 5276 36476
rect 5300 36474 5356 36476
rect 5380 36474 5436 36476
rect 5140 36422 5186 36474
rect 5186 36422 5196 36474
rect 5220 36422 5250 36474
rect 5250 36422 5262 36474
rect 5262 36422 5276 36474
rect 5300 36422 5314 36474
rect 5314 36422 5326 36474
rect 5326 36422 5356 36474
rect 5380 36422 5390 36474
rect 5390 36422 5436 36474
rect 5140 36420 5196 36422
rect 5220 36420 5276 36422
rect 5300 36420 5356 36422
rect 5380 36420 5436 36422
rect 5800 35930 5856 35932
rect 5880 35930 5936 35932
rect 5960 35930 6016 35932
rect 6040 35930 6096 35932
rect 5800 35878 5846 35930
rect 5846 35878 5856 35930
rect 5880 35878 5910 35930
rect 5910 35878 5922 35930
rect 5922 35878 5936 35930
rect 5960 35878 5974 35930
rect 5974 35878 5986 35930
rect 5986 35878 6016 35930
rect 6040 35878 6050 35930
rect 6050 35878 6096 35930
rect 5800 35876 5856 35878
rect 5880 35876 5936 35878
rect 5960 35876 6016 35878
rect 6040 35876 6096 35878
rect 5140 35386 5196 35388
rect 5220 35386 5276 35388
rect 5300 35386 5356 35388
rect 5380 35386 5436 35388
rect 5140 35334 5186 35386
rect 5186 35334 5196 35386
rect 5220 35334 5250 35386
rect 5250 35334 5262 35386
rect 5262 35334 5276 35386
rect 5300 35334 5314 35386
rect 5314 35334 5326 35386
rect 5326 35334 5356 35386
rect 5380 35334 5390 35386
rect 5390 35334 5436 35386
rect 5140 35332 5196 35334
rect 5220 35332 5276 35334
rect 5300 35332 5356 35334
rect 5380 35332 5436 35334
rect 5800 34842 5856 34844
rect 5880 34842 5936 34844
rect 5960 34842 6016 34844
rect 6040 34842 6096 34844
rect 5800 34790 5846 34842
rect 5846 34790 5856 34842
rect 5880 34790 5910 34842
rect 5910 34790 5922 34842
rect 5922 34790 5936 34842
rect 5960 34790 5974 34842
rect 5974 34790 5986 34842
rect 5986 34790 6016 34842
rect 6040 34790 6050 34842
rect 6050 34790 6096 34842
rect 5800 34788 5856 34790
rect 5880 34788 5936 34790
rect 5960 34788 6016 34790
rect 6040 34788 6096 34790
rect 5140 34298 5196 34300
rect 5220 34298 5276 34300
rect 5300 34298 5356 34300
rect 5380 34298 5436 34300
rect 5140 34246 5186 34298
rect 5186 34246 5196 34298
rect 5220 34246 5250 34298
rect 5250 34246 5262 34298
rect 5262 34246 5276 34298
rect 5300 34246 5314 34298
rect 5314 34246 5326 34298
rect 5326 34246 5356 34298
rect 5380 34246 5390 34298
rect 5390 34246 5436 34298
rect 5140 34244 5196 34246
rect 5220 34244 5276 34246
rect 5300 34244 5356 34246
rect 5380 34244 5436 34246
rect 5800 33754 5856 33756
rect 5880 33754 5936 33756
rect 5960 33754 6016 33756
rect 6040 33754 6096 33756
rect 5800 33702 5846 33754
rect 5846 33702 5856 33754
rect 5880 33702 5910 33754
rect 5910 33702 5922 33754
rect 5922 33702 5936 33754
rect 5960 33702 5974 33754
rect 5974 33702 5986 33754
rect 5986 33702 6016 33754
rect 6040 33702 6050 33754
rect 6050 33702 6096 33754
rect 5800 33700 5856 33702
rect 5880 33700 5936 33702
rect 5960 33700 6016 33702
rect 6040 33700 6096 33702
rect 5140 33210 5196 33212
rect 5220 33210 5276 33212
rect 5300 33210 5356 33212
rect 5380 33210 5436 33212
rect 5140 33158 5186 33210
rect 5186 33158 5196 33210
rect 5220 33158 5250 33210
rect 5250 33158 5262 33210
rect 5262 33158 5276 33210
rect 5300 33158 5314 33210
rect 5314 33158 5326 33210
rect 5326 33158 5356 33210
rect 5380 33158 5390 33210
rect 5390 33158 5436 33210
rect 5140 33156 5196 33158
rect 5220 33156 5276 33158
rect 5300 33156 5356 33158
rect 5380 33156 5436 33158
rect 5800 32666 5856 32668
rect 5880 32666 5936 32668
rect 5960 32666 6016 32668
rect 6040 32666 6096 32668
rect 5800 32614 5846 32666
rect 5846 32614 5856 32666
rect 5880 32614 5910 32666
rect 5910 32614 5922 32666
rect 5922 32614 5936 32666
rect 5960 32614 5974 32666
rect 5974 32614 5986 32666
rect 5986 32614 6016 32666
rect 6040 32614 6050 32666
rect 6050 32614 6096 32666
rect 5800 32612 5856 32614
rect 5880 32612 5936 32614
rect 5960 32612 6016 32614
rect 6040 32612 6096 32614
rect 5140 32122 5196 32124
rect 5220 32122 5276 32124
rect 5300 32122 5356 32124
rect 5380 32122 5436 32124
rect 5140 32070 5186 32122
rect 5186 32070 5196 32122
rect 5220 32070 5250 32122
rect 5250 32070 5262 32122
rect 5262 32070 5276 32122
rect 5300 32070 5314 32122
rect 5314 32070 5326 32122
rect 5326 32070 5356 32122
rect 5380 32070 5390 32122
rect 5390 32070 5436 32122
rect 5140 32068 5196 32070
rect 5220 32068 5276 32070
rect 5300 32068 5356 32070
rect 5380 32068 5436 32070
rect 5800 31578 5856 31580
rect 5880 31578 5936 31580
rect 5960 31578 6016 31580
rect 6040 31578 6096 31580
rect 5800 31526 5846 31578
rect 5846 31526 5856 31578
rect 5880 31526 5910 31578
rect 5910 31526 5922 31578
rect 5922 31526 5936 31578
rect 5960 31526 5974 31578
rect 5974 31526 5986 31578
rect 5986 31526 6016 31578
rect 6040 31526 6050 31578
rect 6050 31526 6096 31578
rect 5800 31524 5856 31526
rect 5880 31524 5936 31526
rect 5960 31524 6016 31526
rect 6040 31524 6096 31526
rect 5140 31034 5196 31036
rect 5220 31034 5276 31036
rect 5300 31034 5356 31036
rect 5380 31034 5436 31036
rect 5140 30982 5186 31034
rect 5186 30982 5196 31034
rect 5220 30982 5250 31034
rect 5250 30982 5262 31034
rect 5262 30982 5276 31034
rect 5300 30982 5314 31034
rect 5314 30982 5326 31034
rect 5326 30982 5356 31034
rect 5380 30982 5390 31034
rect 5390 30982 5436 31034
rect 5140 30980 5196 30982
rect 5220 30980 5276 30982
rect 5300 30980 5356 30982
rect 5380 30980 5436 30982
rect 5800 30490 5856 30492
rect 5880 30490 5936 30492
rect 5960 30490 6016 30492
rect 6040 30490 6096 30492
rect 5800 30438 5846 30490
rect 5846 30438 5856 30490
rect 5880 30438 5910 30490
rect 5910 30438 5922 30490
rect 5922 30438 5936 30490
rect 5960 30438 5974 30490
rect 5974 30438 5986 30490
rect 5986 30438 6016 30490
rect 6040 30438 6050 30490
rect 6050 30438 6096 30490
rect 5800 30436 5856 30438
rect 5880 30436 5936 30438
rect 5960 30436 6016 30438
rect 6040 30436 6096 30438
rect 5140 29946 5196 29948
rect 5220 29946 5276 29948
rect 5300 29946 5356 29948
rect 5380 29946 5436 29948
rect 5140 29894 5186 29946
rect 5186 29894 5196 29946
rect 5220 29894 5250 29946
rect 5250 29894 5262 29946
rect 5262 29894 5276 29946
rect 5300 29894 5314 29946
rect 5314 29894 5326 29946
rect 5326 29894 5356 29946
rect 5380 29894 5390 29946
rect 5390 29894 5436 29946
rect 5140 29892 5196 29894
rect 5220 29892 5276 29894
rect 5300 29892 5356 29894
rect 5380 29892 5436 29894
rect 5800 29402 5856 29404
rect 5880 29402 5936 29404
rect 5960 29402 6016 29404
rect 6040 29402 6096 29404
rect 5800 29350 5846 29402
rect 5846 29350 5856 29402
rect 5880 29350 5910 29402
rect 5910 29350 5922 29402
rect 5922 29350 5936 29402
rect 5960 29350 5974 29402
rect 5974 29350 5986 29402
rect 5986 29350 6016 29402
rect 6040 29350 6050 29402
rect 6050 29350 6096 29402
rect 5800 29348 5856 29350
rect 5880 29348 5936 29350
rect 5960 29348 6016 29350
rect 6040 29348 6096 29350
rect 5140 28858 5196 28860
rect 5220 28858 5276 28860
rect 5300 28858 5356 28860
rect 5380 28858 5436 28860
rect 5140 28806 5186 28858
rect 5186 28806 5196 28858
rect 5220 28806 5250 28858
rect 5250 28806 5262 28858
rect 5262 28806 5276 28858
rect 5300 28806 5314 28858
rect 5314 28806 5326 28858
rect 5326 28806 5356 28858
rect 5380 28806 5390 28858
rect 5390 28806 5436 28858
rect 5140 28804 5196 28806
rect 5220 28804 5276 28806
rect 5300 28804 5356 28806
rect 5380 28804 5436 28806
rect 5800 28314 5856 28316
rect 5880 28314 5936 28316
rect 5960 28314 6016 28316
rect 6040 28314 6096 28316
rect 5800 28262 5846 28314
rect 5846 28262 5856 28314
rect 5880 28262 5910 28314
rect 5910 28262 5922 28314
rect 5922 28262 5936 28314
rect 5960 28262 5974 28314
rect 5974 28262 5986 28314
rect 5986 28262 6016 28314
rect 6040 28262 6050 28314
rect 6050 28262 6096 28314
rect 5800 28260 5856 28262
rect 5880 28260 5936 28262
rect 5960 28260 6016 28262
rect 6040 28260 6096 28262
rect 5140 27770 5196 27772
rect 5220 27770 5276 27772
rect 5300 27770 5356 27772
rect 5380 27770 5436 27772
rect 5140 27718 5186 27770
rect 5186 27718 5196 27770
rect 5220 27718 5250 27770
rect 5250 27718 5262 27770
rect 5262 27718 5276 27770
rect 5300 27718 5314 27770
rect 5314 27718 5326 27770
rect 5326 27718 5356 27770
rect 5380 27718 5390 27770
rect 5390 27718 5436 27770
rect 5140 27716 5196 27718
rect 5220 27716 5276 27718
rect 5300 27716 5356 27718
rect 5380 27716 5436 27718
rect 5800 27226 5856 27228
rect 5880 27226 5936 27228
rect 5960 27226 6016 27228
rect 6040 27226 6096 27228
rect 5800 27174 5846 27226
rect 5846 27174 5856 27226
rect 5880 27174 5910 27226
rect 5910 27174 5922 27226
rect 5922 27174 5936 27226
rect 5960 27174 5974 27226
rect 5974 27174 5986 27226
rect 5986 27174 6016 27226
rect 6040 27174 6050 27226
rect 6050 27174 6096 27226
rect 5800 27172 5856 27174
rect 5880 27172 5936 27174
rect 5960 27172 6016 27174
rect 6040 27172 6096 27174
rect 10874 26832 10930 26888
rect 5140 26682 5196 26684
rect 5220 26682 5276 26684
rect 5300 26682 5356 26684
rect 5380 26682 5436 26684
rect 5140 26630 5186 26682
rect 5186 26630 5196 26682
rect 5220 26630 5250 26682
rect 5250 26630 5262 26682
rect 5262 26630 5276 26682
rect 5300 26630 5314 26682
rect 5314 26630 5326 26682
rect 5326 26630 5356 26682
rect 5380 26630 5390 26682
rect 5390 26630 5436 26682
rect 5140 26628 5196 26630
rect 5220 26628 5276 26630
rect 5300 26628 5356 26630
rect 5380 26628 5436 26630
rect 5800 26138 5856 26140
rect 5880 26138 5936 26140
rect 5960 26138 6016 26140
rect 6040 26138 6096 26140
rect 5800 26086 5846 26138
rect 5846 26086 5856 26138
rect 5880 26086 5910 26138
rect 5910 26086 5922 26138
rect 5922 26086 5936 26138
rect 5960 26086 5974 26138
rect 5974 26086 5986 26138
rect 5986 26086 6016 26138
rect 6040 26086 6050 26138
rect 6050 26086 6096 26138
rect 5800 26084 5856 26086
rect 5880 26084 5936 26086
rect 5960 26084 6016 26086
rect 6040 26084 6096 26086
rect 5140 25594 5196 25596
rect 5220 25594 5276 25596
rect 5300 25594 5356 25596
rect 5380 25594 5436 25596
rect 5140 25542 5186 25594
rect 5186 25542 5196 25594
rect 5220 25542 5250 25594
rect 5250 25542 5262 25594
rect 5262 25542 5276 25594
rect 5300 25542 5314 25594
rect 5314 25542 5326 25594
rect 5326 25542 5356 25594
rect 5380 25542 5390 25594
rect 5390 25542 5436 25594
rect 5140 25540 5196 25542
rect 5220 25540 5276 25542
rect 5300 25540 5356 25542
rect 5380 25540 5436 25542
rect 5800 25050 5856 25052
rect 5880 25050 5936 25052
rect 5960 25050 6016 25052
rect 6040 25050 6096 25052
rect 5800 24998 5846 25050
rect 5846 24998 5856 25050
rect 5880 24998 5910 25050
rect 5910 24998 5922 25050
rect 5922 24998 5936 25050
rect 5960 24998 5974 25050
rect 5974 24998 5986 25050
rect 5986 24998 6016 25050
rect 6040 24998 6050 25050
rect 6050 24998 6096 25050
rect 5800 24996 5856 24998
rect 5880 24996 5936 24998
rect 5960 24996 6016 24998
rect 6040 24996 6096 24998
rect 5140 24506 5196 24508
rect 5220 24506 5276 24508
rect 5300 24506 5356 24508
rect 5380 24506 5436 24508
rect 5140 24454 5186 24506
rect 5186 24454 5196 24506
rect 5220 24454 5250 24506
rect 5250 24454 5262 24506
rect 5262 24454 5276 24506
rect 5300 24454 5314 24506
rect 5314 24454 5326 24506
rect 5326 24454 5356 24506
rect 5380 24454 5390 24506
rect 5390 24454 5436 24506
rect 5140 24452 5196 24454
rect 5220 24452 5276 24454
rect 5300 24452 5356 24454
rect 5380 24452 5436 24454
rect 3514 24112 3570 24168
rect 5800 23962 5856 23964
rect 5880 23962 5936 23964
rect 5960 23962 6016 23964
rect 6040 23962 6096 23964
rect 5800 23910 5846 23962
rect 5846 23910 5856 23962
rect 5880 23910 5910 23962
rect 5910 23910 5922 23962
rect 5922 23910 5936 23962
rect 5960 23910 5974 23962
rect 5974 23910 5986 23962
rect 5986 23910 6016 23962
rect 6040 23910 6050 23962
rect 6050 23910 6096 23962
rect 5800 23908 5856 23910
rect 5880 23908 5936 23910
rect 5960 23908 6016 23910
rect 6040 23908 6096 23910
rect 5140 23418 5196 23420
rect 5220 23418 5276 23420
rect 5300 23418 5356 23420
rect 5380 23418 5436 23420
rect 5140 23366 5186 23418
rect 5186 23366 5196 23418
rect 5220 23366 5250 23418
rect 5250 23366 5262 23418
rect 5262 23366 5276 23418
rect 5300 23366 5314 23418
rect 5314 23366 5326 23418
rect 5326 23366 5356 23418
rect 5380 23366 5390 23418
rect 5390 23366 5436 23418
rect 5140 23364 5196 23366
rect 5220 23364 5276 23366
rect 5300 23364 5356 23366
rect 5380 23364 5436 23366
rect 5800 22874 5856 22876
rect 5880 22874 5936 22876
rect 5960 22874 6016 22876
rect 6040 22874 6096 22876
rect 5800 22822 5846 22874
rect 5846 22822 5856 22874
rect 5880 22822 5910 22874
rect 5910 22822 5922 22874
rect 5922 22822 5936 22874
rect 5960 22822 5974 22874
rect 5974 22822 5986 22874
rect 5986 22822 6016 22874
rect 6040 22822 6050 22874
rect 6050 22822 6096 22874
rect 5800 22820 5856 22822
rect 5880 22820 5936 22822
rect 5960 22820 6016 22822
rect 6040 22820 6096 22822
rect 5140 22330 5196 22332
rect 5220 22330 5276 22332
rect 5300 22330 5356 22332
rect 5380 22330 5436 22332
rect 5140 22278 5186 22330
rect 5186 22278 5196 22330
rect 5220 22278 5250 22330
rect 5250 22278 5262 22330
rect 5262 22278 5276 22330
rect 5300 22278 5314 22330
rect 5314 22278 5326 22330
rect 5326 22278 5356 22330
rect 5380 22278 5390 22330
rect 5390 22278 5436 22330
rect 5140 22276 5196 22278
rect 5220 22276 5276 22278
rect 5300 22276 5356 22278
rect 5380 22276 5436 22278
rect 5800 21786 5856 21788
rect 5880 21786 5936 21788
rect 5960 21786 6016 21788
rect 6040 21786 6096 21788
rect 5800 21734 5846 21786
rect 5846 21734 5856 21786
rect 5880 21734 5910 21786
rect 5910 21734 5922 21786
rect 5922 21734 5936 21786
rect 5960 21734 5974 21786
rect 5974 21734 5986 21786
rect 5986 21734 6016 21786
rect 6040 21734 6050 21786
rect 6050 21734 6096 21786
rect 5800 21732 5856 21734
rect 5880 21732 5936 21734
rect 5960 21732 6016 21734
rect 6040 21732 6096 21734
rect 5140 21242 5196 21244
rect 5220 21242 5276 21244
rect 5300 21242 5356 21244
rect 5380 21242 5436 21244
rect 5140 21190 5186 21242
rect 5186 21190 5196 21242
rect 5220 21190 5250 21242
rect 5250 21190 5262 21242
rect 5262 21190 5276 21242
rect 5300 21190 5314 21242
rect 5314 21190 5326 21242
rect 5326 21190 5356 21242
rect 5380 21190 5390 21242
rect 5390 21190 5436 21242
rect 5140 21188 5196 21190
rect 5220 21188 5276 21190
rect 5300 21188 5356 21190
rect 5380 21188 5436 21190
rect 5800 20698 5856 20700
rect 5880 20698 5936 20700
rect 5960 20698 6016 20700
rect 6040 20698 6096 20700
rect 5800 20646 5846 20698
rect 5846 20646 5856 20698
rect 5880 20646 5910 20698
rect 5910 20646 5922 20698
rect 5922 20646 5936 20698
rect 5960 20646 5974 20698
rect 5974 20646 5986 20698
rect 5986 20646 6016 20698
rect 6040 20646 6050 20698
rect 6050 20646 6096 20698
rect 5800 20644 5856 20646
rect 5880 20644 5936 20646
rect 5960 20644 6016 20646
rect 6040 20644 6096 20646
rect 5140 20154 5196 20156
rect 5220 20154 5276 20156
rect 5300 20154 5356 20156
rect 5380 20154 5436 20156
rect 5140 20102 5186 20154
rect 5186 20102 5196 20154
rect 5220 20102 5250 20154
rect 5250 20102 5262 20154
rect 5262 20102 5276 20154
rect 5300 20102 5314 20154
rect 5314 20102 5326 20154
rect 5326 20102 5356 20154
rect 5380 20102 5390 20154
rect 5390 20102 5436 20154
rect 5140 20100 5196 20102
rect 5220 20100 5276 20102
rect 5300 20100 5356 20102
rect 5380 20100 5436 20102
rect 5800 19610 5856 19612
rect 5880 19610 5936 19612
rect 5960 19610 6016 19612
rect 6040 19610 6096 19612
rect 5800 19558 5846 19610
rect 5846 19558 5856 19610
rect 5880 19558 5910 19610
rect 5910 19558 5922 19610
rect 5922 19558 5936 19610
rect 5960 19558 5974 19610
rect 5974 19558 5986 19610
rect 5986 19558 6016 19610
rect 6040 19558 6050 19610
rect 6050 19558 6096 19610
rect 5800 19556 5856 19558
rect 5880 19556 5936 19558
rect 5960 19556 6016 19558
rect 6040 19556 6096 19558
rect 5140 19066 5196 19068
rect 5220 19066 5276 19068
rect 5300 19066 5356 19068
rect 5380 19066 5436 19068
rect 5140 19014 5186 19066
rect 5186 19014 5196 19066
rect 5220 19014 5250 19066
rect 5250 19014 5262 19066
rect 5262 19014 5276 19066
rect 5300 19014 5314 19066
rect 5314 19014 5326 19066
rect 5326 19014 5356 19066
rect 5380 19014 5390 19066
rect 5390 19014 5436 19066
rect 5140 19012 5196 19014
rect 5220 19012 5276 19014
rect 5300 19012 5356 19014
rect 5380 19012 5436 19014
rect 5800 18522 5856 18524
rect 5880 18522 5936 18524
rect 5960 18522 6016 18524
rect 6040 18522 6096 18524
rect 5800 18470 5846 18522
rect 5846 18470 5856 18522
rect 5880 18470 5910 18522
rect 5910 18470 5922 18522
rect 5922 18470 5936 18522
rect 5960 18470 5974 18522
rect 5974 18470 5986 18522
rect 5986 18470 6016 18522
rect 6040 18470 6050 18522
rect 6050 18470 6096 18522
rect 5800 18468 5856 18470
rect 5880 18468 5936 18470
rect 5960 18468 6016 18470
rect 6040 18468 6096 18470
rect 5140 17978 5196 17980
rect 5220 17978 5276 17980
rect 5300 17978 5356 17980
rect 5380 17978 5436 17980
rect 5140 17926 5186 17978
rect 5186 17926 5196 17978
rect 5220 17926 5250 17978
rect 5250 17926 5262 17978
rect 5262 17926 5276 17978
rect 5300 17926 5314 17978
rect 5314 17926 5326 17978
rect 5326 17926 5356 17978
rect 5380 17926 5390 17978
rect 5390 17926 5436 17978
rect 5140 17924 5196 17926
rect 5220 17924 5276 17926
rect 5300 17924 5356 17926
rect 5380 17924 5436 17926
rect 5800 17434 5856 17436
rect 5880 17434 5936 17436
rect 5960 17434 6016 17436
rect 6040 17434 6096 17436
rect 5800 17382 5846 17434
rect 5846 17382 5856 17434
rect 5880 17382 5910 17434
rect 5910 17382 5922 17434
rect 5922 17382 5936 17434
rect 5960 17382 5974 17434
rect 5974 17382 5986 17434
rect 5986 17382 6016 17434
rect 6040 17382 6050 17434
rect 6050 17382 6096 17434
rect 5800 17380 5856 17382
rect 5880 17380 5936 17382
rect 5960 17380 6016 17382
rect 6040 17380 6096 17382
rect 5140 16890 5196 16892
rect 5220 16890 5276 16892
rect 5300 16890 5356 16892
rect 5380 16890 5436 16892
rect 5140 16838 5186 16890
rect 5186 16838 5196 16890
rect 5220 16838 5250 16890
rect 5250 16838 5262 16890
rect 5262 16838 5276 16890
rect 5300 16838 5314 16890
rect 5314 16838 5326 16890
rect 5326 16838 5356 16890
rect 5380 16838 5390 16890
rect 5390 16838 5436 16890
rect 5140 16836 5196 16838
rect 5220 16836 5276 16838
rect 5300 16836 5356 16838
rect 5380 16836 5436 16838
rect 5800 16346 5856 16348
rect 5880 16346 5936 16348
rect 5960 16346 6016 16348
rect 6040 16346 6096 16348
rect 5800 16294 5846 16346
rect 5846 16294 5856 16346
rect 5880 16294 5910 16346
rect 5910 16294 5922 16346
rect 5922 16294 5936 16346
rect 5960 16294 5974 16346
rect 5974 16294 5986 16346
rect 5986 16294 6016 16346
rect 6040 16294 6050 16346
rect 6050 16294 6096 16346
rect 5800 16292 5856 16294
rect 5880 16292 5936 16294
rect 5960 16292 6016 16294
rect 6040 16292 6096 16294
rect 5140 15802 5196 15804
rect 5220 15802 5276 15804
rect 5300 15802 5356 15804
rect 5380 15802 5436 15804
rect 5140 15750 5186 15802
rect 5186 15750 5196 15802
rect 5220 15750 5250 15802
rect 5250 15750 5262 15802
rect 5262 15750 5276 15802
rect 5300 15750 5314 15802
rect 5314 15750 5326 15802
rect 5326 15750 5356 15802
rect 5380 15750 5390 15802
rect 5390 15750 5436 15802
rect 5140 15748 5196 15750
rect 5220 15748 5276 15750
rect 5300 15748 5356 15750
rect 5380 15748 5436 15750
rect 5800 15258 5856 15260
rect 5880 15258 5936 15260
rect 5960 15258 6016 15260
rect 6040 15258 6096 15260
rect 5800 15206 5846 15258
rect 5846 15206 5856 15258
rect 5880 15206 5910 15258
rect 5910 15206 5922 15258
rect 5922 15206 5936 15258
rect 5960 15206 5974 15258
rect 5974 15206 5986 15258
rect 5986 15206 6016 15258
rect 6040 15206 6050 15258
rect 6050 15206 6096 15258
rect 5800 15204 5856 15206
rect 5880 15204 5936 15206
rect 5960 15204 6016 15206
rect 6040 15204 6096 15206
rect 5140 14714 5196 14716
rect 5220 14714 5276 14716
rect 5300 14714 5356 14716
rect 5380 14714 5436 14716
rect 5140 14662 5186 14714
rect 5186 14662 5196 14714
rect 5220 14662 5250 14714
rect 5250 14662 5262 14714
rect 5262 14662 5276 14714
rect 5300 14662 5314 14714
rect 5314 14662 5326 14714
rect 5326 14662 5356 14714
rect 5380 14662 5390 14714
rect 5390 14662 5436 14714
rect 5140 14660 5196 14662
rect 5220 14660 5276 14662
rect 5300 14660 5356 14662
rect 5380 14660 5436 14662
rect 5800 14170 5856 14172
rect 5880 14170 5936 14172
rect 5960 14170 6016 14172
rect 6040 14170 6096 14172
rect 5800 14118 5846 14170
rect 5846 14118 5856 14170
rect 5880 14118 5910 14170
rect 5910 14118 5922 14170
rect 5922 14118 5936 14170
rect 5960 14118 5974 14170
rect 5974 14118 5986 14170
rect 5986 14118 6016 14170
rect 6040 14118 6050 14170
rect 6050 14118 6096 14170
rect 5800 14116 5856 14118
rect 5880 14116 5936 14118
rect 5960 14116 6016 14118
rect 6040 14116 6096 14118
rect 5140 13626 5196 13628
rect 5220 13626 5276 13628
rect 5300 13626 5356 13628
rect 5380 13626 5436 13628
rect 5140 13574 5186 13626
rect 5186 13574 5196 13626
rect 5220 13574 5250 13626
rect 5250 13574 5262 13626
rect 5262 13574 5276 13626
rect 5300 13574 5314 13626
rect 5314 13574 5326 13626
rect 5326 13574 5356 13626
rect 5380 13574 5390 13626
rect 5390 13574 5436 13626
rect 5140 13572 5196 13574
rect 5220 13572 5276 13574
rect 5300 13572 5356 13574
rect 5380 13572 5436 13574
rect 5800 13082 5856 13084
rect 5880 13082 5936 13084
rect 5960 13082 6016 13084
rect 6040 13082 6096 13084
rect 5800 13030 5846 13082
rect 5846 13030 5856 13082
rect 5880 13030 5910 13082
rect 5910 13030 5922 13082
rect 5922 13030 5936 13082
rect 5960 13030 5974 13082
rect 5974 13030 5986 13082
rect 5986 13030 6016 13082
rect 6040 13030 6050 13082
rect 6050 13030 6096 13082
rect 5800 13028 5856 13030
rect 5880 13028 5936 13030
rect 5960 13028 6016 13030
rect 6040 13028 6096 13030
rect 5140 12538 5196 12540
rect 5220 12538 5276 12540
rect 5300 12538 5356 12540
rect 5380 12538 5436 12540
rect 5140 12486 5186 12538
rect 5186 12486 5196 12538
rect 5220 12486 5250 12538
rect 5250 12486 5262 12538
rect 5262 12486 5276 12538
rect 5300 12486 5314 12538
rect 5314 12486 5326 12538
rect 5326 12486 5356 12538
rect 5380 12486 5390 12538
rect 5390 12486 5436 12538
rect 5140 12484 5196 12486
rect 5220 12484 5276 12486
rect 5300 12484 5356 12486
rect 5380 12484 5436 12486
rect 5800 11994 5856 11996
rect 5880 11994 5936 11996
rect 5960 11994 6016 11996
rect 6040 11994 6096 11996
rect 5800 11942 5846 11994
rect 5846 11942 5856 11994
rect 5880 11942 5910 11994
rect 5910 11942 5922 11994
rect 5922 11942 5936 11994
rect 5960 11942 5974 11994
rect 5974 11942 5986 11994
rect 5986 11942 6016 11994
rect 6040 11942 6050 11994
rect 6050 11942 6096 11994
rect 5800 11940 5856 11942
rect 5880 11940 5936 11942
rect 5960 11940 6016 11942
rect 6040 11940 6096 11942
rect 5140 11450 5196 11452
rect 5220 11450 5276 11452
rect 5300 11450 5356 11452
rect 5380 11450 5436 11452
rect 5140 11398 5186 11450
rect 5186 11398 5196 11450
rect 5220 11398 5250 11450
rect 5250 11398 5262 11450
rect 5262 11398 5276 11450
rect 5300 11398 5314 11450
rect 5314 11398 5326 11450
rect 5326 11398 5356 11450
rect 5380 11398 5390 11450
rect 5390 11398 5436 11450
rect 5140 11396 5196 11398
rect 5220 11396 5276 11398
rect 5300 11396 5356 11398
rect 5380 11396 5436 11398
rect 5800 10906 5856 10908
rect 5880 10906 5936 10908
rect 5960 10906 6016 10908
rect 6040 10906 6096 10908
rect 5800 10854 5846 10906
rect 5846 10854 5856 10906
rect 5880 10854 5910 10906
rect 5910 10854 5922 10906
rect 5922 10854 5936 10906
rect 5960 10854 5974 10906
rect 5974 10854 5986 10906
rect 5986 10854 6016 10906
rect 6040 10854 6050 10906
rect 6050 10854 6096 10906
rect 5800 10852 5856 10854
rect 5880 10852 5936 10854
rect 5960 10852 6016 10854
rect 6040 10852 6096 10854
rect 5140 10362 5196 10364
rect 5220 10362 5276 10364
rect 5300 10362 5356 10364
rect 5380 10362 5436 10364
rect 5140 10310 5186 10362
rect 5186 10310 5196 10362
rect 5220 10310 5250 10362
rect 5250 10310 5262 10362
rect 5262 10310 5276 10362
rect 5300 10310 5314 10362
rect 5314 10310 5326 10362
rect 5326 10310 5356 10362
rect 5380 10310 5390 10362
rect 5390 10310 5436 10362
rect 5140 10308 5196 10310
rect 5220 10308 5276 10310
rect 5300 10308 5356 10310
rect 5380 10308 5436 10310
rect 9034 9832 9090 9888
rect 5800 9818 5856 9820
rect 5880 9818 5936 9820
rect 5960 9818 6016 9820
rect 6040 9818 6096 9820
rect 5800 9766 5846 9818
rect 5846 9766 5856 9818
rect 5880 9766 5910 9818
rect 5910 9766 5922 9818
rect 5922 9766 5936 9818
rect 5960 9766 5974 9818
rect 5974 9766 5986 9818
rect 5986 9766 6016 9818
rect 6040 9766 6050 9818
rect 6050 9766 6096 9818
rect 5800 9764 5856 9766
rect 5880 9764 5936 9766
rect 5960 9764 6016 9766
rect 6040 9764 6096 9766
rect 5140 9274 5196 9276
rect 5220 9274 5276 9276
rect 5300 9274 5356 9276
rect 5380 9274 5436 9276
rect 5140 9222 5186 9274
rect 5186 9222 5196 9274
rect 5220 9222 5250 9274
rect 5250 9222 5262 9274
rect 5262 9222 5276 9274
rect 5300 9222 5314 9274
rect 5314 9222 5326 9274
rect 5326 9222 5356 9274
rect 5380 9222 5390 9274
rect 5390 9222 5436 9274
rect 5140 9220 5196 9222
rect 5220 9220 5276 9222
rect 5300 9220 5356 9222
rect 5380 9220 5436 9222
rect 5800 8730 5856 8732
rect 5880 8730 5936 8732
rect 5960 8730 6016 8732
rect 6040 8730 6096 8732
rect 5800 8678 5846 8730
rect 5846 8678 5856 8730
rect 5880 8678 5910 8730
rect 5910 8678 5922 8730
rect 5922 8678 5936 8730
rect 5960 8678 5974 8730
rect 5974 8678 5986 8730
rect 5986 8678 6016 8730
rect 6040 8678 6050 8730
rect 6050 8678 6096 8730
rect 5800 8676 5856 8678
rect 5880 8676 5936 8678
rect 5960 8676 6016 8678
rect 6040 8676 6096 8678
rect 5140 8186 5196 8188
rect 5220 8186 5276 8188
rect 5300 8186 5356 8188
rect 5380 8186 5436 8188
rect 5140 8134 5186 8186
rect 5186 8134 5196 8186
rect 5220 8134 5250 8186
rect 5250 8134 5262 8186
rect 5262 8134 5276 8186
rect 5300 8134 5314 8186
rect 5314 8134 5326 8186
rect 5326 8134 5356 8186
rect 5380 8134 5390 8186
rect 5390 8134 5436 8186
rect 5140 8132 5196 8134
rect 5220 8132 5276 8134
rect 5300 8132 5356 8134
rect 5380 8132 5436 8134
rect 5800 7642 5856 7644
rect 5880 7642 5936 7644
rect 5960 7642 6016 7644
rect 6040 7642 6096 7644
rect 5800 7590 5846 7642
rect 5846 7590 5856 7642
rect 5880 7590 5910 7642
rect 5910 7590 5922 7642
rect 5922 7590 5936 7642
rect 5960 7590 5974 7642
rect 5974 7590 5986 7642
rect 5986 7590 6016 7642
rect 6040 7590 6050 7642
rect 6050 7590 6096 7642
rect 5800 7588 5856 7590
rect 5880 7588 5936 7590
rect 5960 7588 6016 7590
rect 6040 7588 6096 7590
rect 5140 7098 5196 7100
rect 5220 7098 5276 7100
rect 5300 7098 5356 7100
rect 5380 7098 5436 7100
rect 5140 7046 5186 7098
rect 5186 7046 5196 7098
rect 5220 7046 5250 7098
rect 5250 7046 5262 7098
rect 5262 7046 5276 7098
rect 5300 7046 5314 7098
rect 5314 7046 5326 7098
rect 5326 7046 5356 7098
rect 5380 7046 5390 7098
rect 5390 7046 5436 7098
rect 5140 7044 5196 7046
rect 5220 7044 5276 7046
rect 5300 7044 5356 7046
rect 5380 7044 5436 7046
rect 5800 6554 5856 6556
rect 5880 6554 5936 6556
rect 5960 6554 6016 6556
rect 6040 6554 6096 6556
rect 5800 6502 5846 6554
rect 5846 6502 5856 6554
rect 5880 6502 5910 6554
rect 5910 6502 5922 6554
rect 5922 6502 5936 6554
rect 5960 6502 5974 6554
rect 5974 6502 5986 6554
rect 5986 6502 6016 6554
rect 6040 6502 6050 6554
rect 6050 6502 6096 6554
rect 5800 6500 5856 6502
rect 5880 6500 5936 6502
rect 5960 6500 6016 6502
rect 6040 6500 6096 6502
rect 5140 6010 5196 6012
rect 5220 6010 5276 6012
rect 5300 6010 5356 6012
rect 5380 6010 5436 6012
rect 5140 5958 5186 6010
rect 5186 5958 5196 6010
rect 5220 5958 5250 6010
rect 5250 5958 5262 6010
rect 5262 5958 5276 6010
rect 5300 5958 5314 6010
rect 5314 5958 5326 6010
rect 5326 5958 5356 6010
rect 5380 5958 5390 6010
rect 5390 5958 5436 6010
rect 5140 5956 5196 5958
rect 5220 5956 5276 5958
rect 5300 5956 5356 5958
rect 5380 5956 5436 5958
rect 5800 5466 5856 5468
rect 5880 5466 5936 5468
rect 5960 5466 6016 5468
rect 6040 5466 6096 5468
rect 5800 5414 5846 5466
rect 5846 5414 5856 5466
rect 5880 5414 5910 5466
rect 5910 5414 5922 5466
rect 5922 5414 5936 5466
rect 5960 5414 5974 5466
rect 5974 5414 5986 5466
rect 5986 5414 6016 5466
rect 6040 5414 6050 5466
rect 6050 5414 6096 5466
rect 5800 5412 5856 5414
rect 5880 5412 5936 5414
rect 5960 5412 6016 5414
rect 6040 5412 6096 5414
rect 5140 4922 5196 4924
rect 5220 4922 5276 4924
rect 5300 4922 5356 4924
rect 5380 4922 5436 4924
rect 5140 4870 5186 4922
rect 5186 4870 5196 4922
rect 5220 4870 5250 4922
rect 5250 4870 5262 4922
rect 5262 4870 5276 4922
rect 5300 4870 5314 4922
rect 5314 4870 5326 4922
rect 5326 4870 5356 4922
rect 5380 4870 5390 4922
rect 5390 4870 5436 4922
rect 5140 4868 5196 4870
rect 5220 4868 5276 4870
rect 5300 4868 5356 4870
rect 5380 4868 5436 4870
rect 5800 4378 5856 4380
rect 5880 4378 5936 4380
rect 5960 4378 6016 4380
rect 6040 4378 6096 4380
rect 5800 4326 5846 4378
rect 5846 4326 5856 4378
rect 5880 4326 5910 4378
rect 5910 4326 5922 4378
rect 5922 4326 5936 4378
rect 5960 4326 5974 4378
rect 5974 4326 5986 4378
rect 5986 4326 6016 4378
rect 6040 4326 6050 4378
rect 6050 4326 6096 4378
rect 5800 4324 5856 4326
rect 5880 4324 5936 4326
rect 5960 4324 6016 4326
rect 6040 4324 6096 4326
rect 5140 3834 5196 3836
rect 5220 3834 5276 3836
rect 5300 3834 5356 3836
rect 5380 3834 5436 3836
rect 5140 3782 5186 3834
rect 5186 3782 5196 3834
rect 5220 3782 5250 3834
rect 5250 3782 5262 3834
rect 5262 3782 5276 3834
rect 5300 3782 5314 3834
rect 5314 3782 5326 3834
rect 5326 3782 5356 3834
rect 5380 3782 5390 3834
rect 5390 3782 5436 3834
rect 5140 3780 5196 3782
rect 5220 3780 5276 3782
rect 5300 3780 5356 3782
rect 5380 3780 5436 3782
rect 5078 3576 5134 3632
rect 5140 2746 5196 2748
rect 5220 2746 5276 2748
rect 5300 2746 5356 2748
rect 5380 2746 5436 2748
rect 5140 2694 5186 2746
rect 5186 2694 5196 2746
rect 5220 2694 5250 2746
rect 5250 2694 5262 2746
rect 5262 2694 5276 2746
rect 5300 2694 5314 2746
rect 5314 2694 5326 2746
rect 5326 2694 5356 2746
rect 5380 2694 5390 2746
rect 5390 2694 5436 2746
rect 5140 2692 5196 2694
rect 5220 2692 5276 2694
rect 5300 2692 5356 2694
rect 5380 2692 5436 2694
rect 5630 2372 5686 2408
rect 5630 2352 5632 2372
rect 5632 2352 5684 2372
rect 5684 2352 5686 2372
rect 5800 3290 5856 3292
rect 5880 3290 5936 3292
rect 5960 3290 6016 3292
rect 6040 3290 6096 3292
rect 5800 3238 5846 3290
rect 5846 3238 5856 3290
rect 5880 3238 5910 3290
rect 5910 3238 5922 3290
rect 5922 3238 5936 3290
rect 5960 3238 5974 3290
rect 5974 3238 5986 3290
rect 5986 3238 6016 3290
rect 6040 3238 6050 3290
rect 6050 3238 6096 3290
rect 5800 3236 5856 3238
rect 5880 3236 5936 3238
rect 5960 3236 6016 3238
rect 6040 3236 6096 3238
rect 5814 2508 5870 2544
rect 5814 2488 5816 2508
rect 5816 2488 5868 2508
rect 5868 2488 5870 2508
rect 5800 2202 5856 2204
rect 5880 2202 5936 2204
rect 5960 2202 6016 2204
rect 6040 2202 6096 2204
rect 5800 2150 5846 2202
rect 5846 2150 5856 2202
rect 5880 2150 5910 2202
rect 5910 2150 5922 2202
rect 5922 2150 5936 2202
rect 5960 2150 5974 2202
rect 5974 2150 5986 2202
rect 5986 2150 6016 2202
rect 6040 2150 6050 2202
rect 6050 2150 6096 2202
rect 5800 2148 5856 2150
rect 5880 2148 5936 2150
rect 5960 2148 6016 2150
rect 6040 2148 6096 2150
rect 7470 3576 7526 3632
rect 7654 3168 7710 3224
rect 8390 3052 8446 3088
rect 8390 3032 8392 3052
rect 8392 3032 8444 3052
rect 8444 3032 8446 3052
rect 9678 7520 9734 7576
rect 10414 8880 10470 8936
rect 10138 6160 10194 6216
rect 9954 2760 10010 2816
rect 18970 29552 19026 29608
rect 21914 17992 21970 18048
rect 14554 14456 14610 14512
rect 11978 9016 12034 9072
rect 11702 8608 11758 8664
rect 10230 3476 10232 3496
rect 10232 3476 10284 3496
rect 10284 3476 10286 3496
rect 10230 3440 10286 3476
rect 10506 2916 10562 2952
rect 10506 2896 10508 2916
rect 10508 2896 10560 2916
rect 10560 2896 10562 2916
rect 10414 2624 10470 2680
rect 10874 4020 10876 4040
rect 10876 4020 10928 4040
rect 10928 4020 10930 4040
rect 10874 3984 10930 4020
rect 11334 3304 11390 3360
rect 12162 5616 12218 5672
rect 11702 4020 11704 4040
rect 11704 4020 11756 4040
rect 11756 4020 11758 4040
rect 11702 3984 11758 4020
rect 11702 3848 11758 3904
rect 12714 6316 12770 6352
rect 12714 6296 12716 6316
rect 12716 6296 12768 6316
rect 12768 6296 12770 6316
rect 12714 6060 12716 6080
rect 12716 6060 12768 6080
rect 12768 6060 12770 6080
rect 12714 6024 12770 6060
rect 12622 4820 12678 4856
rect 12622 4800 12624 4820
rect 12624 4800 12676 4820
rect 12676 4800 12678 4820
rect 12622 4664 12678 4720
rect 12714 3304 12770 3360
rect 13542 9696 13598 9752
rect 13450 9288 13506 9344
rect 13174 5208 13230 5264
rect 12990 3848 13046 3904
rect 13542 3576 13598 3632
rect 14094 5888 14150 5944
rect 13634 3304 13690 3360
rect 14094 4936 14150 4992
rect 14278 3712 14334 3768
rect 14002 3576 14058 3632
rect 13910 2896 13966 2952
rect 15106 5616 15162 5672
rect 15290 5636 15346 5672
rect 15290 5616 15292 5636
rect 15292 5616 15344 5636
rect 15344 5616 15346 5636
rect 15198 5364 15254 5400
rect 15198 5344 15200 5364
rect 15200 5344 15252 5364
rect 15252 5344 15254 5364
rect 15014 4392 15070 4448
rect 15106 4120 15162 4176
rect 15658 9424 15714 9480
rect 15750 8336 15806 8392
rect 15658 6840 15714 6896
rect 15566 6296 15622 6352
rect 15474 3168 15530 3224
rect 15842 6840 15898 6896
rect 16118 6296 16174 6352
rect 16394 6024 16450 6080
rect 16302 5772 16358 5808
rect 16302 5752 16304 5772
rect 16304 5752 16356 5772
rect 16356 5752 16358 5772
rect 17038 4820 17094 4856
rect 17038 4800 17040 4820
rect 17040 4800 17092 4820
rect 17092 4800 17094 4820
rect 16854 4528 16910 4584
rect 15658 3304 15714 3360
rect 15934 3304 15990 3360
rect 16946 3848 17002 3904
rect 16854 3168 16910 3224
rect 24674 12144 24730 12200
rect 18234 8744 18290 8800
rect 17682 5228 17738 5264
rect 17682 5208 17684 5228
rect 17684 5208 17736 5228
rect 17736 5208 17738 5228
rect 17682 4800 17738 4856
rect 17958 2760 18014 2816
rect 18602 8472 18658 8528
rect 18694 8336 18750 8392
rect 17406 1264 17462 1320
rect 18602 6024 18658 6080
rect 18602 5480 18658 5536
rect 18694 5072 18750 5128
rect 18510 4256 18566 4312
rect 19982 10512 20038 10568
rect 19338 9016 19394 9072
rect 19614 9016 19670 9072
rect 19430 7284 19432 7304
rect 19432 7284 19484 7304
rect 19484 7284 19486 7304
rect 19430 7248 19486 7284
rect 19246 6296 19302 6352
rect 19338 6160 19394 6216
rect 19890 8608 19946 8664
rect 19614 6740 19616 6760
rect 19616 6740 19668 6760
rect 19668 6740 19670 6760
rect 19614 6704 19670 6740
rect 19430 5752 19486 5808
rect 19522 5344 19578 5400
rect 19430 4800 19486 4856
rect 19154 4528 19210 4584
rect 19982 8472 20038 8528
rect 19062 4120 19118 4176
rect 19338 4156 19340 4176
rect 19340 4156 19392 4176
rect 19392 4156 19394 4176
rect 19338 4120 19394 4156
rect 19706 4528 19762 4584
rect 19614 4120 19670 4176
rect 20074 7928 20130 7984
rect 20074 5208 20130 5264
rect 19982 4428 19984 4448
rect 19984 4428 20036 4448
rect 20036 4428 20038 4448
rect 19982 4392 20038 4428
rect 21638 10920 21694 10976
rect 20442 8900 20498 8936
rect 20442 8880 20444 8900
rect 20444 8880 20496 8900
rect 20496 8880 20498 8900
rect 20350 5228 20406 5264
rect 20350 5208 20352 5228
rect 20352 5208 20404 5228
rect 20404 5208 20406 5228
rect 20718 6840 20774 6896
rect 20902 8200 20958 8256
rect 20902 6976 20958 7032
rect 19522 3032 19578 3088
rect 19890 3032 19946 3088
rect 20534 4120 20590 4176
rect 19338 2508 19394 2544
rect 19338 2488 19340 2508
rect 19340 2488 19392 2508
rect 19392 2488 19394 2508
rect 22466 11192 22522 11248
rect 21546 10240 21602 10296
rect 21362 9968 21418 10024
rect 21362 9868 21364 9888
rect 21364 9868 21416 9888
rect 21416 9868 21418 9888
rect 21362 9832 21418 9868
rect 21270 9016 21326 9072
rect 21178 8356 21234 8392
rect 21178 8336 21180 8356
rect 21180 8336 21232 8356
rect 21232 8336 21234 8356
rect 20902 4664 20958 4720
rect 21454 7520 21510 7576
rect 21730 7520 21786 7576
rect 21362 5752 21418 5808
rect 21178 4800 21234 4856
rect 20718 2216 20774 2272
rect 20902 3440 20958 3496
rect 21454 5344 21510 5400
rect 21822 6568 21878 6624
rect 21546 3984 21602 4040
rect 21822 4528 21878 4584
rect 21362 3848 21418 3904
rect 21546 1672 21602 1728
rect 19982 1400 20038 1456
rect 20810 1400 20866 1456
rect 19338 1264 19394 1320
rect 18602 1128 18658 1184
rect 21730 3068 21732 3088
rect 21732 3068 21784 3088
rect 21784 3068 21786 3088
rect 21730 3032 21786 3068
rect 22006 7284 22008 7304
rect 22008 7284 22060 7304
rect 22060 7284 22062 7304
rect 22006 7248 22062 7284
rect 22374 7384 22430 7440
rect 22374 6860 22430 6896
rect 22374 6840 22376 6860
rect 22376 6840 22428 6860
rect 22428 6840 22430 6860
rect 22190 6740 22192 6760
rect 22192 6740 22244 6760
rect 22244 6740 22246 6760
rect 22190 6704 22246 6740
rect 22374 6704 22430 6760
rect 22006 6432 22062 6488
rect 22282 6432 22338 6488
rect 22098 5344 22154 5400
rect 22098 4428 22100 4448
rect 22100 4428 22152 4448
rect 22152 4428 22154 4448
rect 22098 4392 22154 4428
rect 22098 3984 22154 4040
rect 22006 3304 22062 3360
rect 22282 5344 22338 5400
rect 22282 4564 22284 4584
rect 22284 4564 22336 4584
rect 22336 4564 22338 4584
rect 22282 4528 22338 4564
rect 22282 3168 22338 3224
rect 22558 7928 22614 7984
rect 22558 6976 22614 7032
rect 22926 9560 22982 9616
rect 23478 11056 23534 11112
rect 23386 10512 23442 10568
rect 23478 10004 23480 10024
rect 23480 10004 23532 10024
rect 23532 10004 23534 10024
rect 23478 9968 23534 10004
rect 23386 9832 23442 9888
rect 23294 9696 23350 9752
rect 22834 8880 22890 8936
rect 22834 7384 22890 7440
rect 22742 6840 22798 6896
rect 23386 9288 23442 9344
rect 23570 9152 23626 9208
rect 22650 4020 22652 4040
rect 22652 4020 22704 4040
rect 22704 4020 22706 4040
rect 22650 3984 22706 4020
rect 23478 7656 23534 7712
rect 23202 4664 23258 4720
rect 23294 2896 23350 2952
rect 22558 1400 22614 1456
rect 23754 5888 23810 5944
rect 24398 10512 24454 10568
rect 24306 8472 24362 8528
rect 24122 7948 24178 7984
rect 24122 7928 24124 7948
rect 24124 7928 24176 7948
rect 24176 7928 24178 7948
rect 23938 7656 23994 7712
rect 23754 5652 23756 5672
rect 23756 5652 23808 5672
rect 23808 5652 23810 5672
rect 23754 5616 23810 5652
rect 23662 4664 23718 4720
rect 23846 4936 23902 4992
rect 23754 3712 23810 3768
rect 24950 11092 24952 11112
rect 24952 11092 25004 11112
rect 25004 11092 25006 11112
rect 24950 11056 25006 11092
rect 24490 9288 24546 9344
rect 24490 8064 24546 8120
rect 24674 9444 24730 9480
rect 24674 9424 24676 9444
rect 24676 9424 24728 9444
rect 24728 9424 24730 9444
rect 25686 12144 25742 12200
rect 25778 10512 25834 10568
rect 35860 37562 35916 37564
rect 35940 37562 35996 37564
rect 36020 37562 36076 37564
rect 36100 37562 36156 37564
rect 35860 37510 35906 37562
rect 35906 37510 35916 37562
rect 35940 37510 35970 37562
rect 35970 37510 35982 37562
rect 35982 37510 35996 37562
rect 36020 37510 36034 37562
rect 36034 37510 36046 37562
rect 36046 37510 36076 37562
rect 36100 37510 36110 37562
rect 36110 37510 36156 37562
rect 35860 37508 35916 37510
rect 35940 37508 35996 37510
rect 36020 37508 36076 37510
rect 36100 37508 36156 37510
rect 36520 37018 36576 37020
rect 36600 37018 36656 37020
rect 36680 37018 36736 37020
rect 36760 37018 36816 37020
rect 36520 36966 36566 37018
rect 36566 36966 36576 37018
rect 36600 36966 36630 37018
rect 36630 36966 36642 37018
rect 36642 36966 36656 37018
rect 36680 36966 36694 37018
rect 36694 36966 36706 37018
rect 36706 36966 36736 37018
rect 36760 36966 36770 37018
rect 36770 36966 36816 37018
rect 36520 36964 36576 36966
rect 36600 36964 36656 36966
rect 36680 36964 36736 36966
rect 36760 36964 36816 36966
rect 32770 36488 32826 36544
rect 35860 36474 35916 36476
rect 35940 36474 35996 36476
rect 36020 36474 36076 36476
rect 36100 36474 36156 36476
rect 35860 36422 35906 36474
rect 35906 36422 35916 36474
rect 35940 36422 35970 36474
rect 35970 36422 35982 36474
rect 35982 36422 35996 36474
rect 36020 36422 36034 36474
rect 36034 36422 36046 36474
rect 36046 36422 36076 36474
rect 36100 36422 36110 36474
rect 36110 36422 36156 36474
rect 35860 36420 35916 36422
rect 35940 36420 35996 36422
rect 36020 36420 36076 36422
rect 36100 36420 36156 36422
rect 36520 35930 36576 35932
rect 36600 35930 36656 35932
rect 36680 35930 36736 35932
rect 36760 35930 36816 35932
rect 36520 35878 36566 35930
rect 36566 35878 36576 35930
rect 36600 35878 36630 35930
rect 36630 35878 36642 35930
rect 36642 35878 36656 35930
rect 36680 35878 36694 35930
rect 36694 35878 36706 35930
rect 36706 35878 36736 35930
rect 36760 35878 36770 35930
rect 36770 35878 36816 35930
rect 36520 35876 36576 35878
rect 36600 35876 36656 35878
rect 36680 35876 36736 35878
rect 36760 35876 36816 35878
rect 35860 35386 35916 35388
rect 35940 35386 35996 35388
rect 36020 35386 36076 35388
rect 36100 35386 36156 35388
rect 35860 35334 35906 35386
rect 35906 35334 35916 35386
rect 35940 35334 35970 35386
rect 35970 35334 35982 35386
rect 35982 35334 35996 35386
rect 36020 35334 36034 35386
rect 36034 35334 36046 35386
rect 36046 35334 36076 35386
rect 36100 35334 36110 35386
rect 36110 35334 36156 35386
rect 35860 35332 35916 35334
rect 35940 35332 35996 35334
rect 36020 35332 36076 35334
rect 36100 35332 36156 35334
rect 36520 34842 36576 34844
rect 36600 34842 36656 34844
rect 36680 34842 36736 34844
rect 36760 34842 36816 34844
rect 36520 34790 36566 34842
rect 36566 34790 36576 34842
rect 36600 34790 36630 34842
rect 36630 34790 36642 34842
rect 36642 34790 36656 34842
rect 36680 34790 36694 34842
rect 36694 34790 36706 34842
rect 36706 34790 36736 34842
rect 36760 34790 36770 34842
rect 36770 34790 36816 34842
rect 36520 34788 36576 34790
rect 36600 34788 36656 34790
rect 36680 34788 36736 34790
rect 36760 34788 36816 34790
rect 35860 34298 35916 34300
rect 35940 34298 35996 34300
rect 36020 34298 36076 34300
rect 36100 34298 36156 34300
rect 35860 34246 35906 34298
rect 35906 34246 35916 34298
rect 35940 34246 35970 34298
rect 35970 34246 35982 34298
rect 35982 34246 35996 34298
rect 36020 34246 36034 34298
rect 36034 34246 36046 34298
rect 36046 34246 36076 34298
rect 36100 34246 36110 34298
rect 36110 34246 36156 34298
rect 35860 34244 35916 34246
rect 35940 34244 35996 34246
rect 36020 34244 36076 34246
rect 36100 34244 36156 34246
rect 36520 33754 36576 33756
rect 36600 33754 36656 33756
rect 36680 33754 36736 33756
rect 36760 33754 36816 33756
rect 36520 33702 36566 33754
rect 36566 33702 36576 33754
rect 36600 33702 36630 33754
rect 36630 33702 36642 33754
rect 36642 33702 36656 33754
rect 36680 33702 36694 33754
rect 36694 33702 36706 33754
rect 36706 33702 36736 33754
rect 36760 33702 36770 33754
rect 36770 33702 36816 33754
rect 36520 33700 36576 33702
rect 36600 33700 36656 33702
rect 36680 33700 36736 33702
rect 36760 33700 36816 33702
rect 35860 33210 35916 33212
rect 35940 33210 35996 33212
rect 36020 33210 36076 33212
rect 36100 33210 36156 33212
rect 35860 33158 35906 33210
rect 35906 33158 35916 33210
rect 35940 33158 35970 33210
rect 35970 33158 35982 33210
rect 35982 33158 35996 33210
rect 36020 33158 36034 33210
rect 36034 33158 36046 33210
rect 36046 33158 36076 33210
rect 36100 33158 36110 33210
rect 36110 33158 36156 33210
rect 35860 33156 35916 33158
rect 35940 33156 35996 33158
rect 36020 33156 36076 33158
rect 36100 33156 36156 33158
rect 36520 32666 36576 32668
rect 36600 32666 36656 32668
rect 36680 32666 36736 32668
rect 36760 32666 36816 32668
rect 36520 32614 36566 32666
rect 36566 32614 36576 32666
rect 36600 32614 36630 32666
rect 36630 32614 36642 32666
rect 36642 32614 36656 32666
rect 36680 32614 36694 32666
rect 36694 32614 36706 32666
rect 36706 32614 36736 32666
rect 36760 32614 36770 32666
rect 36770 32614 36816 32666
rect 36520 32612 36576 32614
rect 36600 32612 36656 32614
rect 36680 32612 36736 32614
rect 36760 32612 36816 32614
rect 35860 32122 35916 32124
rect 35940 32122 35996 32124
rect 36020 32122 36076 32124
rect 36100 32122 36156 32124
rect 35860 32070 35906 32122
rect 35906 32070 35916 32122
rect 35940 32070 35970 32122
rect 35970 32070 35982 32122
rect 35982 32070 35996 32122
rect 36020 32070 36034 32122
rect 36034 32070 36046 32122
rect 36046 32070 36076 32122
rect 36100 32070 36110 32122
rect 36110 32070 36156 32122
rect 35860 32068 35916 32070
rect 35940 32068 35996 32070
rect 36020 32068 36076 32070
rect 36100 32068 36156 32070
rect 36520 31578 36576 31580
rect 36600 31578 36656 31580
rect 36680 31578 36736 31580
rect 36760 31578 36816 31580
rect 36520 31526 36566 31578
rect 36566 31526 36576 31578
rect 36600 31526 36630 31578
rect 36630 31526 36642 31578
rect 36642 31526 36656 31578
rect 36680 31526 36694 31578
rect 36694 31526 36706 31578
rect 36706 31526 36736 31578
rect 36760 31526 36770 31578
rect 36770 31526 36816 31578
rect 36520 31524 36576 31526
rect 36600 31524 36656 31526
rect 36680 31524 36736 31526
rect 36760 31524 36816 31526
rect 35860 31034 35916 31036
rect 35940 31034 35996 31036
rect 36020 31034 36076 31036
rect 36100 31034 36156 31036
rect 35860 30982 35906 31034
rect 35906 30982 35916 31034
rect 35940 30982 35970 31034
rect 35970 30982 35982 31034
rect 35982 30982 35996 31034
rect 36020 30982 36034 31034
rect 36034 30982 36046 31034
rect 36046 30982 36076 31034
rect 36100 30982 36110 31034
rect 36110 30982 36156 31034
rect 35860 30980 35916 30982
rect 35940 30980 35996 30982
rect 36020 30980 36076 30982
rect 36100 30980 36156 30982
rect 36520 30490 36576 30492
rect 36600 30490 36656 30492
rect 36680 30490 36736 30492
rect 36760 30490 36816 30492
rect 36520 30438 36566 30490
rect 36566 30438 36576 30490
rect 36600 30438 36630 30490
rect 36630 30438 36642 30490
rect 36642 30438 36656 30490
rect 36680 30438 36694 30490
rect 36694 30438 36706 30490
rect 36706 30438 36736 30490
rect 36760 30438 36770 30490
rect 36770 30438 36816 30490
rect 36520 30436 36576 30438
rect 36600 30436 36656 30438
rect 36680 30436 36736 30438
rect 36760 30436 36816 30438
rect 35860 29946 35916 29948
rect 35940 29946 35996 29948
rect 36020 29946 36076 29948
rect 36100 29946 36156 29948
rect 35860 29894 35906 29946
rect 35906 29894 35916 29946
rect 35940 29894 35970 29946
rect 35970 29894 35982 29946
rect 35982 29894 35996 29946
rect 36020 29894 36034 29946
rect 36034 29894 36046 29946
rect 36046 29894 36076 29946
rect 36100 29894 36110 29946
rect 36110 29894 36156 29946
rect 35860 29892 35916 29894
rect 35940 29892 35996 29894
rect 36020 29892 36076 29894
rect 36100 29892 36156 29894
rect 36520 29402 36576 29404
rect 36600 29402 36656 29404
rect 36680 29402 36736 29404
rect 36760 29402 36816 29404
rect 36520 29350 36566 29402
rect 36566 29350 36576 29402
rect 36600 29350 36630 29402
rect 36630 29350 36642 29402
rect 36642 29350 36656 29402
rect 36680 29350 36694 29402
rect 36694 29350 36706 29402
rect 36706 29350 36736 29402
rect 36760 29350 36770 29402
rect 36770 29350 36816 29402
rect 36520 29348 36576 29350
rect 36600 29348 36656 29350
rect 36680 29348 36736 29350
rect 36760 29348 36816 29350
rect 35860 28858 35916 28860
rect 35940 28858 35996 28860
rect 36020 28858 36076 28860
rect 36100 28858 36156 28860
rect 35860 28806 35906 28858
rect 35906 28806 35916 28858
rect 35940 28806 35970 28858
rect 35970 28806 35982 28858
rect 35982 28806 35996 28858
rect 36020 28806 36034 28858
rect 36034 28806 36046 28858
rect 36046 28806 36076 28858
rect 36100 28806 36110 28858
rect 36110 28806 36156 28858
rect 35860 28804 35916 28806
rect 35940 28804 35996 28806
rect 36020 28804 36076 28806
rect 36100 28804 36156 28806
rect 36520 28314 36576 28316
rect 36600 28314 36656 28316
rect 36680 28314 36736 28316
rect 36760 28314 36816 28316
rect 36520 28262 36566 28314
rect 36566 28262 36576 28314
rect 36600 28262 36630 28314
rect 36630 28262 36642 28314
rect 36642 28262 36656 28314
rect 36680 28262 36694 28314
rect 36694 28262 36706 28314
rect 36706 28262 36736 28314
rect 36760 28262 36770 28314
rect 36770 28262 36816 28314
rect 36520 28260 36576 28262
rect 36600 28260 36656 28262
rect 36680 28260 36736 28262
rect 36760 28260 36816 28262
rect 35860 27770 35916 27772
rect 35940 27770 35996 27772
rect 36020 27770 36076 27772
rect 36100 27770 36156 27772
rect 35860 27718 35906 27770
rect 35906 27718 35916 27770
rect 35940 27718 35970 27770
rect 35970 27718 35982 27770
rect 35982 27718 35996 27770
rect 36020 27718 36034 27770
rect 36034 27718 36046 27770
rect 36046 27718 36076 27770
rect 36100 27718 36110 27770
rect 36110 27718 36156 27770
rect 35860 27716 35916 27718
rect 35940 27716 35996 27718
rect 36020 27716 36076 27718
rect 36100 27716 36156 27718
rect 36520 27226 36576 27228
rect 36600 27226 36656 27228
rect 36680 27226 36736 27228
rect 36760 27226 36816 27228
rect 36520 27174 36566 27226
rect 36566 27174 36576 27226
rect 36600 27174 36630 27226
rect 36630 27174 36642 27226
rect 36642 27174 36656 27226
rect 36680 27174 36694 27226
rect 36694 27174 36706 27226
rect 36706 27174 36736 27226
rect 36760 27174 36770 27226
rect 36770 27174 36816 27226
rect 36520 27172 36576 27174
rect 36600 27172 36656 27174
rect 36680 27172 36736 27174
rect 36760 27172 36816 27174
rect 35860 26682 35916 26684
rect 35940 26682 35996 26684
rect 36020 26682 36076 26684
rect 36100 26682 36156 26684
rect 35860 26630 35906 26682
rect 35906 26630 35916 26682
rect 35940 26630 35970 26682
rect 35970 26630 35982 26682
rect 35982 26630 35996 26682
rect 36020 26630 36034 26682
rect 36034 26630 36046 26682
rect 36046 26630 36076 26682
rect 36100 26630 36110 26682
rect 36110 26630 36156 26682
rect 35860 26628 35916 26630
rect 35940 26628 35996 26630
rect 36020 26628 36076 26630
rect 36100 26628 36156 26630
rect 36520 26138 36576 26140
rect 36600 26138 36656 26140
rect 36680 26138 36736 26140
rect 36760 26138 36816 26140
rect 36520 26086 36566 26138
rect 36566 26086 36576 26138
rect 36600 26086 36630 26138
rect 36630 26086 36642 26138
rect 36642 26086 36656 26138
rect 36680 26086 36694 26138
rect 36694 26086 36706 26138
rect 36706 26086 36736 26138
rect 36760 26086 36770 26138
rect 36770 26086 36816 26138
rect 36520 26084 36576 26086
rect 36600 26084 36656 26086
rect 36680 26084 36736 26086
rect 36760 26084 36816 26086
rect 35860 25594 35916 25596
rect 35940 25594 35996 25596
rect 36020 25594 36076 25596
rect 36100 25594 36156 25596
rect 35860 25542 35906 25594
rect 35906 25542 35916 25594
rect 35940 25542 35970 25594
rect 35970 25542 35982 25594
rect 35982 25542 35996 25594
rect 36020 25542 36034 25594
rect 36034 25542 36046 25594
rect 36046 25542 36076 25594
rect 36100 25542 36110 25594
rect 36110 25542 36156 25594
rect 35860 25540 35916 25542
rect 35940 25540 35996 25542
rect 36020 25540 36076 25542
rect 36100 25540 36156 25542
rect 36520 25050 36576 25052
rect 36600 25050 36656 25052
rect 36680 25050 36736 25052
rect 36760 25050 36816 25052
rect 36520 24998 36566 25050
rect 36566 24998 36576 25050
rect 36600 24998 36630 25050
rect 36630 24998 36642 25050
rect 36642 24998 36656 25050
rect 36680 24998 36694 25050
rect 36694 24998 36706 25050
rect 36706 24998 36736 25050
rect 36760 24998 36770 25050
rect 36770 24998 36816 25050
rect 36520 24996 36576 24998
rect 36600 24996 36656 24998
rect 36680 24996 36736 24998
rect 36760 24996 36816 24998
rect 35860 24506 35916 24508
rect 35940 24506 35996 24508
rect 36020 24506 36076 24508
rect 36100 24506 36156 24508
rect 35860 24454 35906 24506
rect 35906 24454 35916 24506
rect 35940 24454 35970 24506
rect 35970 24454 35982 24506
rect 35982 24454 35996 24506
rect 36020 24454 36034 24506
rect 36034 24454 36046 24506
rect 36046 24454 36076 24506
rect 36100 24454 36110 24506
rect 36110 24454 36156 24506
rect 35860 24452 35916 24454
rect 35940 24452 35996 24454
rect 36020 24452 36076 24454
rect 36100 24452 36156 24454
rect 36520 23962 36576 23964
rect 36600 23962 36656 23964
rect 36680 23962 36736 23964
rect 36760 23962 36816 23964
rect 36520 23910 36566 23962
rect 36566 23910 36576 23962
rect 36600 23910 36630 23962
rect 36630 23910 36642 23962
rect 36642 23910 36656 23962
rect 36680 23910 36694 23962
rect 36694 23910 36706 23962
rect 36706 23910 36736 23962
rect 36760 23910 36770 23962
rect 36770 23910 36816 23962
rect 36520 23908 36576 23910
rect 36600 23908 36656 23910
rect 36680 23908 36736 23910
rect 36760 23908 36816 23910
rect 35860 23418 35916 23420
rect 35940 23418 35996 23420
rect 36020 23418 36076 23420
rect 36100 23418 36156 23420
rect 35860 23366 35906 23418
rect 35906 23366 35916 23418
rect 35940 23366 35970 23418
rect 35970 23366 35982 23418
rect 35982 23366 35996 23418
rect 36020 23366 36034 23418
rect 36034 23366 36046 23418
rect 36046 23366 36076 23418
rect 36100 23366 36110 23418
rect 36110 23366 36156 23418
rect 35860 23364 35916 23366
rect 35940 23364 35996 23366
rect 36020 23364 36076 23366
rect 36100 23364 36156 23366
rect 36520 22874 36576 22876
rect 36600 22874 36656 22876
rect 36680 22874 36736 22876
rect 36760 22874 36816 22876
rect 36520 22822 36566 22874
rect 36566 22822 36576 22874
rect 36600 22822 36630 22874
rect 36630 22822 36642 22874
rect 36642 22822 36656 22874
rect 36680 22822 36694 22874
rect 36694 22822 36706 22874
rect 36706 22822 36736 22874
rect 36760 22822 36770 22874
rect 36770 22822 36816 22874
rect 36520 22820 36576 22822
rect 36600 22820 36656 22822
rect 36680 22820 36736 22822
rect 36760 22820 36816 22822
rect 35860 22330 35916 22332
rect 35940 22330 35996 22332
rect 36020 22330 36076 22332
rect 36100 22330 36156 22332
rect 35860 22278 35906 22330
rect 35906 22278 35916 22330
rect 35940 22278 35970 22330
rect 35970 22278 35982 22330
rect 35982 22278 35996 22330
rect 36020 22278 36034 22330
rect 36034 22278 36046 22330
rect 36046 22278 36076 22330
rect 36100 22278 36110 22330
rect 36110 22278 36156 22330
rect 35860 22276 35916 22278
rect 35940 22276 35996 22278
rect 36020 22276 36076 22278
rect 36100 22276 36156 22278
rect 36520 21786 36576 21788
rect 36600 21786 36656 21788
rect 36680 21786 36736 21788
rect 36760 21786 36816 21788
rect 36520 21734 36566 21786
rect 36566 21734 36576 21786
rect 36600 21734 36630 21786
rect 36630 21734 36642 21786
rect 36642 21734 36656 21786
rect 36680 21734 36694 21786
rect 36694 21734 36706 21786
rect 36706 21734 36736 21786
rect 36760 21734 36770 21786
rect 36770 21734 36816 21786
rect 36520 21732 36576 21734
rect 36600 21732 36656 21734
rect 36680 21732 36736 21734
rect 36760 21732 36816 21734
rect 35860 21242 35916 21244
rect 35940 21242 35996 21244
rect 36020 21242 36076 21244
rect 36100 21242 36156 21244
rect 35860 21190 35906 21242
rect 35906 21190 35916 21242
rect 35940 21190 35970 21242
rect 35970 21190 35982 21242
rect 35982 21190 35996 21242
rect 36020 21190 36034 21242
rect 36034 21190 36046 21242
rect 36046 21190 36076 21242
rect 36100 21190 36110 21242
rect 36110 21190 36156 21242
rect 35860 21188 35916 21190
rect 35940 21188 35996 21190
rect 36020 21188 36076 21190
rect 36100 21188 36156 21190
rect 36520 20698 36576 20700
rect 36600 20698 36656 20700
rect 36680 20698 36736 20700
rect 36760 20698 36816 20700
rect 36520 20646 36566 20698
rect 36566 20646 36576 20698
rect 36600 20646 36630 20698
rect 36630 20646 36642 20698
rect 36642 20646 36656 20698
rect 36680 20646 36694 20698
rect 36694 20646 36706 20698
rect 36706 20646 36736 20698
rect 36760 20646 36770 20698
rect 36770 20646 36816 20698
rect 36520 20644 36576 20646
rect 36600 20644 36656 20646
rect 36680 20644 36736 20646
rect 36760 20644 36816 20646
rect 35860 20154 35916 20156
rect 35940 20154 35996 20156
rect 36020 20154 36076 20156
rect 36100 20154 36156 20156
rect 35860 20102 35906 20154
rect 35906 20102 35916 20154
rect 35940 20102 35970 20154
rect 35970 20102 35982 20154
rect 35982 20102 35996 20154
rect 36020 20102 36034 20154
rect 36034 20102 36046 20154
rect 36046 20102 36076 20154
rect 36100 20102 36110 20154
rect 36110 20102 36156 20154
rect 35860 20100 35916 20102
rect 35940 20100 35996 20102
rect 36020 20100 36076 20102
rect 36100 20100 36156 20102
rect 36520 19610 36576 19612
rect 36600 19610 36656 19612
rect 36680 19610 36736 19612
rect 36760 19610 36816 19612
rect 36520 19558 36566 19610
rect 36566 19558 36576 19610
rect 36600 19558 36630 19610
rect 36630 19558 36642 19610
rect 36642 19558 36656 19610
rect 36680 19558 36694 19610
rect 36694 19558 36706 19610
rect 36706 19558 36736 19610
rect 36760 19558 36770 19610
rect 36770 19558 36816 19610
rect 36520 19556 36576 19558
rect 36600 19556 36656 19558
rect 36680 19556 36736 19558
rect 36760 19556 36816 19558
rect 35860 19066 35916 19068
rect 35940 19066 35996 19068
rect 36020 19066 36076 19068
rect 36100 19066 36156 19068
rect 35860 19014 35906 19066
rect 35906 19014 35916 19066
rect 35940 19014 35970 19066
rect 35970 19014 35982 19066
rect 35982 19014 35996 19066
rect 36020 19014 36034 19066
rect 36034 19014 36046 19066
rect 36046 19014 36076 19066
rect 36100 19014 36110 19066
rect 36110 19014 36156 19066
rect 35860 19012 35916 19014
rect 35940 19012 35996 19014
rect 36020 19012 36076 19014
rect 36100 19012 36156 19014
rect 36520 18522 36576 18524
rect 36600 18522 36656 18524
rect 36680 18522 36736 18524
rect 36760 18522 36816 18524
rect 36520 18470 36566 18522
rect 36566 18470 36576 18522
rect 36600 18470 36630 18522
rect 36630 18470 36642 18522
rect 36642 18470 36656 18522
rect 36680 18470 36694 18522
rect 36694 18470 36706 18522
rect 36706 18470 36736 18522
rect 36760 18470 36770 18522
rect 36770 18470 36816 18522
rect 36520 18468 36576 18470
rect 36600 18468 36656 18470
rect 36680 18468 36736 18470
rect 36760 18468 36816 18470
rect 35860 17978 35916 17980
rect 35940 17978 35996 17980
rect 36020 17978 36076 17980
rect 36100 17978 36156 17980
rect 35860 17926 35906 17978
rect 35906 17926 35916 17978
rect 35940 17926 35970 17978
rect 35970 17926 35982 17978
rect 35982 17926 35996 17978
rect 36020 17926 36034 17978
rect 36034 17926 36046 17978
rect 36046 17926 36076 17978
rect 36100 17926 36110 17978
rect 36110 17926 36156 17978
rect 35860 17924 35916 17926
rect 35940 17924 35996 17926
rect 36020 17924 36076 17926
rect 36100 17924 36156 17926
rect 36520 17434 36576 17436
rect 36600 17434 36656 17436
rect 36680 17434 36736 17436
rect 36760 17434 36816 17436
rect 36520 17382 36566 17434
rect 36566 17382 36576 17434
rect 36600 17382 36630 17434
rect 36630 17382 36642 17434
rect 36642 17382 36656 17434
rect 36680 17382 36694 17434
rect 36694 17382 36706 17434
rect 36706 17382 36736 17434
rect 36760 17382 36770 17434
rect 36770 17382 36816 17434
rect 36520 17380 36576 17382
rect 36600 17380 36656 17382
rect 36680 17380 36736 17382
rect 36760 17380 36816 17382
rect 35860 16890 35916 16892
rect 35940 16890 35996 16892
rect 36020 16890 36076 16892
rect 36100 16890 36156 16892
rect 35860 16838 35906 16890
rect 35906 16838 35916 16890
rect 35940 16838 35970 16890
rect 35970 16838 35982 16890
rect 35982 16838 35996 16890
rect 36020 16838 36034 16890
rect 36034 16838 36046 16890
rect 36046 16838 36076 16890
rect 36100 16838 36110 16890
rect 36110 16838 36156 16890
rect 35860 16836 35916 16838
rect 35940 16836 35996 16838
rect 36020 16836 36076 16838
rect 36100 16836 36156 16838
rect 26238 10548 26240 10568
rect 26240 10548 26292 10568
rect 26292 10548 26294 10568
rect 26238 10512 26294 10548
rect 25594 9696 25650 9752
rect 25042 8472 25098 8528
rect 25042 7520 25098 7576
rect 24398 2624 24454 2680
rect 23662 1400 23718 1456
rect 23846 1128 23902 1184
rect 24582 3052 24638 3088
rect 24582 3032 24584 3052
rect 24584 3032 24636 3052
rect 24636 3032 24638 3052
rect 24858 3576 24914 3632
rect 25042 5072 25098 5128
rect 25042 3440 25098 3496
rect 25502 8336 25558 8392
rect 25318 6840 25374 6896
rect 25410 5208 25466 5264
rect 25410 4972 25412 4992
rect 25412 4972 25464 4992
rect 25464 4972 25466 4992
rect 25410 4936 25466 4972
rect 25318 3712 25374 3768
rect 25502 4120 25558 4176
rect 25686 5752 25742 5808
rect 25134 3032 25190 3088
rect 25226 2796 25228 2816
rect 25228 2796 25280 2816
rect 25280 2796 25282 2816
rect 25226 2760 25282 2796
rect 25410 3340 25412 3360
rect 25412 3340 25464 3360
rect 25464 3340 25466 3360
rect 25410 3304 25466 3340
rect 25410 3032 25466 3088
rect 25318 2488 25374 2544
rect 24582 2388 24584 2408
rect 24584 2388 24636 2408
rect 24636 2388 24638 2408
rect 24582 2352 24638 2388
rect 25962 4020 25964 4040
rect 25964 4020 26016 4040
rect 26016 4020 26018 4040
rect 25962 3984 26018 4020
rect 26238 8608 26294 8664
rect 26330 8472 26386 8528
rect 26238 6432 26294 6488
rect 26330 5344 26386 5400
rect 26514 6316 26570 6352
rect 26514 6296 26516 6316
rect 26516 6296 26568 6316
rect 26568 6296 26570 6316
rect 27710 12416 27766 12472
rect 26974 9696 27030 9752
rect 26882 8508 26884 8528
rect 26884 8508 26936 8528
rect 26936 8508 26938 8528
rect 26882 8472 26938 8508
rect 27066 8472 27122 8528
rect 26974 7656 27030 7712
rect 27158 8336 27214 8392
rect 27158 8064 27214 8120
rect 27158 7384 27214 7440
rect 26238 2216 26294 2272
rect 27158 7112 27214 7168
rect 26790 6976 26846 7032
rect 26698 4004 26754 4040
rect 26698 3984 26700 4004
rect 26700 3984 26752 4004
rect 26752 3984 26754 4004
rect 27158 5208 27214 5264
rect 26698 3340 26700 3360
rect 26700 3340 26752 3360
rect 26752 3340 26754 3360
rect 26698 3304 26754 3340
rect 25778 992 25834 1048
rect 27066 3576 27122 3632
rect 27986 11328 28042 11384
rect 27986 9968 28042 10024
rect 27434 8900 27490 8936
rect 27434 8880 27436 8900
rect 27436 8880 27488 8900
rect 27488 8880 27490 8900
rect 27710 8744 27766 8800
rect 27710 8336 27766 8392
rect 27526 8200 27582 8256
rect 27618 7928 27674 7984
rect 27434 7656 27490 7712
rect 27526 7520 27582 7576
rect 27434 5208 27490 5264
rect 28170 11464 28226 11520
rect 28170 10920 28226 10976
rect 27710 5480 27766 5536
rect 27342 3052 27398 3088
rect 27342 3032 27344 3052
rect 27344 3032 27396 3052
rect 27396 3032 27398 3052
rect 28630 10412 28632 10432
rect 28632 10412 28684 10432
rect 28684 10412 28686 10432
rect 28630 10376 28686 10412
rect 28170 7792 28226 7848
rect 28078 7248 28134 7304
rect 27986 6568 28042 6624
rect 27986 5208 28042 5264
rect 28262 5888 28318 5944
rect 28078 3576 28134 3632
rect 28630 9016 28686 9072
rect 28630 7928 28686 7984
rect 28814 10784 28870 10840
rect 28446 6160 28502 6216
rect 28446 4256 28502 4312
rect 28078 1808 28134 1864
rect 28630 6432 28686 6488
rect 29182 10376 29238 10432
rect 28998 9560 29054 9616
rect 29182 8744 29238 8800
rect 29090 5752 29146 5808
rect 28998 4936 29054 4992
rect 28906 4800 28962 4856
rect 28722 3168 28778 3224
rect 28814 2372 28870 2408
rect 28814 2352 28816 2372
rect 28816 2352 28868 2372
rect 28868 2352 28870 2372
rect 29274 5344 29330 5400
rect 29642 9016 29698 9072
rect 29550 7384 29606 7440
rect 29642 5480 29698 5536
rect 29550 5108 29552 5128
rect 29552 5108 29604 5128
rect 29604 5108 29606 5128
rect 29550 5072 29606 5108
rect 30194 9696 30250 9752
rect 30194 8472 30250 8528
rect 30562 9424 30618 9480
rect 30102 7248 30158 7304
rect 30102 6704 30158 6760
rect 30102 6568 30158 6624
rect 30654 8064 30710 8120
rect 30654 7828 30656 7848
rect 30656 7828 30708 7848
rect 30708 7828 30710 7848
rect 30654 7792 30710 7828
rect 30654 6976 30710 7032
rect 30562 5616 30618 5672
rect 31206 10684 31208 10704
rect 31208 10684 31260 10704
rect 31260 10684 31262 10704
rect 31206 10648 31262 10684
rect 31206 10124 31262 10160
rect 31206 10104 31208 10124
rect 31208 10104 31260 10124
rect 31260 10104 31262 10124
rect 36520 16346 36576 16348
rect 36600 16346 36656 16348
rect 36680 16346 36736 16348
rect 36760 16346 36816 16348
rect 36520 16294 36566 16346
rect 36566 16294 36576 16346
rect 36600 16294 36630 16346
rect 36630 16294 36642 16346
rect 36642 16294 36656 16346
rect 36680 16294 36694 16346
rect 36694 16294 36706 16346
rect 36706 16294 36736 16346
rect 36760 16294 36770 16346
rect 36770 16294 36816 16346
rect 36520 16292 36576 16294
rect 36600 16292 36656 16294
rect 36680 16292 36736 16294
rect 36760 16292 36816 16294
rect 35860 15802 35916 15804
rect 35940 15802 35996 15804
rect 36020 15802 36076 15804
rect 36100 15802 36156 15804
rect 35860 15750 35906 15802
rect 35906 15750 35916 15802
rect 35940 15750 35970 15802
rect 35970 15750 35982 15802
rect 35982 15750 35996 15802
rect 36020 15750 36034 15802
rect 36034 15750 36046 15802
rect 36046 15750 36076 15802
rect 36100 15750 36110 15802
rect 36110 15750 36156 15802
rect 35860 15748 35916 15750
rect 35940 15748 35996 15750
rect 36020 15748 36076 15750
rect 36100 15748 36156 15750
rect 36520 15258 36576 15260
rect 36600 15258 36656 15260
rect 36680 15258 36736 15260
rect 36760 15258 36816 15260
rect 36520 15206 36566 15258
rect 36566 15206 36576 15258
rect 36600 15206 36630 15258
rect 36630 15206 36642 15258
rect 36642 15206 36656 15258
rect 36680 15206 36694 15258
rect 36694 15206 36706 15258
rect 36706 15206 36736 15258
rect 36760 15206 36770 15258
rect 36770 15206 36816 15258
rect 36520 15204 36576 15206
rect 36600 15204 36656 15206
rect 36680 15204 36736 15206
rect 36760 15204 36816 15206
rect 35860 14714 35916 14716
rect 35940 14714 35996 14716
rect 36020 14714 36076 14716
rect 36100 14714 36156 14716
rect 35860 14662 35906 14714
rect 35906 14662 35916 14714
rect 35940 14662 35970 14714
rect 35970 14662 35982 14714
rect 35982 14662 35996 14714
rect 36020 14662 36034 14714
rect 36034 14662 36046 14714
rect 36046 14662 36076 14714
rect 36100 14662 36110 14714
rect 36110 14662 36156 14714
rect 35860 14660 35916 14662
rect 35940 14660 35996 14662
rect 36020 14660 36076 14662
rect 36100 14660 36156 14662
rect 39118 14456 39174 14512
rect 66580 37562 66636 37564
rect 66660 37562 66716 37564
rect 66740 37562 66796 37564
rect 66820 37562 66876 37564
rect 66580 37510 66626 37562
rect 66626 37510 66636 37562
rect 66660 37510 66690 37562
rect 66690 37510 66702 37562
rect 66702 37510 66716 37562
rect 66740 37510 66754 37562
rect 66754 37510 66766 37562
rect 66766 37510 66796 37562
rect 66820 37510 66830 37562
rect 66830 37510 66876 37562
rect 66580 37508 66636 37510
rect 66660 37508 66716 37510
rect 66740 37508 66796 37510
rect 66820 37508 66876 37510
rect 67240 37018 67296 37020
rect 67320 37018 67376 37020
rect 67400 37018 67456 37020
rect 67480 37018 67536 37020
rect 67240 36966 67286 37018
rect 67286 36966 67296 37018
rect 67320 36966 67350 37018
rect 67350 36966 67362 37018
rect 67362 36966 67376 37018
rect 67400 36966 67414 37018
rect 67414 36966 67426 37018
rect 67426 36966 67456 37018
rect 67480 36966 67490 37018
rect 67490 36966 67536 37018
rect 67240 36964 67296 36966
rect 67320 36964 67376 36966
rect 67400 36964 67456 36966
rect 67480 36964 67536 36966
rect 66580 36474 66636 36476
rect 66660 36474 66716 36476
rect 66740 36474 66796 36476
rect 66820 36474 66876 36476
rect 66580 36422 66626 36474
rect 66626 36422 66636 36474
rect 66660 36422 66690 36474
rect 66690 36422 66702 36474
rect 66702 36422 66716 36474
rect 66740 36422 66754 36474
rect 66754 36422 66766 36474
rect 66766 36422 66796 36474
rect 66820 36422 66830 36474
rect 66830 36422 66876 36474
rect 66580 36420 66636 36422
rect 66660 36420 66716 36422
rect 66740 36420 66796 36422
rect 66820 36420 66876 36422
rect 67240 35930 67296 35932
rect 67320 35930 67376 35932
rect 67400 35930 67456 35932
rect 67480 35930 67536 35932
rect 67240 35878 67286 35930
rect 67286 35878 67296 35930
rect 67320 35878 67350 35930
rect 67350 35878 67362 35930
rect 67362 35878 67376 35930
rect 67400 35878 67414 35930
rect 67414 35878 67426 35930
rect 67426 35878 67456 35930
rect 67480 35878 67490 35930
rect 67490 35878 67536 35930
rect 67240 35876 67296 35878
rect 67320 35876 67376 35878
rect 67400 35876 67456 35878
rect 67480 35876 67536 35878
rect 66580 35386 66636 35388
rect 66660 35386 66716 35388
rect 66740 35386 66796 35388
rect 66820 35386 66876 35388
rect 66580 35334 66626 35386
rect 66626 35334 66636 35386
rect 66660 35334 66690 35386
rect 66690 35334 66702 35386
rect 66702 35334 66716 35386
rect 66740 35334 66754 35386
rect 66754 35334 66766 35386
rect 66766 35334 66796 35386
rect 66820 35334 66830 35386
rect 66830 35334 66876 35386
rect 66580 35332 66636 35334
rect 66660 35332 66716 35334
rect 66740 35332 66796 35334
rect 66820 35332 66876 35334
rect 67240 34842 67296 34844
rect 67320 34842 67376 34844
rect 67400 34842 67456 34844
rect 67480 34842 67536 34844
rect 67240 34790 67286 34842
rect 67286 34790 67296 34842
rect 67320 34790 67350 34842
rect 67350 34790 67362 34842
rect 67362 34790 67376 34842
rect 67400 34790 67414 34842
rect 67414 34790 67426 34842
rect 67426 34790 67456 34842
rect 67480 34790 67490 34842
rect 67490 34790 67536 34842
rect 67240 34788 67296 34790
rect 67320 34788 67376 34790
rect 67400 34788 67456 34790
rect 67480 34788 67536 34790
rect 66580 34298 66636 34300
rect 66660 34298 66716 34300
rect 66740 34298 66796 34300
rect 66820 34298 66876 34300
rect 66580 34246 66626 34298
rect 66626 34246 66636 34298
rect 66660 34246 66690 34298
rect 66690 34246 66702 34298
rect 66702 34246 66716 34298
rect 66740 34246 66754 34298
rect 66754 34246 66766 34298
rect 66766 34246 66796 34298
rect 66820 34246 66830 34298
rect 66830 34246 66876 34298
rect 66580 34244 66636 34246
rect 66660 34244 66716 34246
rect 66740 34244 66796 34246
rect 66820 34244 66876 34246
rect 67240 33754 67296 33756
rect 67320 33754 67376 33756
rect 67400 33754 67456 33756
rect 67480 33754 67536 33756
rect 67240 33702 67286 33754
rect 67286 33702 67296 33754
rect 67320 33702 67350 33754
rect 67350 33702 67362 33754
rect 67362 33702 67376 33754
rect 67400 33702 67414 33754
rect 67414 33702 67426 33754
rect 67426 33702 67456 33754
rect 67480 33702 67490 33754
rect 67490 33702 67536 33754
rect 67240 33700 67296 33702
rect 67320 33700 67376 33702
rect 67400 33700 67456 33702
rect 67480 33700 67536 33702
rect 66580 33210 66636 33212
rect 66660 33210 66716 33212
rect 66740 33210 66796 33212
rect 66820 33210 66876 33212
rect 66580 33158 66626 33210
rect 66626 33158 66636 33210
rect 66660 33158 66690 33210
rect 66690 33158 66702 33210
rect 66702 33158 66716 33210
rect 66740 33158 66754 33210
rect 66754 33158 66766 33210
rect 66766 33158 66796 33210
rect 66820 33158 66830 33210
rect 66830 33158 66876 33210
rect 66580 33156 66636 33158
rect 66660 33156 66716 33158
rect 66740 33156 66796 33158
rect 66820 33156 66876 33158
rect 67240 32666 67296 32668
rect 67320 32666 67376 32668
rect 67400 32666 67456 32668
rect 67480 32666 67536 32668
rect 67240 32614 67286 32666
rect 67286 32614 67296 32666
rect 67320 32614 67350 32666
rect 67350 32614 67362 32666
rect 67362 32614 67376 32666
rect 67400 32614 67414 32666
rect 67414 32614 67426 32666
rect 67426 32614 67456 32666
rect 67480 32614 67490 32666
rect 67490 32614 67536 32666
rect 67240 32612 67296 32614
rect 67320 32612 67376 32614
rect 67400 32612 67456 32614
rect 67480 32612 67536 32614
rect 66580 32122 66636 32124
rect 66660 32122 66716 32124
rect 66740 32122 66796 32124
rect 66820 32122 66876 32124
rect 66580 32070 66626 32122
rect 66626 32070 66636 32122
rect 66660 32070 66690 32122
rect 66690 32070 66702 32122
rect 66702 32070 66716 32122
rect 66740 32070 66754 32122
rect 66754 32070 66766 32122
rect 66766 32070 66796 32122
rect 66820 32070 66830 32122
rect 66830 32070 66876 32122
rect 66580 32068 66636 32070
rect 66660 32068 66716 32070
rect 66740 32068 66796 32070
rect 66820 32068 66876 32070
rect 67240 31578 67296 31580
rect 67320 31578 67376 31580
rect 67400 31578 67456 31580
rect 67480 31578 67536 31580
rect 67240 31526 67286 31578
rect 67286 31526 67296 31578
rect 67320 31526 67350 31578
rect 67350 31526 67362 31578
rect 67362 31526 67376 31578
rect 67400 31526 67414 31578
rect 67414 31526 67426 31578
rect 67426 31526 67456 31578
rect 67480 31526 67490 31578
rect 67490 31526 67536 31578
rect 67240 31524 67296 31526
rect 67320 31524 67376 31526
rect 67400 31524 67456 31526
rect 67480 31524 67536 31526
rect 66580 31034 66636 31036
rect 66660 31034 66716 31036
rect 66740 31034 66796 31036
rect 66820 31034 66876 31036
rect 66580 30982 66626 31034
rect 66626 30982 66636 31034
rect 66660 30982 66690 31034
rect 66690 30982 66702 31034
rect 66702 30982 66716 31034
rect 66740 30982 66754 31034
rect 66754 30982 66766 31034
rect 66766 30982 66796 31034
rect 66820 30982 66830 31034
rect 66830 30982 66876 31034
rect 66580 30980 66636 30982
rect 66660 30980 66716 30982
rect 66740 30980 66796 30982
rect 66820 30980 66876 30982
rect 67240 30490 67296 30492
rect 67320 30490 67376 30492
rect 67400 30490 67456 30492
rect 67480 30490 67536 30492
rect 67240 30438 67286 30490
rect 67286 30438 67296 30490
rect 67320 30438 67350 30490
rect 67350 30438 67362 30490
rect 67362 30438 67376 30490
rect 67400 30438 67414 30490
rect 67414 30438 67426 30490
rect 67426 30438 67456 30490
rect 67480 30438 67490 30490
rect 67490 30438 67536 30490
rect 67240 30436 67296 30438
rect 67320 30436 67376 30438
rect 67400 30436 67456 30438
rect 67480 30436 67536 30438
rect 66580 29946 66636 29948
rect 66660 29946 66716 29948
rect 66740 29946 66796 29948
rect 66820 29946 66876 29948
rect 66580 29894 66626 29946
rect 66626 29894 66636 29946
rect 66660 29894 66690 29946
rect 66690 29894 66702 29946
rect 66702 29894 66716 29946
rect 66740 29894 66754 29946
rect 66754 29894 66766 29946
rect 66766 29894 66796 29946
rect 66820 29894 66830 29946
rect 66830 29894 66876 29946
rect 66580 29892 66636 29894
rect 66660 29892 66716 29894
rect 66740 29892 66796 29894
rect 66820 29892 66876 29894
rect 67240 29402 67296 29404
rect 67320 29402 67376 29404
rect 67400 29402 67456 29404
rect 67480 29402 67536 29404
rect 67240 29350 67286 29402
rect 67286 29350 67296 29402
rect 67320 29350 67350 29402
rect 67350 29350 67362 29402
rect 67362 29350 67376 29402
rect 67400 29350 67414 29402
rect 67414 29350 67426 29402
rect 67426 29350 67456 29402
rect 67480 29350 67490 29402
rect 67490 29350 67536 29402
rect 67240 29348 67296 29350
rect 67320 29348 67376 29350
rect 67400 29348 67456 29350
rect 67480 29348 67536 29350
rect 66580 28858 66636 28860
rect 66660 28858 66716 28860
rect 66740 28858 66796 28860
rect 66820 28858 66876 28860
rect 66580 28806 66626 28858
rect 66626 28806 66636 28858
rect 66660 28806 66690 28858
rect 66690 28806 66702 28858
rect 66702 28806 66716 28858
rect 66740 28806 66754 28858
rect 66754 28806 66766 28858
rect 66766 28806 66796 28858
rect 66820 28806 66830 28858
rect 66830 28806 66876 28858
rect 66580 28804 66636 28806
rect 66660 28804 66716 28806
rect 66740 28804 66796 28806
rect 66820 28804 66876 28806
rect 67240 28314 67296 28316
rect 67320 28314 67376 28316
rect 67400 28314 67456 28316
rect 67480 28314 67536 28316
rect 67240 28262 67286 28314
rect 67286 28262 67296 28314
rect 67320 28262 67350 28314
rect 67350 28262 67362 28314
rect 67362 28262 67376 28314
rect 67400 28262 67414 28314
rect 67414 28262 67426 28314
rect 67426 28262 67456 28314
rect 67480 28262 67490 28314
rect 67490 28262 67536 28314
rect 67240 28260 67296 28262
rect 67320 28260 67376 28262
rect 67400 28260 67456 28262
rect 67480 28260 67536 28262
rect 66580 27770 66636 27772
rect 66660 27770 66716 27772
rect 66740 27770 66796 27772
rect 66820 27770 66876 27772
rect 66580 27718 66626 27770
rect 66626 27718 66636 27770
rect 66660 27718 66690 27770
rect 66690 27718 66702 27770
rect 66702 27718 66716 27770
rect 66740 27718 66754 27770
rect 66754 27718 66766 27770
rect 66766 27718 66796 27770
rect 66820 27718 66830 27770
rect 66830 27718 66876 27770
rect 66580 27716 66636 27718
rect 66660 27716 66716 27718
rect 66740 27716 66796 27718
rect 66820 27716 66876 27718
rect 67240 27226 67296 27228
rect 67320 27226 67376 27228
rect 67400 27226 67456 27228
rect 67480 27226 67536 27228
rect 67240 27174 67286 27226
rect 67286 27174 67296 27226
rect 67320 27174 67350 27226
rect 67350 27174 67362 27226
rect 67362 27174 67376 27226
rect 67400 27174 67414 27226
rect 67414 27174 67426 27226
rect 67426 27174 67456 27226
rect 67480 27174 67490 27226
rect 67490 27174 67536 27226
rect 67240 27172 67296 27174
rect 67320 27172 67376 27174
rect 67400 27172 67456 27174
rect 67480 27172 67536 27174
rect 66580 26682 66636 26684
rect 66660 26682 66716 26684
rect 66740 26682 66796 26684
rect 66820 26682 66876 26684
rect 66580 26630 66626 26682
rect 66626 26630 66636 26682
rect 66660 26630 66690 26682
rect 66690 26630 66702 26682
rect 66702 26630 66716 26682
rect 66740 26630 66754 26682
rect 66754 26630 66766 26682
rect 66766 26630 66796 26682
rect 66820 26630 66830 26682
rect 66830 26630 66876 26682
rect 66580 26628 66636 26630
rect 66660 26628 66716 26630
rect 66740 26628 66796 26630
rect 66820 26628 66876 26630
rect 67240 26138 67296 26140
rect 67320 26138 67376 26140
rect 67400 26138 67456 26140
rect 67480 26138 67536 26140
rect 67240 26086 67286 26138
rect 67286 26086 67296 26138
rect 67320 26086 67350 26138
rect 67350 26086 67362 26138
rect 67362 26086 67376 26138
rect 67400 26086 67414 26138
rect 67414 26086 67426 26138
rect 67426 26086 67456 26138
rect 67480 26086 67490 26138
rect 67490 26086 67536 26138
rect 67240 26084 67296 26086
rect 67320 26084 67376 26086
rect 67400 26084 67456 26086
rect 67480 26084 67536 26086
rect 66580 25594 66636 25596
rect 66660 25594 66716 25596
rect 66740 25594 66796 25596
rect 66820 25594 66876 25596
rect 66580 25542 66626 25594
rect 66626 25542 66636 25594
rect 66660 25542 66690 25594
rect 66690 25542 66702 25594
rect 66702 25542 66716 25594
rect 66740 25542 66754 25594
rect 66754 25542 66766 25594
rect 66766 25542 66796 25594
rect 66820 25542 66830 25594
rect 66830 25542 66876 25594
rect 66580 25540 66636 25542
rect 66660 25540 66716 25542
rect 66740 25540 66796 25542
rect 66820 25540 66876 25542
rect 67240 25050 67296 25052
rect 67320 25050 67376 25052
rect 67400 25050 67456 25052
rect 67480 25050 67536 25052
rect 67240 24998 67286 25050
rect 67286 24998 67296 25050
rect 67320 24998 67350 25050
rect 67350 24998 67362 25050
rect 67362 24998 67376 25050
rect 67400 24998 67414 25050
rect 67414 24998 67426 25050
rect 67426 24998 67456 25050
rect 67480 24998 67490 25050
rect 67490 24998 67536 25050
rect 67240 24996 67296 24998
rect 67320 24996 67376 24998
rect 67400 24996 67456 24998
rect 67480 24996 67536 24998
rect 66580 24506 66636 24508
rect 66660 24506 66716 24508
rect 66740 24506 66796 24508
rect 66820 24506 66876 24508
rect 66580 24454 66626 24506
rect 66626 24454 66636 24506
rect 66660 24454 66690 24506
rect 66690 24454 66702 24506
rect 66702 24454 66716 24506
rect 66740 24454 66754 24506
rect 66754 24454 66766 24506
rect 66766 24454 66796 24506
rect 66820 24454 66830 24506
rect 66830 24454 66876 24506
rect 66580 24452 66636 24454
rect 66660 24452 66716 24454
rect 66740 24452 66796 24454
rect 66820 24452 66876 24454
rect 67240 23962 67296 23964
rect 67320 23962 67376 23964
rect 67400 23962 67456 23964
rect 67480 23962 67536 23964
rect 67240 23910 67286 23962
rect 67286 23910 67296 23962
rect 67320 23910 67350 23962
rect 67350 23910 67362 23962
rect 67362 23910 67376 23962
rect 67400 23910 67414 23962
rect 67414 23910 67426 23962
rect 67426 23910 67456 23962
rect 67480 23910 67490 23962
rect 67490 23910 67536 23962
rect 67240 23908 67296 23910
rect 67320 23908 67376 23910
rect 67400 23908 67456 23910
rect 67480 23908 67536 23910
rect 66580 23418 66636 23420
rect 66660 23418 66716 23420
rect 66740 23418 66796 23420
rect 66820 23418 66876 23420
rect 66580 23366 66626 23418
rect 66626 23366 66636 23418
rect 66660 23366 66690 23418
rect 66690 23366 66702 23418
rect 66702 23366 66716 23418
rect 66740 23366 66754 23418
rect 66754 23366 66766 23418
rect 66766 23366 66796 23418
rect 66820 23366 66830 23418
rect 66830 23366 66876 23418
rect 66580 23364 66636 23366
rect 66660 23364 66716 23366
rect 66740 23364 66796 23366
rect 66820 23364 66876 23366
rect 67240 22874 67296 22876
rect 67320 22874 67376 22876
rect 67400 22874 67456 22876
rect 67480 22874 67536 22876
rect 67240 22822 67286 22874
rect 67286 22822 67296 22874
rect 67320 22822 67350 22874
rect 67350 22822 67362 22874
rect 67362 22822 67376 22874
rect 67400 22822 67414 22874
rect 67414 22822 67426 22874
rect 67426 22822 67456 22874
rect 67480 22822 67490 22874
rect 67490 22822 67536 22874
rect 67240 22820 67296 22822
rect 67320 22820 67376 22822
rect 67400 22820 67456 22822
rect 67480 22820 67536 22822
rect 66580 22330 66636 22332
rect 66660 22330 66716 22332
rect 66740 22330 66796 22332
rect 66820 22330 66876 22332
rect 66580 22278 66626 22330
rect 66626 22278 66636 22330
rect 66660 22278 66690 22330
rect 66690 22278 66702 22330
rect 66702 22278 66716 22330
rect 66740 22278 66754 22330
rect 66754 22278 66766 22330
rect 66766 22278 66796 22330
rect 66820 22278 66830 22330
rect 66830 22278 66876 22330
rect 66580 22276 66636 22278
rect 66660 22276 66716 22278
rect 66740 22276 66796 22278
rect 66820 22276 66876 22278
rect 67240 21786 67296 21788
rect 67320 21786 67376 21788
rect 67400 21786 67456 21788
rect 67480 21786 67536 21788
rect 67240 21734 67286 21786
rect 67286 21734 67296 21786
rect 67320 21734 67350 21786
rect 67350 21734 67362 21786
rect 67362 21734 67376 21786
rect 67400 21734 67414 21786
rect 67414 21734 67426 21786
rect 67426 21734 67456 21786
rect 67480 21734 67490 21786
rect 67490 21734 67536 21786
rect 67240 21732 67296 21734
rect 67320 21732 67376 21734
rect 67400 21732 67456 21734
rect 67480 21732 67536 21734
rect 66580 21242 66636 21244
rect 66660 21242 66716 21244
rect 66740 21242 66796 21244
rect 66820 21242 66876 21244
rect 66580 21190 66626 21242
rect 66626 21190 66636 21242
rect 66660 21190 66690 21242
rect 66690 21190 66702 21242
rect 66702 21190 66716 21242
rect 66740 21190 66754 21242
rect 66754 21190 66766 21242
rect 66766 21190 66796 21242
rect 66820 21190 66830 21242
rect 66830 21190 66876 21242
rect 66580 21188 66636 21190
rect 66660 21188 66716 21190
rect 66740 21188 66796 21190
rect 66820 21188 66876 21190
rect 67240 20698 67296 20700
rect 67320 20698 67376 20700
rect 67400 20698 67456 20700
rect 67480 20698 67536 20700
rect 67240 20646 67286 20698
rect 67286 20646 67296 20698
rect 67320 20646 67350 20698
rect 67350 20646 67362 20698
rect 67362 20646 67376 20698
rect 67400 20646 67414 20698
rect 67414 20646 67426 20698
rect 67426 20646 67456 20698
rect 67480 20646 67490 20698
rect 67490 20646 67536 20698
rect 67240 20644 67296 20646
rect 67320 20644 67376 20646
rect 67400 20644 67456 20646
rect 67480 20644 67536 20646
rect 66580 20154 66636 20156
rect 66660 20154 66716 20156
rect 66740 20154 66796 20156
rect 66820 20154 66876 20156
rect 66580 20102 66626 20154
rect 66626 20102 66636 20154
rect 66660 20102 66690 20154
rect 66690 20102 66702 20154
rect 66702 20102 66716 20154
rect 66740 20102 66754 20154
rect 66754 20102 66766 20154
rect 66766 20102 66796 20154
rect 66820 20102 66830 20154
rect 66830 20102 66876 20154
rect 66580 20100 66636 20102
rect 66660 20100 66716 20102
rect 66740 20100 66796 20102
rect 66820 20100 66876 20102
rect 67240 19610 67296 19612
rect 67320 19610 67376 19612
rect 67400 19610 67456 19612
rect 67480 19610 67536 19612
rect 67240 19558 67286 19610
rect 67286 19558 67296 19610
rect 67320 19558 67350 19610
rect 67350 19558 67362 19610
rect 67362 19558 67376 19610
rect 67400 19558 67414 19610
rect 67414 19558 67426 19610
rect 67426 19558 67456 19610
rect 67480 19558 67490 19610
rect 67490 19558 67536 19610
rect 67240 19556 67296 19558
rect 67320 19556 67376 19558
rect 67400 19556 67456 19558
rect 67480 19556 67536 19558
rect 66580 19066 66636 19068
rect 66660 19066 66716 19068
rect 66740 19066 66796 19068
rect 66820 19066 66876 19068
rect 66580 19014 66626 19066
rect 66626 19014 66636 19066
rect 66660 19014 66690 19066
rect 66690 19014 66702 19066
rect 66702 19014 66716 19066
rect 66740 19014 66754 19066
rect 66754 19014 66766 19066
rect 66766 19014 66796 19066
rect 66820 19014 66830 19066
rect 66830 19014 66876 19066
rect 66580 19012 66636 19014
rect 66660 19012 66716 19014
rect 66740 19012 66796 19014
rect 66820 19012 66876 19014
rect 67240 18522 67296 18524
rect 67320 18522 67376 18524
rect 67400 18522 67456 18524
rect 67480 18522 67536 18524
rect 67240 18470 67286 18522
rect 67286 18470 67296 18522
rect 67320 18470 67350 18522
rect 67350 18470 67362 18522
rect 67362 18470 67376 18522
rect 67400 18470 67414 18522
rect 67414 18470 67426 18522
rect 67426 18470 67456 18522
rect 67480 18470 67490 18522
rect 67490 18470 67536 18522
rect 67240 18468 67296 18470
rect 67320 18468 67376 18470
rect 67400 18468 67456 18470
rect 67480 18468 67536 18470
rect 66580 17978 66636 17980
rect 66660 17978 66716 17980
rect 66740 17978 66796 17980
rect 66820 17978 66876 17980
rect 66580 17926 66626 17978
rect 66626 17926 66636 17978
rect 66660 17926 66690 17978
rect 66690 17926 66702 17978
rect 66702 17926 66716 17978
rect 66740 17926 66754 17978
rect 66754 17926 66766 17978
rect 66766 17926 66796 17978
rect 66820 17926 66830 17978
rect 66830 17926 66876 17978
rect 66580 17924 66636 17926
rect 66660 17924 66716 17926
rect 66740 17924 66796 17926
rect 66820 17924 66876 17926
rect 67240 17434 67296 17436
rect 67320 17434 67376 17436
rect 67400 17434 67456 17436
rect 67480 17434 67536 17436
rect 67240 17382 67286 17434
rect 67286 17382 67296 17434
rect 67320 17382 67350 17434
rect 67350 17382 67362 17434
rect 67362 17382 67376 17434
rect 67400 17382 67414 17434
rect 67414 17382 67426 17434
rect 67426 17382 67456 17434
rect 67480 17382 67490 17434
rect 67490 17382 67536 17434
rect 67240 17380 67296 17382
rect 67320 17380 67376 17382
rect 67400 17380 67456 17382
rect 67480 17380 67536 17382
rect 66580 16890 66636 16892
rect 66660 16890 66716 16892
rect 66740 16890 66796 16892
rect 66820 16890 66876 16892
rect 66580 16838 66626 16890
rect 66626 16838 66636 16890
rect 66660 16838 66690 16890
rect 66690 16838 66702 16890
rect 66702 16838 66716 16890
rect 66740 16838 66754 16890
rect 66754 16838 66766 16890
rect 66766 16838 66796 16890
rect 66820 16838 66830 16890
rect 66830 16838 66876 16890
rect 66580 16836 66636 16838
rect 66660 16836 66716 16838
rect 66740 16836 66796 16838
rect 66820 16836 66876 16838
rect 67240 16346 67296 16348
rect 67320 16346 67376 16348
rect 67400 16346 67456 16348
rect 67480 16346 67536 16348
rect 67240 16294 67286 16346
rect 67286 16294 67296 16346
rect 67320 16294 67350 16346
rect 67350 16294 67362 16346
rect 67362 16294 67376 16346
rect 67400 16294 67414 16346
rect 67414 16294 67426 16346
rect 67426 16294 67456 16346
rect 67480 16294 67490 16346
rect 67490 16294 67536 16346
rect 67240 16292 67296 16294
rect 67320 16292 67376 16294
rect 67400 16292 67456 16294
rect 67480 16292 67536 16294
rect 66580 15802 66636 15804
rect 66660 15802 66716 15804
rect 66740 15802 66796 15804
rect 66820 15802 66876 15804
rect 66580 15750 66626 15802
rect 66626 15750 66636 15802
rect 66660 15750 66690 15802
rect 66690 15750 66702 15802
rect 66702 15750 66716 15802
rect 66740 15750 66754 15802
rect 66754 15750 66766 15802
rect 66766 15750 66796 15802
rect 66820 15750 66830 15802
rect 66830 15750 66876 15802
rect 66580 15748 66636 15750
rect 66660 15748 66716 15750
rect 66740 15748 66796 15750
rect 66820 15748 66876 15750
rect 67240 15258 67296 15260
rect 67320 15258 67376 15260
rect 67400 15258 67456 15260
rect 67480 15258 67536 15260
rect 67240 15206 67286 15258
rect 67286 15206 67296 15258
rect 67320 15206 67350 15258
rect 67350 15206 67362 15258
rect 67362 15206 67376 15258
rect 67400 15206 67414 15258
rect 67414 15206 67426 15258
rect 67426 15206 67456 15258
rect 67480 15206 67490 15258
rect 67490 15206 67536 15258
rect 67240 15204 67296 15206
rect 67320 15204 67376 15206
rect 67400 15204 67456 15206
rect 67480 15204 67536 15206
rect 66580 14714 66636 14716
rect 66660 14714 66716 14716
rect 66740 14714 66796 14716
rect 66820 14714 66876 14716
rect 66580 14662 66626 14714
rect 66626 14662 66636 14714
rect 66660 14662 66690 14714
rect 66690 14662 66702 14714
rect 66702 14662 66716 14714
rect 66740 14662 66754 14714
rect 66754 14662 66766 14714
rect 66766 14662 66796 14714
rect 66820 14662 66830 14714
rect 66830 14662 66876 14714
rect 66580 14660 66636 14662
rect 66660 14660 66716 14662
rect 66740 14660 66796 14662
rect 66820 14660 66876 14662
rect 36520 14170 36576 14172
rect 36600 14170 36656 14172
rect 36680 14170 36736 14172
rect 36760 14170 36816 14172
rect 36520 14118 36566 14170
rect 36566 14118 36576 14170
rect 36600 14118 36630 14170
rect 36630 14118 36642 14170
rect 36642 14118 36656 14170
rect 36680 14118 36694 14170
rect 36694 14118 36706 14170
rect 36706 14118 36736 14170
rect 36760 14118 36770 14170
rect 36770 14118 36816 14170
rect 36520 14116 36576 14118
rect 36600 14116 36656 14118
rect 36680 14116 36736 14118
rect 36760 14116 36816 14118
rect 67240 14170 67296 14172
rect 67320 14170 67376 14172
rect 67400 14170 67456 14172
rect 67480 14170 67536 14172
rect 67240 14118 67286 14170
rect 67286 14118 67296 14170
rect 67320 14118 67350 14170
rect 67350 14118 67362 14170
rect 67362 14118 67376 14170
rect 67400 14118 67414 14170
rect 67414 14118 67426 14170
rect 67426 14118 67456 14170
rect 67480 14118 67490 14170
rect 67490 14118 67536 14170
rect 67240 14116 67296 14118
rect 67320 14116 67376 14118
rect 67400 14116 67456 14118
rect 67480 14116 67536 14118
rect 35860 13626 35916 13628
rect 35940 13626 35996 13628
rect 36020 13626 36076 13628
rect 36100 13626 36156 13628
rect 35860 13574 35906 13626
rect 35906 13574 35916 13626
rect 35940 13574 35970 13626
rect 35970 13574 35982 13626
rect 35982 13574 35996 13626
rect 36020 13574 36034 13626
rect 36034 13574 36046 13626
rect 36046 13574 36076 13626
rect 36100 13574 36110 13626
rect 36110 13574 36156 13626
rect 35860 13572 35916 13574
rect 35940 13572 35996 13574
rect 36020 13572 36076 13574
rect 36100 13572 36156 13574
rect 66580 13626 66636 13628
rect 66660 13626 66716 13628
rect 66740 13626 66796 13628
rect 66820 13626 66876 13628
rect 66580 13574 66626 13626
rect 66626 13574 66636 13626
rect 66660 13574 66690 13626
rect 66690 13574 66702 13626
rect 66702 13574 66716 13626
rect 66740 13574 66754 13626
rect 66754 13574 66766 13626
rect 66766 13574 66796 13626
rect 66820 13574 66830 13626
rect 66830 13574 66876 13626
rect 66580 13572 66636 13574
rect 66660 13572 66716 13574
rect 66740 13572 66796 13574
rect 66820 13572 66876 13574
rect 36520 13082 36576 13084
rect 36600 13082 36656 13084
rect 36680 13082 36736 13084
rect 36760 13082 36816 13084
rect 36520 13030 36566 13082
rect 36566 13030 36576 13082
rect 36600 13030 36630 13082
rect 36630 13030 36642 13082
rect 36642 13030 36656 13082
rect 36680 13030 36694 13082
rect 36694 13030 36706 13082
rect 36706 13030 36736 13082
rect 36760 13030 36770 13082
rect 36770 13030 36816 13082
rect 36520 13028 36576 13030
rect 36600 13028 36656 13030
rect 36680 13028 36736 13030
rect 36760 13028 36816 13030
rect 67240 13082 67296 13084
rect 67320 13082 67376 13084
rect 67400 13082 67456 13084
rect 67480 13082 67536 13084
rect 67240 13030 67286 13082
rect 67286 13030 67296 13082
rect 67320 13030 67350 13082
rect 67350 13030 67362 13082
rect 67362 13030 67376 13082
rect 67400 13030 67414 13082
rect 67414 13030 67426 13082
rect 67426 13030 67456 13082
rect 67480 13030 67490 13082
rect 67490 13030 67536 13082
rect 67240 13028 67296 13030
rect 67320 13028 67376 13030
rect 67400 13028 67456 13030
rect 67480 13028 67536 13030
rect 35860 12538 35916 12540
rect 35940 12538 35996 12540
rect 36020 12538 36076 12540
rect 36100 12538 36156 12540
rect 35860 12486 35906 12538
rect 35906 12486 35916 12538
rect 35940 12486 35970 12538
rect 35970 12486 35982 12538
rect 35982 12486 35996 12538
rect 36020 12486 36034 12538
rect 36034 12486 36046 12538
rect 36046 12486 36076 12538
rect 36100 12486 36110 12538
rect 36110 12486 36156 12538
rect 35860 12484 35916 12486
rect 35940 12484 35996 12486
rect 36020 12484 36076 12486
rect 36100 12484 36156 12486
rect 36520 11994 36576 11996
rect 36600 11994 36656 11996
rect 36680 11994 36736 11996
rect 36760 11994 36816 11996
rect 36520 11942 36566 11994
rect 36566 11942 36576 11994
rect 36600 11942 36630 11994
rect 36630 11942 36642 11994
rect 36642 11942 36656 11994
rect 36680 11942 36694 11994
rect 36694 11942 36706 11994
rect 36706 11942 36736 11994
rect 36760 11942 36770 11994
rect 36770 11942 36816 11994
rect 36520 11940 36576 11942
rect 36600 11940 36656 11942
rect 36680 11940 36736 11942
rect 36760 11940 36816 11942
rect 35860 11450 35916 11452
rect 35940 11450 35996 11452
rect 36020 11450 36076 11452
rect 36100 11450 36156 11452
rect 35860 11398 35906 11450
rect 35906 11398 35916 11450
rect 35940 11398 35970 11450
rect 35970 11398 35982 11450
rect 35982 11398 35996 11450
rect 36020 11398 36034 11450
rect 36034 11398 36046 11450
rect 36046 11398 36076 11450
rect 36100 11398 36110 11450
rect 36110 11398 36156 11450
rect 35860 11396 35916 11398
rect 35940 11396 35996 11398
rect 36020 11396 36076 11398
rect 36100 11396 36156 11398
rect 31850 10104 31906 10160
rect 31850 9560 31906 9616
rect 31114 6840 31170 6896
rect 30930 6432 30986 6488
rect 30930 6160 30986 6216
rect 30838 4800 30894 4856
rect 30838 4256 30894 4312
rect 31206 6160 31262 6216
rect 31206 5344 31262 5400
rect 31390 8336 31446 8392
rect 31390 8064 31446 8120
rect 31482 7928 31538 7984
rect 31758 8336 31814 8392
rect 31666 7928 31722 7984
rect 31758 7828 31760 7848
rect 31760 7828 31812 7848
rect 31812 7828 31814 7848
rect 31758 7792 31814 7828
rect 31666 7656 31722 7712
rect 31942 7384 31998 7440
rect 31850 6976 31906 7032
rect 31666 6160 31722 6216
rect 31666 5752 31722 5808
rect 31574 5208 31630 5264
rect 31850 5480 31906 5536
rect 32218 8608 32274 8664
rect 32402 8200 32458 8256
rect 32310 7792 32366 7848
rect 32310 7692 32312 7712
rect 32312 7692 32364 7712
rect 32364 7692 32366 7712
rect 32310 7656 32366 7692
rect 32218 7268 32274 7304
rect 32218 7248 32220 7268
rect 32220 7248 32272 7268
rect 32272 7248 32274 7268
rect 32310 6976 32366 7032
rect 32126 6024 32182 6080
rect 32218 5888 32274 5944
rect 32126 5616 32182 5672
rect 32218 5208 32274 5264
rect 32402 6432 32458 6488
rect 32126 4800 32182 4856
rect 32402 4936 32458 4992
rect 31758 3168 31814 3224
rect 33046 9580 33102 9616
rect 33046 9560 33048 9580
rect 33048 9560 33100 9580
rect 33100 9560 33102 9580
rect 33230 9424 33286 9480
rect 33046 8744 33102 8800
rect 33138 8608 33194 8664
rect 33138 8064 33194 8120
rect 33322 8336 33378 8392
rect 33046 6160 33102 6216
rect 33322 6568 33378 6624
rect 32862 3440 32918 3496
rect 33046 3848 33102 3904
rect 33322 4528 33378 4584
rect 33046 2916 33102 2952
rect 33046 2896 33048 2916
rect 33048 2896 33100 2916
rect 33100 2896 33102 2916
rect 33506 4392 33562 4448
rect 33690 9288 33746 9344
rect 33874 8064 33930 8120
rect 33782 7520 33838 7576
rect 33782 6432 33838 6488
rect 34334 6568 34390 6624
rect 33966 5616 34022 5672
rect 34150 5616 34206 5672
rect 34058 3576 34114 3632
rect 33782 3440 33838 3496
rect 33782 3304 33838 3360
rect 33874 3168 33930 3224
rect 34242 5344 34298 5400
rect 34334 3576 34390 3632
rect 34702 8200 34758 8256
rect 34610 5228 34666 5264
rect 34610 5208 34612 5228
rect 34612 5208 34664 5228
rect 34664 5208 34666 5228
rect 34886 6840 34942 6896
rect 35254 8472 35310 8528
rect 35162 6740 35164 6760
rect 35164 6740 35216 6760
rect 35216 6740 35218 6760
rect 35162 6704 35218 6740
rect 35162 6160 35218 6216
rect 35254 4256 35310 4312
rect 35162 3304 35218 3360
rect 35860 10362 35916 10364
rect 35940 10362 35996 10364
rect 36020 10362 36076 10364
rect 36100 10362 36156 10364
rect 35860 10310 35906 10362
rect 35906 10310 35916 10362
rect 35940 10310 35970 10362
rect 35970 10310 35982 10362
rect 35982 10310 35996 10362
rect 36020 10310 36034 10362
rect 36034 10310 36046 10362
rect 36046 10310 36076 10362
rect 36100 10310 36110 10362
rect 36110 10310 36156 10362
rect 35860 10308 35916 10310
rect 35940 10308 35996 10310
rect 36020 10308 36076 10310
rect 36100 10308 36156 10310
rect 36520 10906 36576 10908
rect 36600 10906 36656 10908
rect 36680 10906 36736 10908
rect 36760 10906 36816 10908
rect 36520 10854 36566 10906
rect 36566 10854 36576 10906
rect 36600 10854 36630 10906
rect 36630 10854 36642 10906
rect 36642 10854 36656 10906
rect 36680 10854 36694 10906
rect 36694 10854 36706 10906
rect 36706 10854 36736 10906
rect 36760 10854 36770 10906
rect 36770 10854 36816 10906
rect 36520 10852 36576 10854
rect 36600 10852 36656 10854
rect 36680 10852 36736 10854
rect 36760 10852 36816 10854
rect 36520 9818 36576 9820
rect 36600 9818 36656 9820
rect 36680 9818 36736 9820
rect 36760 9818 36816 9820
rect 36520 9766 36566 9818
rect 36566 9766 36576 9818
rect 36600 9766 36630 9818
rect 36630 9766 36642 9818
rect 36642 9766 36656 9818
rect 36680 9766 36694 9818
rect 36694 9766 36706 9818
rect 36706 9766 36736 9818
rect 36760 9766 36770 9818
rect 36770 9766 36816 9818
rect 36520 9764 36576 9766
rect 36600 9764 36656 9766
rect 36680 9764 36736 9766
rect 36760 9764 36816 9766
rect 35714 9424 35770 9480
rect 35860 9274 35916 9276
rect 35940 9274 35996 9276
rect 36020 9274 36076 9276
rect 36100 9274 36156 9276
rect 35860 9222 35906 9274
rect 35906 9222 35916 9274
rect 35940 9222 35970 9274
rect 35970 9222 35982 9274
rect 35982 9222 35996 9274
rect 36020 9222 36034 9274
rect 36034 9222 36046 9274
rect 36046 9222 36076 9274
rect 36100 9222 36110 9274
rect 36110 9222 36156 9274
rect 35860 9220 35916 9222
rect 35940 9220 35996 9222
rect 36020 9220 36076 9222
rect 36100 9220 36156 9222
rect 35860 8186 35916 8188
rect 35940 8186 35996 8188
rect 36020 8186 36076 8188
rect 36100 8186 36156 8188
rect 35860 8134 35906 8186
rect 35906 8134 35916 8186
rect 35940 8134 35970 8186
rect 35970 8134 35982 8186
rect 35982 8134 35996 8186
rect 36020 8134 36034 8186
rect 36034 8134 36046 8186
rect 36046 8134 36076 8186
rect 36100 8134 36110 8186
rect 36110 8134 36156 8186
rect 35860 8132 35916 8134
rect 35940 8132 35996 8134
rect 36020 8132 36076 8134
rect 36100 8132 36156 8134
rect 36266 7656 36322 7712
rect 35990 7520 36046 7576
rect 35860 7098 35916 7100
rect 35940 7098 35996 7100
rect 36020 7098 36076 7100
rect 36100 7098 36156 7100
rect 35860 7046 35906 7098
rect 35906 7046 35916 7098
rect 35940 7046 35970 7098
rect 35970 7046 35982 7098
rect 35982 7046 35996 7098
rect 36020 7046 36034 7098
rect 36034 7046 36046 7098
rect 36046 7046 36076 7098
rect 36100 7046 36110 7098
rect 36110 7046 36156 7098
rect 35860 7044 35916 7046
rect 35940 7044 35996 7046
rect 36020 7044 36076 7046
rect 36100 7044 36156 7046
rect 35806 6740 35808 6760
rect 35808 6740 35860 6760
rect 35860 6740 35862 6760
rect 36520 8730 36576 8732
rect 36600 8730 36656 8732
rect 36680 8730 36736 8732
rect 36760 8730 36816 8732
rect 36520 8678 36566 8730
rect 36566 8678 36576 8730
rect 36600 8678 36630 8730
rect 36630 8678 36642 8730
rect 36642 8678 36656 8730
rect 36680 8678 36694 8730
rect 36694 8678 36706 8730
rect 36706 8678 36736 8730
rect 36760 8678 36770 8730
rect 36770 8678 36816 8730
rect 36520 8676 36576 8678
rect 36600 8676 36656 8678
rect 36680 8676 36736 8678
rect 36760 8676 36816 8678
rect 36520 7642 36576 7644
rect 36600 7642 36656 7644
rect 36680 7642 36736 7644
rect 36760 7642 36816 7644
rect 36520 7590 36566 7642
rect 36566 7590 36576 7642
rect 36600 7590 36630 7642
rect 36630 7590 36642 7642
rect 36642 7590 36656 7642
rect 36680 7590 36694 7642
rect 36694 7590 36706 7642
rect 36706 7590 36736 7642
rect 36760 7590 36770 7642
rect 36770 7590 36816 7642
rect 36520 7588 36576 7590
rect 36600 7588 36656 7590
rect 36680 7588 36736 7590
rect 36760 7588 36816 7590
rect 35806 6704 35862 6740
rect 35898 6604 35900 6624
rect 35900 6604 35952 6624
rect 35952 6604 35954 6624
rect 35898 6568 35954 6604
rect 36520 6554 36576 6556
rect 36600 6554 36656 6556
rect 36680 6554 36736 6556
rect 36760 6554 36816 6556
rect 36520 6502 36566 6554
rect 36566 6502 36576 6554
rect 36600 6502 36630 6554
rect 36630 6502 36642 6554
rect 36642 6502 36656 6554
rect 36680 6502 36694 6554
rect 36694 6502 36706 6554
rect 36706 6502 36736 6554
rect 36760 6502 36770 6554
rect 36770 6502 36816 6554
rect 36520 6500 36576 6502
rect 36600 6500 36656 6502
rect 36680 6500 36736 6502
rect 36760 6500 36816 6502
rect 35714 6024 35770 6080
rect 35860 6010 35916 6012
rect 35940 6010 35996 6012
rect 36020 6010 36076 6012
rect 36100 6010 36156 6012
rect 35860 5958 35906 6010
rect 35906 5958 35916 6010
rect 35940 5958 35970 6010
rect 35970 5958 35982 6010
rect 35982 5958 35996 6010
rect 36020 5958 36034 6010
rect 36034 5958 36046 6010
rect 36046 5958 36076 6010
rect 36100 5958 36110 6010
rect 36110 5958 36156 6010
rect 35860 5956 35916 5958
rect 35940 5956 35996 5958
rect 36020 5956 36076 5958
rect 36100 5956 36156 5958
rect 35860 4922 35916 4924
rect 35940 4922 35996 4924
rect 36020 4922 36076 4924
rect 36100 4922 36156 4924
rect 35860 4870 35906 4922
rect 35906 4870 35916 4922
rect 35940 4870 35970 4922
rect 35970 4870 35982 4922
rect 35982 4870 35996 4922
rect 36020 4870 36034 4922
rect 36034 4870 36046 4922
rect 36046 4870 36076 4922
rect 36100 4870 36110 4922
rect 36110 4870 36156 4922
rect 35860 4868 35916 4870
rect 35940 4868 35996 4870
rect 36020 4868 36076 4870
rect 36100 4868 36156 4870
rect 35714 4120 35770 4176
rect 35860 3834 35916 3836
rect 35940 3834 35996 3836
rect 36020 3834 36076 3836
rect 36100 3834 36156 3836
rect 35860 3782 35906 3834
rect 35906 3782 35916 3834
rect 35940 3782 35970 3834
rect 35970 3782 35982 3834
rect 35982 3782 35996 3834
rect 36020 3782 36034 3834
rect 36034 3782 36046 3834
rect 36046 3782 36076 3834
rect 36100 3782 36110 3834
rect 36110 3782 36156 3834
rect 35860 3780 35916 3782
rect 35940 3780 35996 3782
rect 36020 3780 36076 3782
rect 36100 3780 36156 3782
rect 36266 2760 36322 2816
rect 35860 2746 35916 2748
rect 35940 2746 35996 2748
rect 36020 2746 36076 2748
rect 36100 2746 36156 2748
rect 35860 2694 35906 2746
rect 35906 2694 35916 2746
rect 35940 2694 35970 2746
rect 35970 2694 35982 2746
rect 35982 2694 35996 2746
rect 36020 2694 36034 2746
rect 36034 2694 36046 2746
rect 36046 2694 36076 2746
rect 36100 2694 36110 2746
rect 36110 2694 36156 2746
rect 35860 2692 35916 2694
rect 35940 2692 35996 2694
rect 36020 2692 36076 2694
rect 36100 2692 36156 2694
rect 36082 1400 36138 1456
rect 36450 5908 36506 5944
rect 36450 5888 36452 5908
rect 36452 5888 36504 5908
rect 36504 5888 36506 5908
rect 36520 5466 36576 5468
rect 36600 5466 36656 5468
rect 36680 5466 36736 5468
rect 36760 5466 36816 5468
rect 36520 5414 36566 5466
rect 36566 5414 36576 5466
rect 36600 5414 36630 5466
rect 36630 5414 36642 5466
rect 36642 5414 36656 5466
rect 36680 5414 36694 5466
rect 36694 5414 36706 5466
rect 36706 5414 36736 5466
rect 36760 5414 36770 5466
rect 36770 5414 36816 5466
rect 36520 5412 36576 5414
rect 36600 5412 36656 5414
rect 36680 5412 36736 5414
rect 36760 5412 36816 5414
rect 36818 4936 36874 4992
rect 36520 4378 36576 4380
rect 36600 4378 36656 4380
rect 36680 4378 36736 4380
rect 36760 4378 36816 4380
rect 36520 4326 36566 4378
rect 36566 4326 36576 4378
rect 36600 4326 36630 4378
rect 36630 4326 36642 4378
rect 36642 4326 36656 4378
rect 36680 4326 36694 4378
rect 36694 4326 36706 4378
rect 36706 4326 36736 4378
rect 36760 4326 36770 4378
rect 36770 4326 36816 4378
rect 36520 4324 36576 4326
rect 36600 4324 36656 4326
rect 36680 4324 36736 4326
rect 36760 4324 36816 4326
rect 37370 8900 37426 8936
rect 37370 8880 37372 8900
rect 37372 8880 37424 8900
rect 37424 8880 37426 8900
rect 37186 8472 37242 8528
rect 37278 5616 37334 5672
rect 36520 3290 36576 3292
rect 36600 3290 36656 3292
rect 36680 3290 36736 3292
rect 36760 3290 36816 3292
rect 36520 3238 36566 3290
rect 36566 3238 36576 3290
rect 36600 3238 36630 3290
rect 36630 3238 36642 3290
rect 36642 3238 36656 3290
rect 36680 3238 36694 3290
rect 36694 3238 36706 3290
rect 36706 3238 36736 3290
rect 36760 3238 36770 3290
rect 36770 3238 36816 3290
rect 36520 3236 36576 3238
rect 36600 3236 36656 3238
rect 36680 3236 36736 3238
rect 36760 3236 36816 3238
rect 36910 2896 36966 2952
rect 36520 2202 36576 2204
rect 36600 2202 36656 2204
rect 36680 2202 36736 2204
rect 36760 2202 36816 2204
rect 36520 2150 36566 2202
rect 36566 2150 36576 2202
rect 36600 2150 36630 2202
rect 36630 2150 36642 2202
rect 36642 2150 36656 2202
rect 36680 2150 36694 2202
rect 36694 2150 36706 2202
rect 36706 2150 36736 2202
rect 36760 2150 36770 2202
rect 36770 2150 36816 2202
rect 36520 2148 36576 2150
rect 36600 2148 36656 2150
rect 36680 2148 36736 2150
rect 36760 2148 36816 2150
rect 37278 1400 37334 1456
rect 37554 4936 37610 4992
rect 37830 6432 37886 6488
rect 37830 6160 37886 6216
rect 37738 4664 37794 4720
rect 37922 5072 37978 5128
rect 37922 3576 37978 3632
rect 37554 2760 37610 2816
rect 66580 12538 66636 12540
rect 66660 12538 66716 12540
rect 66740 12538 66796 12540
rect 66820 12538 66876 12540
rect 66580 12486 66626 12538
rect 66626 12486 66636 12538
rect 66660 12486 66690 12538
rect 66690 12486 66702 12538
rect 66702 12486 66716 12538
rect 66740 12486 66754 12538
rect 66754 12486 66766 12538
rect 66766 12486 66796 12538
rect 66820 12486 66830 12538
rect 66830 12486 66876 12538
rect 66580 12484 66636 12486
rect 66660 12484 66716 12486
rect 66740 12484 66796 12486
rect 66820 12484 66876 12486
rect 67240 11994 67296 11996
rect 67320 11994 67376 11996
rect 67400 11994 67456 11996
rect 67480 11994 67536 11996
rect 67240 11942 67286 11994
rect 67286 11942 67296 11994
rect 67320 11942 67350 11994
rect 67350 11942 67362 11994
rect 67362 11942 67376 11994
rect 67400 11942 67414 11994
rect 67414 11942 67426 11994
rect 67426 11942 67456 11994
rect 67480 11942 67490 11994
rect 67490 11942 67536 11994
rect 67240 11940 67296 11942
rect 67320 11940 67376 11942
rect 67400 11940 67456 11942
rect 67480 11940 67536 11942
rect 38198 7928 38254 7984
rect 38106 6704 38162 6760
rect 38658 8336 38714 8392
rect 38566 6568 38622 6624
rect 38474 6432 38530 6488
rect 38474 6160 38530 6216
rect 38566 5888 38622 5944
rect 38658 3440 38714 3496
rect 38290 1808 38346 1864
rect 66580 11450 66636 11452
rect 66660 11450 66716 11452
rect 66740 11450 66796 11452
rect 66820 11450 66876 11452
rect 66580 11398 66626 11450
rect 66626 11398 66636 11450
rect 66660 11398 66690 11450
rect 66690 11398 66702 11450
rect 66702 11398 66716 11450
rect 66740 11398 66754 11450
rect 66754 11398 66766 11450
rect 66766 11398 66796 11450
rect 66820 11398 66830 11450
rect 66830 11398 66876 11450
rect 66580 11396 66636 11398
rect 66660 11396 66716 11398
rect 66740 11396 66796 11398
rect 66820 11396 66876 11398
rect 67240 10906 67296 10908
rect 67320 10906 67376 10908
rect 67400 10906 67456 10908
rect 67480 10906 67536 10908
rect 67240 10854 67286 10906
rect 67286 10854 67296 10906
rect 67320 10854 67350 10906
rect 67350 10854 67362 10906
rect 67362 10854 67376 10906
rect 67400 10854 67414 10906
rect 67414 10854 67426 10906
rect 67426 10854 67456 10906
rect 67480 10854 67490 10906
rect 67490 10854 67536 10906
rect 67240 10852 67296 10854
rect 67320 10852 67376 10854
rect 67400 10852 67456 10854
rect 67480 10852 67536 10854
rect 66580 10362 66636 10364
rect 66660 10362 66716 10364
rect 66740 10362 66796 10364
rect 66820 10362 66876 10364
rect 66580 10310 66626 10362
rect 66626 10310 66636 10362
rect 66660 10310 66690 10362
rect 66690 10310 66702 10362
rect 66702 10310 66716 10362
rect 66740 10310 66754 10362
rect 66754 10310 66766 10362
rect 66766 10310 66796 10362
rect 66820 10310 66830 10362
rect 66830 10310 66876 10362
rect 66580 10308 66636 10310
rect 66660 10308 66716 10310
rect 66740 10308 66796 10310
rect 66820 10308 66876 10310
rect 67240 9818 67296 9820
rect 67320 9818 67376 9820
rect 67400 9818 67456 9820
rect 67480 9818 67536 9820
rect 67240 9766 67286 9818
rect 67286 9766 67296 9818
rect 67320 9766 67350 9818
rect 67350 9766 67362 9818
rect 67362 9766 67376 9818
rect 67400 9766 67414 9818
rect 67414 9766 67426 9818
rect 67426 9766 67456 9818
rect 67480 9766 67490 9818
rect 67490 9766 67536 9818
rect 67240 9764 67296 9766
rect 67320 9764 67376 9766
rect 67400 9764 67456 9766
rect 67480 9764 67536 9766
rect 66580 9274 66636 9276
rect 66660 9274 66716 9276
rect 66740 9274 66796 9276
rect 66820 9274 66876 9276
rect 66580 9222 66626 9274
rect 66626 9222 66636 9274
rect 66660 9222 66690 9274
rect 66690 9222 66702 9274
rect 66702 9222 66716 9274
rect 66740 9222 66754 9274
rect 66754 9222 66766 9274
rect 66766 9222 66796 9274
rect 66820 9222 66830 9274
rect 66830 9222 66876 9274
rect 66580 9220 66636 9222
rect 66660 9220 66716 9222
rect 66740 9220 66796 9222
rect 66820 9220 66876 9222
rect 67240 8730 67296 8732
rect 67320 8730 67376 8732
rect 67400 8730 67456 8732
rect 67480 8730 67536 8732
rect 67240 8678 67286 8730
rect 67286 8678 67296 8730
rect 67320 8678 67350 8730
rect 67350 8678 67362 8730
rect 67362 8678 67376 8730
rect 67400 8678 67414 8730
rect 67414 8678 67426 8730
rect 67426 8678 67456 8730
rect 67480 8678 67490 8730
rect 67490 8678 67536 8730
rect 67240 8676 67296 8678
rect 67320 8676 67376 8678
rect 67400 8676 67456 8678
rect 67480 8676 67536 8678
rect 38934 6332 38936 6352
rect 38936 6332 38988 6352
rect 38988 6332 38990 6352
rect 38934 6296 38990 6332
rect 39394 6860 39450 6896
rect 39394 6840 39396 6860
rect 39396 6840 39448 6860
rect 39448 6840 39450 6860
rect 39486 6296 39542 6352
rect 40222 5752 40278 5808
rect 66580 8186 66636 8188
rect 66660 8186 66716 8188
rect 66740 8186 66796 8188
rect 66820 8186 66876 8188
rect 66580 8134 66626 8186
rect 66626 8134 66636 8186
rect 66660 8134 66690 8186
rect 66690 8134 66702 8186
rect 66702 8134 66716 8186
rect 66740 8134 66754 8186
rect 66754 8134 66766 8186
rect 66766 8134 66796 8186
rect 66820 8134 66830 8186
rect 66830 8134 66876 8186
rect 66580 8132 66636 8134
rect 66660 8132 66716 8134
rect 66740 8132 66796 8134
rect 66820 8132 66876 8134
rect 67240 7642 67296 7644
rect 67320 7642 67376 7644
rect 67400 7642 67456 7644
rect 67480 7642 67536 7644
rect 67240 7590 67286 7642
rect 67286 7590 67296 7642
rect 67320 7590 67350 7642
rect 67350 7590 67362 7642
rect 67362 7590 67376 7642
rect 67400 7590 67414 7642
rect 67414 7590 67426 7642
rect 67426 7590 67456 7642
rect 67480 7590 67490 7642
rect 67490 7590 67536 7642
rect 67240 7588 67296 7590
rect 67320 7588 67376 7590
rect 67400 7588 67456 7590
rect 67480 7588 67536 7590
rect 66580 7098 66636 7100
rect 66660 7098 66716 7100
rect 66740 7098 66796 7100
rect 66820 7098 66876 7100
rect 66580 7046 66626 7098
rect 66626 7046 66636 7098
rect 66660 7046 66690 7098
rect 66690 7046 66702 7098
rect 66702 7046 66716 7098
rect 66740 7046 66754 7098
rect 66754 7046 66766 7098
rect 66766 7046 66796 7098
rect 66820 7046 66830 7098
rect 66830 7046 66876 7098
rect 66580 7044 66636 7046
rect 66660 7044 66716 7046
rect 66740 7044 66796 7046
rect 66820 7044 66876 7046
rect 42982 3068 42984 3088
rect 42984 3068 43036 3088
rect 43036 3068 43038 3088
rect 42982 3032 43038 3068
rect 41786 2352 41842 2408
rect 67240 6554 67296 6556
rect 67320 6554 67376 6556
rect 67400 6554 67456 6556
rect 67480 6554 67536 6556
rect 67240 6502 67286 6554
rect 67286 6502 67296 6554
rect 67320 6502 67350 6554
rect 67350 6502 67362 6554
rect 67362 6502 67376 6554
rect 67400 6502 67414 6554
rect 67414 6502 67426 6554
rect 67426 6502 67456 6554
rect 67480 6502 67490 6554
rect 67490 6502 67536 6554
rect 67240 6500 67296 6502
rect 67320 6500 67376 6502
rect 67400 6500 67456 6502
rect 67480 6500 67536 6502
rect 66580 6010 66636 6012
rect 66660 6010 66716 6012
rect 66740 6010 66796 6012
rect 66820 6010 66876 6012
rect 66580 5958 66626 6010
rect 66626 5958 66636 6010
rect 66660 5958 66690 6010
rect 66690 5958 66702 6010
rect 66702 5958 66716 6010
rect 66740 5958 66754 6010
rect 66754 5958 66766 6010
rect 66766 5958 66796 6010
rect 66820 5958 66830 6010
rect 66830 5958 66876 6010
rect 66580 5956 66636 5958
rect 66660 5956 66716 5958
rect 66740 5956 66796 5958
rect 66820 5956 66876 5958
rect 44914 5208 44970 5264
rect 67240 5466 67296 5468
rect 67320 5466 67376 5468
rect 67400 5466 67456 5468
rect 67480 5466 67536 5468
rect 67240 5414 67286 5466
rect 67286 5414 67296 5466
rect 67320 5414 67350 5466
rect 67350 5414 67362 5466
rect 67362 5414 67376 5466
rect 67400 5414 67414 5466
rect 67414 5414 67426 5466
rect 67426 5414 67456 5466
rect 67480 5414 67490 5466
rect 67490 5414 67536 5466
rect 67240 5412 67296 5414
rect 67320 5412 67376 5414
rect 67400 5412 67456 5414
rect 67480 5412 67536 5414
rect 66580 4922 66636 4924
rect 66660 4922 66716 4924
rect 66740 4922 66796 4924
rect 66820 4922 66876 4924
rect 66580 4870 66626 4922
rect 66626 4870 66636 4922
rect 66660 4870 66690 4922
rect 66690 4870 66702 4922
rect 66702 4870 66716 4922
rect 66740 4870 66754 4922
rect 66754 4870 66766 4922
rect 66766 4870 66796 4922
rect 66820 4870 66830 4922
rect 66830 4870 66876 4922
rect 66580 4868 66636 4870
rect 66660 4868 66716 4870
rect 66740 4868 66796 4870
rect 66820 4868 66876 4870
rect 51078 4664 51134 4720
rect 67240 4378 67296 4380
rect 67320 4378 67376 4380
rect 67400 4378 67456 4380
rect 67480 4378 67536 4380
rect 67240 4326 67286 4378
rect 67286 4326 67296 4378
rect 67320 4326 67350 4378
rect 67350 4326 67362 4378
rect 67362 4326 67376 4378
rect 67400 4326 67414 4378
rect 67414 4326 67426 4378
rect 67426 4326 67456 4378
rect 67480 4326 67490 4378
rect 67490 4326 67536 4378
rect 67240 4324 67296 4326
rect 67320 4324 67376 4326
rect 67400 4324 67456 4326
rect 67480 4324 67536 4326
rect 52642 4156 52644 4176
rect 52644 4156 52696 4176
rect 52696 4156 52698 4176
rect 52642 4120 52698 4156
rect 66580 3834 66636 3836
rect 66660 3834 66716 3836
rect 66740 3834 66796 3836
rect 66820 3834 66876 3836
rect 66580 3782 66626 3834
rect 66626 3782 66636 3834
rect 66660 3782 66690 3834
rect 66690 3782 66702 3834
rect 66702 3782 66716 3834
rect 66740 3782 66754 3834
rect 66754 3782 66766 3834
rect 66766 3782 66796 3834
rect 66820 3782 66830 3834
rect 66830 3782 66876 3834
rect 66580 3780 66636 3782
rect 66660 3780 66716 3782
rect 66740 3780 66796 3782
rect 66820 3780 66876 3782
rect 67240 3290 67296 3292
rect 67320 3290 67376 3292
rect 67400 3290 67456 3292
rect 67480 3290 67536 3292
rect 67240 3238 67286 3290
rect 67286 3238 67296 3290
rect 67320 3238 67350 3290
rect 67350 3238 67362 3290
rect 67362 3238 67376 3290
rect 67400 3238 67414 3290
rect 67414 3238 67426 3290
rect 67426 3238 67456 3290
rect 67480 3238 67490 3290
rect 67490 3238 67536 3290
rect 67240 3236 67296 3238
rect 67320 3236 67376 3238
rect 67400 3236 67456 3238
rect 67480 3236 67536 3238
rect 66580 2746 66636 2748
rect 66660 2746 66716 2748
rect 66740 2746 66796 2748
rect 66820 2746 66876 2748
rect 66580 2694 66626 2746
rect 66626 2694 66636 2746
rect 66660 2694 66690 2746
rect 66690 2694 66702 2746
rect 66702 2694 66716 2746
rect 66740 2694 66754 2746
rect 66754 2694 66766 2746
rect 66766 2694 66796 2746
rect 66820 2694 66830 2746
rect 66830 2694 66876 2746
rect 66580 2692 66636 2694
rect 66660 2692 66716 2694
rect 66740 2692 66796 2694
rect 66820 2692 66876 2694
rect 74078 3712 74134 3768
rect 67240 2202 67296 2204
rect 67320 2202 67376 2204
rect 67400 2202 67456 2204
rect 67480 2202 67536 2204
rect 67240 2150 67286 2202
rect 67286 2150 67296 2202
rect 67320 2150 67350 2202
rect 67350 2150 67362 2202
rect 67362 2150 67376 2202
rect 67400 2150 67414 2202
rect 67414 2150 67426 2202
rect 67426 2150 67456 2202
rect 67480 2150 67490 2202
rect 67490 2150 67536 2202
rect 67240 2148 67296 2150
rect 67320 2148 67376 2150
rect 67400 2148 67456 2150
rect 67480 2148 67536 2150
<< metal3 >>
rect 5130 37568 5446 37569
rect 5130 37504 5136 37568
rect 5200 37504 5216 37568
rect 5280 37504 5296 37568
rect 5360 37504 5376 37568
rect 5440 37504 5446 37568
rect 5130 37503 5446 37504
rect 35850 37568 36166 37569
rect 35850 37504 35856 37568
rect 35920 37504 35936 37568
rect 36000 37504 36016 37568
rect 36080 37504 36096 37568
rect 36160 37504 36166 37568
rect 35850 37503 36166 37504
rect 66570 37568 66886 37569
rect 66570 37504 66576 37568
rect 66640 37504 66656 37568
rect 66720 37504 66736 37568
rect 66800 37504 66816 37568
rect 66880 37504 66886 37568
rect 66570 37503 66886 37504
rect 5790 37024 6106 37025
rect 5790 36960 5796 37024
rect 5860 36960 5876 37024
rect 5940 36960 5956 37024
rect 6020 36960 6036 37024
rect 6100 36960 6106 37024
rect 5790 36959 6106 36960
rect 36510 37024 36826 37025
rect 36510 36960 36516 37024
rect 36580 36960 36596 37024
rect 36660 36960 36676 37024
rect 36740 36960 36756 37024
rect 36820 36960 36826 37024
rect 36510 36959 36826 36960
rect 67230 37024 67546 37025
rect 67230 36960 67236 37024
rect 67300 36960 67316 37024
rect 67380 36960 67396 37024
rect 67460 36960 67476 37024
rect 67540 36960 67546 37024
rect 67230 36959 67546 36960
rect 7005 36548 7071 36549
rect 32765 36548 32831 36549
rect 7005 36544 7052 36548
rect 7116 36546 7122 36548
rect 7005 36488 7010 36544
rect 7005 36484 7052 36488
rect 7116 36486 7162 36546
rect 32765 36544 32812 36548
rect 32876 36546 32882 36548
rect 32765 36488 32770 36544
rect 7116 36484 7122 36486
rect 32765 36484 32812 36488
rect 32876 36486 32922 36546
rect 32876 36484 32882 36486
rect 7005 36483 7071 36484
rect 32765 36483 32831 36484
rect 5130 36480 5446 36481
rect 5130 36416 5136 36480
rect 5200 36416 5216 36480
rect 5280 36416 5296 36480
rect 5360 36416 5376 36480
rect 5440 36416 5446 36480
rect 5130 36415 5446 36416
rect 35850 36480 36166 36481
rect 35850 36416 35856 36480
rect 35920 36416 35936 36480
rect 36000 36416 36016 36480
rect 36080 36416 36096 36480
rect 36160 36416 36166 36480
rect 35850 36415 36166 36416
rect 66570 36480 66886 36481
rect 66570 36416 66576 36480
rect 66640 36416 66656 36480
rect 66720 36416 66736 36480
rect 66800 36416 66816 36480
rect 66880 36416 66886 36480
rect 66570 36415 66886 36416
rect 5790 35936 6106 35937
rect 5790 35872 5796 35936
rect 5860 35872 5876 35936
rect 5940 35872 5956 35936
rect 6020 35872 6036 35936
rect 6100 35872 6106 35936
rect 5790 35871 6106 35872
rect 36510 35936 36826 35937
rect 36510 35872 36516 35936
rect 36580 35872 36596 35936
rect 36660 35872 36676 35936
rect 36740 35872 36756 35936
rect 36820 35872 36826 35936
rect 36510 35871 36826 35872
rect 67230 35936 67546 35937
rect 67230 35872 67236 35936
rect 67300 35872 67316 35936
rect 67380 35872 67396 35936
rect 67460 35872 67476 35936
rect 67540 35872 67546 35936
rect 67230 35871 67546 35872
rect 5130 35392 5446 35393
rect 5130 35328 5136 35392
rect 5200 35328 5216 35392
rect 5280 35328 5296 35392
rect 5360 35328 5376 35392
rect 5440 35328 5446 35392
rect 5130 35327 5446 35328
rect 35850 35392 36166 35393
rect 35850 35328 35856 35392
rect 35920 35328 35936 35392
rect 36000 35328 36016 35392
rect 36080 35328 36096 35392
rect 36160 35328 36166 35392
rect 35850 35327 36166 35328
rect 66570 35392 66886 35393
rect 66570 35328 66576 35392
rect 66640 35328 66656 35392
rect 66720 35328 66736 35392
rect 66800 35328 66816 35392
rect 66880 35328 66886 35392
rect 66570 35327 66886 35328
rect 5790 34848 6106 34849
rect 5790 34784 5796 34848
rect 5860 34784 5876 34848
rect 5940 34784 5956 34848
rect 6020 34784 6036 34848
rect 6100 34784 6106 34848
rect 5790 34783 6106 34784
rect 36510 34848 36826 34849
rect 36510 34784 36516 34848
rect 36580 34784 36596 34848
rect 36660 34784 36676 34848
rect 36740 34784 36756 34848
rect 36820 34784 36826 34848
rect 36510 34783 36826 34784
rect 67230 34848 67546 34849
rect 67230 34784 67236 34848
rect 67300 34784 67316 34848
rect 67380 34784 67396 34848
rect 67460 34784 67476 34848
rect 67540 34784 67546 34848
rect 67230 34783 67546 34784
rect 5130 34304 5446 34305
rect 5130 34240 5136 34304
rect 5200 34240 5216 34304
rect 5280 34240 5296 34304
rect 5360 34240 5376 34304
rect 5440 34240 5446 34304
rect 5130 34239 5446 34240
rect 35850 34304 36166 34305
rect 35850 34240 35856 34304
rect 35920 34240 35936 34304
rect 36000 34240 36016 34304
rect 36080 34240 36096 34304
rect 36160 34240 36166 34304
rect 35850 34239 36166 34240
rect 66570 34304 66886 34305
rect 66570 34240 66576 34304
rect 66640 34240 66656 34304
rect 66720 34240 66736 34304
rect 66800 34240 66816 34304
rect 66880 34240 66886 34304
rect 66570 34239 66886 34240
rect 5790 33760 6106 33761
rect 5790 33696 5796 33760
rect 5860 33696 5876 33760
rect 5940 33696 5956 33760
rect 6020 33696 6036 33760
rect 6100 33696 6106 33760
rect 5790 33695 6106 33696
rect 36510 33760 36826 33761
rect 36510 33696 36516 33760
rect 36580 33696 36596 33760
rect 36660 33696 36676 33760
rect 36740 33696 36756 33760
rect 36820 33696 36826 33760
rect 36510 33695 36826 33696
rect 67230 33760 67546 33761
rect 67230 33696 67236 33760
rect 67300 33696 67316 33760
rect 67380 33696 67396 33760
rect 67460 33696 67476 33760
rect 67540 33696 67546 33760
rect 67230 33695 67546 33696
rect 5130 33216 5446 33217
rect 5130 33152 5136 33216
rect 5200 33152 5216 33216
rect 5280 33152 5296 33216
rect 5360 33152 5376 33216
rect 5440 33152 5446 33216
rect 5130 33151 5446 33152
rect 35850 33216 36166 33217
rect 35850 33152 35856 33216
rect 35920 33152 35936 33216
rect 36000 33152 36016 33216
rect 36080 33152 36096 33216
rect 36160 33152 36166 33216
rect 35850 33151 36166 33152
rect 66570 33216 66886 33217
rect 66570 33152 66576 33216
rect 66640 33152 66656 33216
rect 66720 33152 66736 33216
rect 66800 33152 66816 33216
rect 66880 33152 66886 33216
rect 66570 33151 66886 33152
rect 5790 32672 6106 32673
rect 5790 32608 5796 32672
rect 5860 32608 5876 32672
rect 5940 32608 5956 32672
rect 6020 32608 6036 32672
rect 6100 32608 6106 32672
rect 5790 32607 6106 32608
rect 36510 32672 36826 32673
rect 36510 32608 36516 32672
rect 36580 32608 36596 32672
rect 36660 32608 36676 32672
rect 36740 32608 36756 32672
rect 36820 32608 36826 32672
rect 36510 32607 36826 32608
rect 67230 32672 67546 32673
rect 67230 32608 67236 32672
rect 67300 32608 67316 32672
rect 67380 32608 67396 32672
rect 67460 32608 67476 32672
rect 67540 32608 67546 32672
rect 67230 32607 67546 32608
rect 5130 32128 5446 32129
rect 5130 32064 5136 32128
rect 5200 32064 5216 32128
rect 5280 32064 5296 32128
rect 5360 32064 5376 32128
rect 5440 32064 5446 32128
rect 5130 32063 5446 32064
rect 35850 32128 36166 32129
rect 35850 32064 35856 32128
rect 35920 32064 35936 32128
rect 36000 32064 36016 32128
rect 36080 32064 36096 32128
rect 36160 32064 36166 32128
rect 35850 32063 36166 32064
rect 66570 32128 66886 32129
rect 66570 32064 66576 32128
rect 66640 32064 66656 32128
rect 66720 32064 66736 32128
rect 66800 32064 66816 32128
rect 66880 32064 66886 32128
rect 66570 32063 66886 32064
rect 5790 31584 6106 31585
rect 5790 31520 5796 31584
rect 5860 31520 5876 31584
rect 5940 31520 5956 31584
rect 6020 31520 6036 31584
rect 6100 31520 6106 31584
rect 5790 31519 6106 31520
rect 36510 31584 36826 31585
rect 36510 31520 36516 31584
rect 36580 31520 36596 31584
rect 36660 31520 36676 31584
rect 36740 31520 36756 31584
rect 36820 31520 36826 31584
rect 36510 31519 36826 31520
rect 67230 31584 67546 31585
rect 67230 31520 67236 31584
rect 67300 31520 67316 31584
rect 67380 31520 67396 31584
rect 67460 31520 67476 31584
rect 67540 31520 67546 31584
rect 67230 31519 67546 31520
rect 5130 31040 5446 31041
rect 5130 30976 5136 31040
rect 5200 30976 5216 31040
rect 5280 30976 5296 31040
rect 5360 30976 5376 31040
rect 5440 30976 5446 31040
rect 5130 30975 5446 30976
rect 35850 31040 36166 31041
rect 35850 30976 35856 31040
rect 35920 30976 35936 31040
rect 36000 30976 36016 31040
rect 36080 30976 36096 31040
rect 36160 30976 36166 31040
rect 35850 30975 36166 30976
rect 66570 31040 66886 31041
rect 66570 30976 66576 31040
rect 66640 30976 66656 31040
rect 66720 30976 66736 31040
rect 66800 30976 66816 31040
rect 66880 30976 66886 31040
rect 66570 30975 66886 30976
rect 5790 30496 6106 30497
rect 5790 30432 5796 30496
rect 5860 30432 5876 30496
rect 5940 30432 5956 30496
rect 6020 30432 6036 30496
rect 6100 30432 6106 30496
rect 5790 30431 6106 30432
rect 36510 30496 36826 30497
rect 36510 30432 36516 30496
rect 36580 30432 36596 30496
rect 36660 30432 36676 30496
rect 36740 30432 36756 30496
rect 36820 30432 36826 30496
rect 36510 30431 36826 30432
rect 67230 30496 67546 30497
rect 67230 30432 67236 30496
rect 67300 30432 67316 30496
rect 67380 30432 67396 30496
rect 67460 30432 67476 30496
rect 67540 30432 67546 30496
rect 67230 30431 67546 30432
rect 5130 29952 5446 29953
rect 5130 29888 5136 29952
rect 5200 29888 5216 29952
rect 5280 29888 5296 29952
rect 5360 29888 5376 29952
rect 5440 29888 5446 29952
rect 5130 29887 5446 29888
rect 35850 29952 36166 29953
rect 35850 29888 35856 29952
rect 35920 29888 35936 29952
rect 36000 29888 36016 29952
rect 36080 29888 36096 29952
rect 36160 29888 36166 29952
rect 35850 29887 36166 29888
rect 66570 29952 66886 29953
rect 66570 29888 66576 29952
rect 66640 29888 66656 29952
rect 66720 29888 66736 29952
rect 66800 29888 66816 29952
rect 66880 29888 66886 29952
rect 66570 29887 66886 29888
rect 18965 29610 19031 29613
rect 27470 29610 27476 29612
rect 18965 29608 27476 29610
rect 18965 29552 18970 29608
rect 19026 29552 27476 29608
rect 18965 29550 27476 29552
rect 18965 29547 19031 29550
rect 27470 29548 27476 29550
rect 27540 29548 27546 29612
rect 5790 29408 6106 29409
rect 5790 29344 5796 29408
rect 5860 29344 5876 29408
rect 5940 29344 5956 29408
rect 6020 29344 6036 29408
rect 6100 29344 6106 29408
rect 5790 29343 6106 29344
rect 36510 29408 36826 29409
rect 36510 29344 36516 29408
rect 36580 29344 36596 29408
rect 36660 29344 36676 29408
rect 36740 29344 36756 29408
rect 36820 29344 36826 29408
rect 36510 29343 36826 29344
rect 67230 29408 67546 29409
rect 67230 29344 67236 29408
rect 67300 29344 67316 29408
rect 67380 29344 67396 29408
rect 67460 29344 67476 29408
rect 67540 29344 67546 29408
rect 67230 29343 67546 29344
rect 5130 28864 5446 28865
rect 5130 28800 5136 28864
rect 5200 28800 5216 28864
rect 5280 28800 5296 28864
rect 5360 28800 5376 28864
rect 5440 28800 5446 28864
rect 5130 28799 5446 28800
rect 35850 28864 36166 28865
rect 35850 28800 35856 28864
rect 35920 28800 35936 28864
rect 36000 28800 36016 28864
rect 36080 28800 36096 28864
rect 36160 28800 36166 28864
rect 35850 28799 36166 28800
rect 66570 28864 66886 28865
rect 66570 28800 66576 28864
rect 66640 28800 66656 28864
rect 66720 28800 66736 28864
rect 66800 28800 66816 28864
rect 66880 28800 66886 28864
rect 66570 28799 66886 28800
rect 5790 28320 6106 28321
rect 5790 28256 5796 28320
rect 5860 28256 5876 28320
rect 5940 28256 5956 28320
rect 6020 28256 6036 28320
rect 6100 28256 6106 28320
rect 5790 28255 6106 28256
rect 36510 28320 36826 28321
rect 36510 28256 36516 28320
rect 36580 28256 36596 28320
rect 36660 28256 36676 28320
rect 36740 28256 36756 28320
rect 36820 28256 36826 28320
rect 36510 28255 36826 28256
rect 67230 28320 67546 28321
rect 67230 28256 67236 28320
rect 67300 28256 67316 28320
rect 67380 28256 67396 28320
rect 67460 28256 67476 28320
rect 67540 28256 67546 28320
rect 67230 28255 67546 28256
rect 5130 27776 5446 27777
rect 5130 27712 5136 27776
rect 5200 27712 5216 27776
rect 5280 27712 5296 27776
rect 5360 27712 5376 27776
rect 5440 27712 5446 27776
rect 5130 27711 5446 27712
rect 35850 27776 36166 27777
rect 35850 27712 35856 27776
rect 35920 27712 35936 27776
rect 36000 27712 36016 27776
rect 36080 27712 36096 27776
rect 36160 27712 36166 27776
rect 35850 27711 36166 27712
rect 66570 27776 66886 27777
rect 66570 27712 66576 27776
rect 66640 27712 66656 27776
rect 66720 27712 66736 27776
rect 66800 27712 66816 27776
rect 66880 27712 66886 27776
rect 66570 27711 66886 27712
rect 5790 27232 6106 27233
rect 5790 27168 5796 27232
rect 5860 27168 5876 27232
rect 5940 27168 5956 27232
rect 6020 27168 6036 27232
rect 6100 27168 6106 27232
rect 5790 27167 6106 27168
rect 36510 27232 36826 27233
rect 36510 27168 36516 27232
rect 36580 27168 36596 27232
rect 36660 27168 36676 27232
rect 36740 27168 36756 27232
rect 36820 27168 36826 27232
rect 36510 27167 36826 27168
rect 67230 27232 67546 27233
rect 67230 27168 67236 27232
rect 67300 27168 67316 27232
rect 67380 27168 67396 27232
rect 67460 27168 67476 27232
rect 67540 27168 67546 27232
rect 67230 27167 67546 27168
rect 10869 26890 10935 26893
rect 28390 26890 28396 26892
rect 10869 26888 28396 26890
rect 10869 26832 10874 26888
rect 10930 26832 28396 26888
rect 10869 26830 28396 26832
rect 10869 26827 10935 26830
rect 28390 26828 28396 26830
rect 28460 26828 28466 26892
rect 5130 26688 5446 26689
rect 5130 26624 5136 26688
rect 5200 26624 5216 26688
rect 5280 26624 5296 26688
rect 5360 26624 5376 26688
rect 5440 26624 5446 26688
rect 5130 26623 5446 26624
rect 35850 26688 36166 26689
rect 35850 26624 35856 26688
rect 35920 26624 35936 26688
rect 36000 26624 36016 26688
rect 36080 26624 36096 26688
rect 36160 26624 36166 26688
rect 35850 26623 36166 26624
rect 66570 26688 66886 26689
rect 66570 26624 66576 26688
rect 66640 26624 66656 26688
rect 66720 26624 66736 26688
rect 66800 26624 66816 26688
rect 66880 26624 66886 26688
rect 66570 26623 66886 26624
rect 5790 26144 6106 26145
rect 5790 26080 5796 26144
rect 5860 26080 5876 26144
rect 5940 26080 5956 26144
rect 6020 26080 6036 26144
rect 6100 26080 6106 26144
rect 5790 26079 6106 26080
rect 36510 26144 36826 26145
rect 36510 26080 36516 26144
rect 36580 26080 36596 26144
rect 36660 26080 36676 26144
rect 36740 26080 36756 26144
rect 36820 26080 36826 26144
rect 36510 26079 36826 26080
rect 67230 26144 67546 26145
rect 67230 26080 67236 26144
rect 67300 26080 67316 26144
rect 67380 26080 67396 26144
rect 67460 26080 67476 26144
rect 67540 26080 67546 26144
rect 67230 26079 67546 26080
rect 5130 25600 5446 25601
rect 5130 25536 5136 25600
rect 5200 25536 5216 25600
rect 5280 25536 5296 25600
rect 5360 25536 5376 25600
rect 5440 25536 5446 25600
rect 5130 25535 5446 25536
rect 35850 25600 36166 25601
rect 35850 25536 35856 25600
rect 35920 25536 35936 25600
rect 36000 25536 36016 25600
rect 36080 25536 36096 25600
rect 36160 25536 36166 25600
rect 35850 25535 36166 25536
rect 66570 25600 66886 25601
rect 66570 25536 66576 25600
rect 66640 25536 66656 25600
rect 66720 25536 66736 25600
rect 66800 25536 66816 25600
rect 66880 25536 66886 25600
rect 66570 25535 66886 25536
rect 5790 25056 6106 25057
rect 5790 24992 5796 25056
rect 5860 24992 5876 25056
rect 5940 24992 5956 25056
rect 6020 24992 6036 25056
rect 6100 24992 6106 25056
rect 5790 24991 6106 24992
rect 36510 25056 36826 25057
rect 36510 24992 36516 25056
rect 36580 24992 36596 25056
rect 36660 24992 36676 25056
rect 36740 24992 36756 25056
rect 36820 24992 36826 25056
rect 36510 24991 36826 24992
rect 67230 25056 67546 25057
rect 67230 24992 67236 25056
rect 67300 24992 67316 25056
rect 67380 24992 67396 25056
rect 67460 24992 67476 25056
rect 67540 24992 67546 25056
rect 67230 24991 67546 24992
rect 5130 24512 5446 24513
rect 5130 24448 5136 24512
rect 5200 24448 5216 24512
rect 5280 24448 5296 24512
rect 5360 24448 5376 24512
rect 5440 24448 5446 24512
rect 5130 24447 5446 24448
rect 35850 24512 36166 24513
rect 35850 24448 35856 24512
rect 35920 24448 35936 24512
rect 36000 24448 36016 24512
rect 36080 24448 36096 24512
rect 36160 24448 36166 24512
rect 35850 24447 36166 24448
rect 66570 24512 66886 24513
rect 66570 24448 66576 24512
rect 66640 24448 66656 24512
rect 66720 24448 66736 24512
rect 66800 24448 66816 24512
rect 66880 24448 66886 24512
rect 66570 24447 66886 24448
rect 3509 24170 3575 24173
rect 35014 24170 35020 24172
rect 3509 24168 35020 24170
rect 3509 24112 3514 24168
rect 3570 24112 35020 24168
rect 3509 24110 35020 24112
rect 3509 24107 3575 24110
rect 35014 24108 35020 24110
rect 35084 24108 35090 24172
rect 5790 23968 6106 23969
rect 5790 23904 5796 23968
rect 5860 23904 5876 23968
rect 5940 23904 5956 23968
rect 6020 23904 6036 23968
rect 6100 23904 6106 23968
rect 5790 23903 6106 23904
rect 36510 23968 36826 23969
rect 36510 23904 36516 23968
rect 36580 23904 36596 23968
rect 36660 23904 36676 23968
rect 36740 23904 36756 23968
rect 36820 23904 36826 23968
rect 36510 23903 36826 23904
rect 67230 23968 67546 23969
rect 67230 23904 67236 23968
rect 67300 23904 67316 23968
rect 67380 23904 67396 23968
rect 67460 23904 67476 23968
rect 67540 23904 67546 23968
rect 67230 23903 67546 23904
rect 5130 23424 5446 23425
rect 5130 23360 5136 23424
rect 5200 23360 5216 23424
rect 5280 23360 5296 23424
rect 5360 23360 5376 23424
rect 5440 23360 5446 23424
rect 5130 23359 5446 23360
rect 35850 23424 36166 23425
rect 35850 23360 35856 23424
rect 35920 23360 35936 23424
rect 36000 23360 36016 23424
rect 36080 23360 36096 23424
rect 36160 23360 36166 23424
rect 35850 23359 36166 23360
rect 66570 23424 66886 23425
rect 66570 23360 66576 23424
rect 66640 23360 66656 23424
rect 66720 23360 66736 23424
rect 66800 23360 66816 23424
rect 66880 23360 66886 23424
rect 66570 23359 66886 23360
rect 5790 22880 6106 22881
rect 5790 22816 5796 22880
rect 5860 22816 5876 22880
rect 5940 22816 5956 22880
rect 6020 22816 6036 22880
rect 6100 22816 6106 22880
rect 5790 22815 6106 22816
rect 36510 22880 36826 22881
rect 36510 22816 36516 22880
rect 36580 22816 36596 22880
rect 36660 22816 36676 22880
rect 36740 22816 36756 22880
rect 36820 22816 36826 22880
rect 36510 22815 36826 22816
rect 67230 22880 67546 22881
rect 67230 22816 67236 22880
rect 67300 22816 67316 22880
rect 67380 22816 67396 22880
rect 67460 22816 67476 22880
rect 67540 22816 67546 22880
rect 67230 22815 67546 22816
rect 5130 22336 5446 22337
rect 5130 22272 5136 22336
rect 5200 22272 5216 22336
rect 5280 22272 5296 22336
rect 5360 22272 5376 22336
rect 5440 22272 5446 22336
rect 5130 22271 5446 22272
rect 35850 22336 36166 22337
rect 35850 22272 35856 22336
rect 35920 22272 35936 22336
rect 36000 22272 36016 22336
rect 36080 22272 36096 22336
rect 36160 22272 36166 22336
rect 35850 22271 36166 22272
rect 66570 22336 66886 22337
rect 66570 22272 66576 22336
rect 66640 22272 66656 22336
rect 66720 22272 66736 22336
rect 66800 22272 66816 22336
rect 66880 22272 66886 22336
rect 66570 22271 66886 22272
rect 5790 21792 6106 21793
rect 5790 21728 5796 21792
rect 5860 21728 5876 21792
rect 5940 21728 5956 21792
rect 6020 21728 6036 21792
rect 6100 21728 6106 21792
rect 5790 21727 6106 21728
rect 36510 21792 36826 21793
rect 36510 21728 36516 21792
rect 36580 21728 36596 21792
rect 36660 21728 36676 21792
rect 36740 21728 36756 21792
rect 36820 21728 36826 21792
rect 36510 21727 36826 21728
rect 67230 21792 67546 21793
rect 67230 21728 67236 21792
rect 67300 21728 67316 21792
rect 67380 21728 67396 21792
rect 67460 21728 67476 21792
rect 67540 21728 67546 21792
rect 67230 21727 67546 21728
rect 5130 21248 5446 21249
rect 5130 21184 5136 21248
rect 5200 21184 5216 21248
rect 5280 21184 5296 21248
rect 5360 21184 5376 21248
rect 5440 21184 5446 21248
rect 5130 21183 5446 21184
rect 35850 21248 36166 21249
rect 35850 21184 35856 21248
rect 35920 21184 35936 21248
rect 36000 21184 36016 21248
rect 36080 21184 36096 21248
rect 36160 21184 36166 21248
rect 35850 21183 36166 21184
rect 66570 21248 66886 21249
rect 66570 21184 66576 21248
rect 66640 21184 66656 21248
rect 66720 21184 66736 21248
rect 66800 21184 66816 21248
rect 66880 21184 66886 21248
rect 66570 21183 66886 21184
rect 5790 20704 6106 20705
rect 5790 20640 5796 20704
rect 5860 20640 5876 20704
rect 5940 20640 5956 20704
rect 6020 20640 6036 20704
rect 6100 20640 6106 20704
rect 5790 20639 6106 20640
rect 36510 20704 36826 20705
rect 36510 20640 36516 20704
rect 36580 20640 36596 20704
rect 36660 20640 36676 20704
rect 36740 20640 36756 20704
rect 36820 20640 36826 20704
rect 36510 20639 36826 20640
rect 67230 20704 67546 20705
rect 67230 20640 67236 20704
rect 67300 20640 67316 20704
rect 67380 20640 67396 20704
rect 67460 20640 67476 20704
rect 67540 20640 67546 20704
rect 67230 20639 67546 20640
rect 5130 20160 5446 20161
rect 5130 20096 5136 20160
rect 5200 20096 5216 20160
rect 5280 20096 5296 20160
rect 5360 20096 5376 20160
rect 5440 20096 5446 20160
rect 5130 20095 5446 20096
rect 35850 20160 36166 20161
rect 35850 20096 35856 20160
rect 35920 20096 35936 20160
rect 36000 20096 36016 20160
rect 36080 20096 36096 20160
rect 36160 20096 36166 20160
rect 35850 20095 36166 20096
rect 66570 20160 66886 20161
rect 66570 20096 66576 20160
rect 66640 20096 66656 20160
rect 66720 20096 66736 20160
rect 66800 20096 66816 20160
rect 66880 20096 66886 20160
rect 66570 20095 66886 20096
rect 5790 19616 6106 19617
rect 5790 19552 5796 19616
rect 5860 19552 5876 19616
rect 5940 19552 5956 19616
rect 6020 19552 6036 19616
rect 6100 19552 6106 19616
rect 5790 19551 6106 19552
rect 36510 19616 36826 19617
rect 36510 19552 36516 19616
rect 36580 19552 36596 19616
rect 36660 19552 36676 19616
rect 36740 19552 36756 19616
rect 36820 19552 36826 19616
rect 36510 19551 36826 19552
rect 67230 19616 67546 19617
rect 67230 19552 67236 19616
rect 67300 19552 67316 19616
rect 67380 19552 67396 19616
rect 67460 19552 67476 19616
rect 67540 19552 67546 19616
rect 67230 19551 67546 19552
rect 5130 19072 5446 19073
rect 5130 19008 5136 19072
rect 5200 19008 5216 19072
rect 5280 19008 5296 19072
rect 5360 19008 5376 19072
rect 5440 19008 5446 19072
rect 5130 19007 5446 19008
rect 35850 19072 36166 19073
rect 35850 19008 35856 19072
rect 35920 19008 35936 19072
rect 36000 19008 36016 19072
rect 36080 19008 36096 19072
rect 36160 19008 36166 19072
rect 35850 19007 36166 19008
rect 66570 19072 66886 19073
rect 66570 19008 66576 19072
rect 66640 19008 66656 19072
rect 66720 19008 66736 19072
rect 66800 19008 66816 19072
rect 66880 19008 66886 19072
rect 66570 19007 66886 19008
rect 5790 18528 6106 18529
rect 5790 18464 5796 18528
rect 5860 18464 5876 18528
rect 5940 18464 5956 18528
rect 6020 18464 6036 18528
rect 6100 18464 6106 18528
rect 5790 18463 6106 18464
rect 36510 18528 36826 18529
rect 36510 18464 36516 18528
rect 36580 18464 36596 18528
rect 36660 18464 36676 18528
rect 36740 18464 36756 18528
rect 36820 18464 36826 18528
rect 36510 18463 36826 18464
rect 67230 18528 67546 18529
rect 67230 18464 67236 18528
rect 67300 18464 67316 18528
rect 67380 18464 67396 18528
rect 67460 18464 67476 18528
rect 67540 18464 67546 18528
rect 67230 18463 67546 18464
rect 21909 18050 21975 18053
rect 27286 18050 27292 18052
rect 21909 18048 27292 18050
rect 21909 17992 21914 18048
rect 21970 17992 27292 18048
rect 21909 17990 27292 17992
rect 21909 17987 21975 17990
rect 27286 17988 27292 17990
rect 27356 17988 27362 18052
rect 5130 17984 5446 17985
rect 5130 17920 5136 17984
rect 5200 17920 5216 17984
rect 5280 17920 5296 17984
rect 5360 17920 5376 17984
rect 5440 17920 5446 17984
rect 5130 17919 5446 17920
rect 35850 17984 36166 17985
rect 35850 17920 35856 17984
rect 35920 17920 35936 17984
rect 36000 17920 36016 17984
rect 36080 17920 36096 17984
rect 36160 17920 36166 17984
rect 35850 17919 36166 17920
rect 66570 17984 66886 17985
rect 66570 17920 66576 17984
rect 66640 17920 66656 17984
rect 66720 17920 66736 17984
rect 66800 17920 66816 17984
rect 66880 17920 66886 17984
rect 66570 17919 66886 17920
rect 5790 17440 6106 17441
rect 5790 17376 5796 17440
rect 5860 17376 5876 17440
rect 5940 17376 5956 17440
rect 6020 17376 6036 17440
rect 6100 17376 6106 17440
rect 5790 17375 6106 17376
rect 36510 17440 36826 17441
rect 36510 17376 36516 17440
rect 36580 17376 36596 17440
rect 36660 17376 36676 17440
rect 36740 17376 36756 17440
rect 36820 17376 36826 17440
rect 36510 17375 36826 17376
rect 67230 17440 67546 17441
rect 67230 17376 67236 17440
rect 67300 17376 67316 17440
rect 67380 17376 67396 17440
rect 67460 17376 67476 17440
rect 67540 17376 67546 17440
rect 67230 17375 67546 17376
rect 5130 16896 5446 16897
rect 5130 16832 5136 16896
rect 5200 16832 5216 16896
rect 5280 16832 5296 16896
rect 5360 16832 5376 16896
rect 5440 16832 5446 16896
rect 5130 16831 5446 16832
rect 35850 16896 36166 16897
rect 35850 16832 35856 16896
rect 35920 16832 35936 16896
rect 36000 16832 36016 16896
rect 36080 16832 36096 16896
rect 36160 16832 36166 16896
rect 35850 16831 36166 16832
rect 66570 16896 66886 16897
rect 66570 16832 66576 16896
rect 66640 16832 66656 16896
rect 66720 16832 66736 16896
rect 66800 16832 66816 16896
rect 66880 16832 66886 16896
rect 66570 16831 66886 16832
rect 5790 16352 6106 16353
rect 5790 16288 5796 16352
rect 5860 16288 5876 16352
rect 5940 16288 5956 16352
rect 6020 16288 6036 16352
rect 6100 16288 6106 16352
rect 5790 16287 6106 16288
rect 36510 16352 36826 16353
rect 36510 16288 36516 16352
rect 36580 16288 36596 16352
rect 36660 16288 36676 16352
rect 36740 16288 36756 16352
rect 36820 16288 36826 16352
rect 36510 16287 36826 16288
rect 67230 16352 67546 16353
rect 67230 16288 67236 16352
rect 67300 16288 67316 16352
rect 67380 16288 67396 16352
rect 67460 16288 67476 16352
rect 67540 16288 67546 16352
rect 67230 16287 67546 16288
rect 5130 15808 5446 15809
rect 5130 15744 5136 15808
rect 5200 15744 5216 15808
rect 5280 15744 5296 15808
rect 5360 15744 5376 15808
rect 5440 15744 5446 15808
rect 5130 15743 5446 15744
rect 35850 15808 36166 15809
rect 35850 15744 35856 15808
rect 35920 15744 35936 15808
rect 36000 15744 36016 15808
rect 36080 15744 36096 15808
rect 36160 15744 36166 15808
rect 35850 15743 36166 15744
rect 66570 15808 66886 15809
rect 66570 15744 66576 15808
rect 66640 15744 66656 15808
rect 66720 15744 66736 15808
rect 66800 15744 66816 15808
rect 66880 15744 66886 15808
rect 66570 15743 66886 15744
rect 5790 15264 6106 15265
rect 5790 15200 5796 15264
rect 5860 15200 5876 15264
rect 5940 15200 5956 15264
rect 6020 15200 6036 15264
rect 6100 15200 6106 15264
rect 5790 15199 6106 15200
rect 36510 15264 36826 15265
rect 36510 15200 36516 15264
rect 36580 15200 36596 15264
rect 36660 15200 36676 15264
rect 36740 15200 36756 15264
rect 36820 15200 36826 15264
rect 36510 15199 36826 15200
rect 67230 15264 67546 15265
rect 67230 15200 67236 15264
rect 67300 15200 67316 15264
rect 67380 15200 67396 15264
rect 67460 15200 67476 15264
rect 67540 15200 67546 15264
rect 67230 15199 67546 15200
rect 5130 14720 5446 14721
rect 5130 14656 5136 14720
rect 5200 14656 5216 14720
rect 5280 14656 5296 14720
rect 5360 14656 5376 14720
rect 5440 14656 5446 14720
rect 5130 14655 5446 14656
rect 35850 14720 36166 14721
rect 35850 14656 35856 14720
rect 35920 14656 35936 14720
rect 36000 14656 36016 14720
rect 36080 14656 36096 14720
rect 36160 14656 36166 14720
rect 35850 14655 36166 14656
rect 66570 14720 66886 14721
rect 66570 14656 66576 14720
rect 66640 14656 66656 14720
rect 66720 14656 66736 14720
rect 66800 14656 66816 14720
rect 66880 14656 66886 14720
rect 66570 14655 66886 14656
rect 14549 14514 14615 14517
rect 28574 14514 28580 14516
rect 14549 14512 28580 14514
rect 14549 14456 14554 14512
rect 14610 14456 28580 14512
rect 14549 14454 28580 14456
rect 14549 14451 14615 14454
rect 28574 14452 28580 14454
rect 28644 14452 28650 14516
rect 39113 14514 39179 14517
rect 35850 14512 39179 14514
rect 35850 14456 39118 14512
rect 39174 14456 39179 14512
rect 35850 14454 39179 14456
rect 28206 14316 28212 14380
rect 28276 14378 28282 14380
rect 35850 14378 35910 14454
rect 39113 14451 39179 14454
rect 28276 14318 35910 14378
rect 28276 14316 28282 14318
rect 5790 14176 6106 14177
rect 5790 14112 5796 14176
rect 5860 14112 5876 14176
rect 5940 14112 5956 14176
rect 6020 14112 6036 14176
rect 6100 14112 6106 14176
rect 5790 14111 6106 14112
rect 36510 14176 36826 14177
rect 36510 14112 36516 14176
rect 36580 14112 36596 14176
rect 36660 14112 36676 14176
rect 36740 14112 36756 14176
rect 36820 14112 36826 14176
rect 36510 14111 36826 14112
rect 67230 14176 67546 14177
rect 67230 14112 67236 14176
rect 67300 14112 67316 14176
rect 67380 14112 67396 14176
rect 67460 14112 67476 14176
rect 67540 14112 67546 14176
rect 67230 14111 67546 14112
rect 5130 13632 5446 13633
rect 5130 13568 5136 13632
rect 5200 13568 5216 13632
rect 5280 13568 5296 13632
rect 5360 13568 5376 13632
rect 5440 13568 5446 13632
rect 5130 13567 5446 13568
rect 35850 13632 36166 13633
rect 35850 13568 35856 13632
rect 35920 13568 35936 13632
rect 36000 13568 36016 13632
rect 36080 13568 36096 13632
rect 36160 13568 36166 13632
rect 35850 13567 36166 13568
rect 66570 13632 66886 13633
rect 66570 13568 66576 13632
rect 66640 13568 66656 13632
rect 66720 13568 66736 13632
rect 66800 13568 66816 13632
rect 66880 13568 66886 13632
rect 66570 13567 66886 13568
rect 5790 13088 6106 13089
rect 5790 13024 5796 13088
rect 5860 13024 5876 13088
rect 5940 13024 5956 13088
rect 6020 13024 6036 13088
rect 6100 13024 6106 13088
rect 5790 13023 6106 13024
rect 36510 13088 36826 13089
rect 36510 13024 36516 13088
rect 36580 13024 36596 13088
rect 36660 13024 36676 13088
rect 36740 13024 36756 13088
rect 36820 13024 36826 13088
rect 36510 13023 36826 13024
rect 67230 13088 67546 13089
rect 67230 13024 67236 13088
rect 67300 13024 67316 13088
rect 67380 13024 67396 13088
rect 67460 13024 67476 13088
rect 67540 13024 67546 13088
rect 67230 13023 67546 13024
rect 5130 12544 5446 12545
rect 5130 12480 5136 12544
rect 5200 12480 5216 12544
rect 5280 12480 5296 12544
rect 5360 12480 5376 12544
rect 5440 12480 5446 12544
rect 5130 12479 5446 12480
rect 35850 12544 36166 12545
rect 35850 12480 35856 12544
rect 35920 12480 35936 12544
rect 36000 12480 36016 12544
rect 36080 12480 36096 12544
rect 36160 12480 36166 12544
rect 35850 12479 36166 12480
rect 66570 12544 66886 12545
rect 66570 12480 66576 12544
rect 66640 12480 66656 12544
rect 66720 12480 66736 12544
rect 66800 12480 66816 12544
rect 66880 12480 66886 12544
rect 66570 12479 66886 12480
rect 12750 12412 12756 12476
rect 12820 12474 12826 12476
rect 27705 12474 27771 12477
rect 12820 12472 27771 12474
rect 12820 12416 27710 12472
rect 27766 12416 27771 12472
rect 12820 12414 27771 12416
rect 12820 12412 12826 12414
rect 27705 12411 27771 12414
rect 24669 12202 24735 12205
rect 25681 12202 25747 12205
rect 24669 12200 25747 12202
rect 24669 12144 24674 12200
rect 24730 12144 25686 12200
rect 25742 12144 25747 12200
rect 24669 12142 25747 12144
rect 24669 12139 24735 12142
rect 25681 12139 25747 12142
rect 5790 12000 6106 12001
rect 5790 11936 5796 12000
rect 5860 11936 5876 12000
rect 5940 11936 5956 12000
rect 6020 11936 6036 12000
rect 6100 11936 6106 12000
rect 5790 11935 6106 11936
rect 36510 12000 36826 12001
rect 36510 11936 36516 12000
rect 36580 11936 36596 12000
rect 36660 11936 36676 12000
rect 36740 11936 36756 12000
rect 36820 11936 36826 12000
rect 36510 11935 36826 11936
rect 67230 12000 67546 12001
rect 67230 11936 67236 12000
rect 67300 11936 67316 12000
rect 67380 11936 67396 12000
rect 67460 11936 67476 12000
rect 67540 11936 67546 12000
rect 67230 11935 67546 11936
rect 19926 11460 19932 11524
rect 19996 11522 20002 11524
rect 28165 11522 28231 11525
rect 19996 11520 28231 11522
rect 19996 11464 28170 11520
rect 28226 11464 28231 11520
rect 19996 11462 28231 11464
rect 19996 11460 20002 11462
rect 28165 11459 28231 11462
rect 5130 11456 5446 11457
rect 5130 11392 5136 11456
rect 5200 11392 5216 11456
rect 5280 11392 5296 11456
rect 5360 11392 5376 11456
rect 5440 11392 5446 11456
rect 5130 11391 5446 11392
rect 35850 11456 36166 11457
rect 35850 11392 35856 11456
rect 35920 11392 35936 11456
rect 36000 11392 36016 11456
rect 36080 11392 36096 11456
rect 36160 11392 36166 11456
rect 35850 11391 36166 11392
rect 66570 11456 66886 11457
rect 66570 11392 66576 11456
rect 66640 11392 66656 11456
rect 66720 11392 66736 11456
rect 66800 11392 66816 11456
rect 66880 11392 66886 11456
rect 66570 11391 66886 11392
rect 17718 11324 17724 11388
rect 17788 11386 17794 11388
rect 27981 11386 28047 11389
rect 17788 11384 28047 11386
rect 17788 11328 27986 11384
rect 28042 11328 28047 11384
rect 17788 11326 28047 11328
rect 17788 11324 17794 11326
rect 27981 11323 28047 11326
rect 15326 11188 15332 11252
rect 15396 11250 15402 11252
rect 22461 11250 22527 11253
rect 15396 11248 22527 11250
rect 15396 11192 22466 11248
rect 22522 11192 22527 11248
rect 15396 11190 22527 11192
rect 15396 11188 15402 11190
rect 22461 11187 22527 11190
rect 13302 11052 13308 11116
rect 13372 11114 13378 11116
rect 23473 11114 23539 11117
rect 13372 11112 23539 11114
rect 13372 11056 23478 11112
rect 23534 11056 23539 11112
rect 13372 11054 23539 11056
rect 13372 11052 13378 11054
rect 23473 11051 23539 11054
rect 24945 11114 25011 11117
rect 26550 11114 26556 11116
rect 24945 11112 26556 11114
rect 24945 11056 24950 11112
rect 25006 11056 26556 11112
rect 24945 11054 26556 11056
rect 24945 11051 25011 11054
rect 26550 11052 26556 11054
rect 26620 11052 26626 11116
rect 21633 10978 21699 10981
rect 28165 10978 28231 10981
rect 21633 10976 28231 10978
rect 21633 10920 21638 10976
rect 21694 10920 28170 10976
rect 28226 10920 28231 10976
rect 21633 10918 28231 10920
rect 21633 10915 21699 10918
rect 28165 10915 28231 10918
rect 5790 10912 6106 10913
rect 5790 10848 5796 10912
rect 5860 10848 5876 10912
rect 5940 10848 5956 10912
rect 6020 10848 6036 10912
rect 6100 10848 6106 10912
rect 5790 10847 6106 10848
rect 36510 10912 36826 10913
rect 36510 10848 36516 10912
rect 36580 10848 36596 10912
rect 36660 10848 36676 10912
rect 36740 10848 36756 10912
rect 36820 10848 36826 10912
rect 36510 10847 36826 10848
rect 67230 10912 67546 10913
rect 67230 10848 67236 10912
rect 67300 10848 67316 10912
rect 67380 10848 67396 10912
rect 67460 10848 67476 10912
rect 67540 10848 67546 10912
rect 67230 10847 67546 10848
rect 17350 10780 17356 10844
rect 17420 10842 17426 10844
rect 28809 10842 28875 10845
rect 17420 10840 28875 10842
rect 17420 10784 28814 10840
rect 28870 10784 28875 10840
rect 17420 10782 28875 10784
rect 17420 10780 17426 10782
rect 28809 10779 28875 10782
rect 10726 10644 10732 10708
rect 10796 10706 10802 10708
rect 31201 10706 31267 10709
rect 10796 10704 31267 10706
rect 10796 10648 31206 10704
rect 31262 10648 31267 10704
rect 10796 10646 31267 10648
rect 10796 10644 10802 10646
rect 31201 10643 31267 10646
rect 19977 10570 20043 10573
rect 23381 10570 23447 10573
rect 19977 10568 23447 10570
rect 19977 10512 19982 10568
rect 20038 10512 23386 10568
rect 23442 10512 23447 10568
rect 19977 10510 23447 10512
rect 19977 10507 20043 10510
rect 23381 10507 23447 10510
rect 24393 10570 24459 10573
rect 25773 10570 25839 10573
rect 26233 10572 26299 10573
rect 26182 10570 26188 10572
rect 24393 10568 25839 10570
rect 24393 10512 24398 10568
rect 24454 10512 25778 10568
rect 25834 10512 25839 10568
rect 24393 10510 25839 10512
rect 26142 10510 26188 10570
rect 26252 10568 26299 10572
rect 26294 10512 26299 10568
rect 24393 10507 24459 10510
rect 25773 10507 25839 10510
rect 26182 10508 26188 10510
rect 26252 10508 26299 10512
rect 26233 10507 26299 10508
rect 16430 10372 16436 10436
rect 16500 10434 16506 10436
rect 28625 10434 28691 10437
rect 16500 10432 28691 10434
rect 16500 10376 28630 10432
rect 28686 10376 28691 10432
rect 16500 10374 28691 10376
rect 16500 10372 16506 10374
rect 28625 10371 28691 10374
rect 29177 10434 29243 10437
rect 30966 10434 30972 10436
rect 29177 10432 30972 10434
rect 29177 10376 29182 10432
rect 29238 10376 30972 10432
rect 29177 10374 30972 10376
rect 29177 10371 29243 10374
rect 30966 10372 30972 10374
rect 31036 10372 31042 10436
rect 5130 10368 5446 10369
rect 5130 10304 5136 10368
rect 5200 10304 5216 10368
rect 5280 10304 5296 10368
rect 5360 10304 5376 10368
rect 5440 10304 5446 10368
rect 5130 10303 5446 10304
rect 35850 10368 36166 10369
rect 35850 10304 35856 10368
rect 35920 10304 35936 10368
rect 36000 10304 36016 10368
rect 36080 10304 36096 10368
rect 36160 10304 36166 10368
rect 35850 10303 36166 10304
rect 66570 10368 66886 10369
rect 66570 10304 66576 10368
rect 66640 10304 66656 10368
rect 66720 10304 66736 10368
rect 66800 10304 66816 10368
rect 66880 10304 66886 10368
rect 66570 10303 66886 10304
rect 10910 10236 10916 10300
rect 10980 10298 10986 10300
rect 21541 10298 21607 10301
rect 10980 10296 21607 10298
rect 10980 10240 21546 10296
rect 21602 10240 21607 10296
rect 10980 10238 21607 10240
rect 10980 10236 10986 10238
rect 21541 10235 21607 10238
rect 23054 10236 23060 10300
rect 23124 10298 23130 10300
rect 23124 10238 31770 10298
rect 23124 10236 23130 10238
rect 18086 10100 18092 10164
rect 18156 10162 18162 10164
rect 31201 10162 31267 10165
rect 18156 10160 31267 10162
rect 18156 10104 31206 10160
rect 31262 10104 31267 10160
rect 18156 10102 31267 10104
rect 31710 10162 31770 10238
rect 31845 10162 31911 10165
rect 31710 10160 31911 10162
rect 31710 10104 31850 10160
rect 31906 10104 31911 10160
rect 31710 10102 31911 10104
rect 18156 10100 18162 10102
rect 31201 10099 31267 10102
rect 31845 10099 31911 10102
rect 21357 10026 21423 10029
rect 21766 10026 21772 10028
rect 21357 10024 21772 10026
rect 21357 9968 21362 10024
rect 21418 9968 21772 10024
rect 21357 9966 21772 9968
rect 21357 9963 21423 9966
rect 21766 9964 21772 9966
rect 21836 9964 21842 10028
rect 22686 9964 22692 10028
rect 22756 10026 22762 10028
rect 23473 10026 23539 10029
rect 22756 10024 23539 10026
rect 22756 9968 23478 10024
rect 23534 9968 23539 10024
rect 22756 9966 23539 9968
rect 22756 9964 22762 9966
rect 23473 9963 23539 9966
rect 23790 9964 23796 10028
rect 23860 10026 23866 10028
rect 27981 10026 28047 10029
rect 23860 10024 28047 10026
rect 23860 9968 27986 10024
rect 28042 9968 28047 10024
rect 23860 9966 28047 9968
rect 23860 9964 23866 9966
rect 27981 9963 28047 9966
rect 9029 9890 9095 9893
rect 21357 9890 21423 9893
rect 9029 9888 21423 9890
rect 9029 9832 9034 9888
rect 9090 9832 21362 9888
rect 21418 9832 21423 9888
rect 9029 9830 21423 9832
rect 9029 9827 9095 9830
rect 21357 9827 21423 9830
rect 23381 9890 23447 9893
rect 23381 9888 23490 9890
rect 23381 9832 23386 9888
rect 23442 9832 23490 9888
rect 23381 9827 23490 9832
rect 5790 9824 6106 9825
rect 5790 9760 5796 9824
rect 5860 9760 5876 9824
rect 5940 9760 5956 9824
rect 6020 9760 6036 9824
rect 6100 9760 6106 9824
rect 5790 9759 6106 9760
rect 13537 9754 13603 9757
rect 23289 9754 23355 9757
rect 13537 9752 23355 9754
rect 13537 9696 13542 9752
rect 13598 9696 23294 9752
rect 23350 9696 23355 9752
rect 13537 9694 23355 9696
rect 13537 9691 13603 9694
rect 23289 9691 23355 9694
rect 19742 9556 19748 9620
rect 19812 9618 19818 9620
rect 22921 9618 22987 9621
rect 19812 9616 22987 9618
rect 19812 9560 22926 9616
rect 22982 9560 22987 9616
rect 19812 9558 22987 9560
rect 23430 9618 23490 9827
rect 36510 9824 36826 9825
rect 36510 9760 36516 9824
rect 36580 9760 36596 9824
rect 36660 9760 36676 9824
rect 36740 9760 36756 9824
rect 36820 9760 36826 9824
rect 36510 9759 36826 9760
rect 67230 9824 67546 9825
rect 67230 9760 67236 9824
rect 67300 9760 67316 9824
rect 67380 9760 67396 9824
rect 67460 9760 67476 9824
rect 67540 9760 67546 9824
rect 67230 9759 67546 9760
rect 24894 9692 24900 9756
rect 24964 9754 24970 9756
rect 25589 9754 25655 9757
rect 24964 9752 25655 9754
rect 24964 9696 25594 9752
rect 25650 9696 25655 9752
rect 24964 9694 25655 9696
rect 24964 9692 24970 9694
rect 25589 9691 25655 9694
rect 26969 9754 27035 9757
rect 30189 9756 30255 9757
rect 29126 9754 29132 9756
rect 26969 9752 29132 9754
rect 26969 9696 26974 9752
rect 27030 9696 29132 9752
rect 26969 9694 29132 9696
rect 26969 9691 27035 9694
rect 29126 9692 29132 9694
rect 29196 9692 29202 9756
rect 30189 9752 30236 9756
rect 30300 9754 30306 9756
rect 30189 9696 30194 9752
rect 30189 9692 30236 9696
rect 30300 9694 30346 9754
rect 30300 9692 30306 9694
rect 30189 9691 30255 9692
rect 28993 9620 29059 9621
rect 23430 9558 25330 9618
rect 19812 9556 19818 9558
rect 22921 9555 22987 9558
rect 15653 9482 15719 9485
rect 24669 9482 24735 9485
rect 15653 9480 24735 9482
rect 15653 9424 15658 9480
rect 15714 9424 24674 9480
rect 24730 9424 24735 9480
rect 15653 9422 24735 9424
rect 15653 9419 15719 9422
rect 24669 9419 24735 9422
rect 13445 9346 13511 9349
rect 23381 9346 23447 9349
rect 13445 9344 23447 9346
rect 13445 9288 13450 9344
rect 13506 9288 23386 9344
rect 23442 9288 23447 9344
rect 13445 9286 23447 9288
rect 13445 9283 13511 9286
rect 23381 9283 23447 9286
rect 24158 9284 24164 9348
rect 24228 9346 24234 9348
rect 24485 9346 24551 9349
rect 24228 9344 24551 9346
rect 24228 9288 24490 9344
rect 24546 9288 24551 9344
rect 24228 9286 24551 9288
rect 25270 9346 25330 9558
rect 28942 9556 28948 9620
rect 29012 9618 29059 9620
rect 31845 9618 31911 9621
rect 33041 9618 33107 9621
rect 29012 9616 29104 9618
rect 29054 9560 29104 9616
rect 29012 9558 29104 9560
rect 31845 9616 33107 9618
rect 31845 9560 31850 9616
rect 31906 9560 33046 9616
rect 33102 9560 33107 9616
rect 31845 9558 33107 9560
rect 29012 9556 29059 9558
rect 28993 9555 29059 9556
rect 31845 9555 31911 9558
rect 33041 9555 33107 9558
rect 30557 9482 30623 9485
rect 33225 9482 33291 9485
rect 35709 9482 35775 9485
rect 30557 9480 35775 9482
rect 30557 9424 30562 9480
rect 30618 9424 33230 9480
rect 33286 9424 35714 9480
rect 35770 9424 35775 9480
rect 30557 9422 35775 9424
rect 30557 9419 30623 9422
rect 33225 9419 33291 9422
rect 35709 9419 35775 9422
rect 33685 9346 33751 9349
rect 25270 9344 33751 9346
rect 25270 9288 33690 9344
rect 33746 9288 33751 9344
rect 25270 9286 33751 9288
rect 24228 9284 24234 9286
rect 24485 9283 24551 9286
rect 33685 9283 33751 9286
rect 5130 9280 5446 9281
rect 5130 9216 5136 9280
rect 5200 9216 5216 9280
rect 5280 9216 5296 9280
rect 5360 9216 5376 9280
rect 5440 9216 5446 9280
rect 5130 9215 5446 9216
rect 35850 9280 36166 9281
rect 35850 9216 35856 9280
rect 35920 9216 35936 9280
rect 36000 9216 36016 9280
rect 36080 9216 36096 9280
rect 36160 9216 36166 9280
rect 35850 9215 36166 9216
rect 66570 9280 66886 9281
rect 66570 9216 66576 9280
rect 66640 9216 66656 9280
rect 66720 9216 66736 9280
rect 66800 9216 66816 9280
rect 66880 9216 66886 9280
rect 66570 9215 66886 9216
rect 23565 9210 23631 9213
rect 12390 9208 23631 9210
rect 12390 9152 23570 9208
rect 23626 9152 23631 9208
rect 12390 9150 23631 9152
rect 11973 9074 12039 9077
rect 12390 9074 12450 9150
rect 23565 9147 23631 9150
rect 11973 9072 12450 9074
rect 11973 9016 11978 9072
rect 12034 9016 12450 9072
rect 11973 9014 12450 9016
rect 19333 9074 19399 9077
rect 19609 9074 19675 9077
rect 21265 9074 21331 9077
rect 19333 9072 21331 9074
rect 19333 9016 19338 9072
rect 19394 9016 19614 9072
rect 19670 9016 21270 9072
rect 21326 9016 21331 9072
rect 19333 9014 21331 9016
rect 11973 9011 12039 9014
rect 19333 9011 19399 9014
rect 19609 9011 19675 9014
rect 21265 9011 21331 9014
rect 24710 9012 24716 9076
rect 24780 9074 24786 9076
rect 28625 9074 28691 9077
rect 24780 9072 28691 9074
rect 24780 9016 28630 9072
rect 28686 9016 28691 9072
rect 24780 9014 28691 9016
rect 24780 9012 24786 9014
rect 28625 9011 28691 9014
rect 29310 9012 29316 9076
rect 29380 9074 29386 9076
rect 29637 9074 29703 9077
rect 29380 9072 29703 9074
rect 29380 9016 29642 9072
rect 29698 9016 29703 9072
rect 29380 9014 29703 9016
rect 29380 9012 29386 9014
rect 29637 9011 29703 9014
rect 10409 8938 10475 8941
rect 20437 8938 20503 8941
rect 10409 8936 20503 8938
rect 10409 8880 10414 8936
rect 10470 8880 20442 8936
rect 20498 8880 20503 8936
rect 10409 8878 20503 8880
rect 10409 8875 10475 8878
rect 20437 8875 20503 8878
rect 22829 8938 22895 8941
rect 27429 8938 27495 8941
rect 22829 8936 27495 8938
rect 22829 8880 22834 8936
rect 22890 8880 27434 8936
rect 27490 8880 27495 8936
rect 22829 8878 27495 8880
rect 22829 8875 22895 8878
rect 27429 8875 27495 8878
rect 28758 8876 28764 8940
rect 28828 8938 28834 8940
rect 37365 8938 37431 8941
rect 28828 8936 37431 8938
rect 28828 8880 37370 8936
rect 37426 8880 37431 8936
rect 28828 8878 37431 8880
rect 28828 8876 28834 8878
rect 37365 8875 37431 8878
rect 17902 8740 17908 8804
rect 17972 8802 17978 8804
rect 18229 8802 18295 8805
rect 17972 8800 18295 8802
rect 17972 8744 18234 8800
rect 18290 8744 18295 8800
rect 17972 8742 18295 8744
rect 17972 8740 17978 8742
rect 18229 8739 18295 8742
rect 18638 8740 18644 8804
rect 18708 8802 18714 8804
rect 27705 8802 27771 8805
rect 18708 8800 27771 8802
rect 18708 8744 27710 8800
rect 27766 8744 27771 8800
rect 18708 8742 27771 8744
rect 18708 8740 18714 8742
rect 27705 8739 27771 8742
rect 29177 8802 29243 8805
rect 33041 8802 33107 8805
rect 29177 8800 33107 8802
rect 29177 8744 29182 8800
rect 29238 8744 33046 8800
rect 33102 8744 33107 8800
rect 29177 8742 33107 8744
rect 29177 8739 29243 8742
rect 33041 8739 33107 8742
rect 5790 8736 6106 8737
rect 5790 8672 5796 8736
rect 5860 8672 5876 8736
rect 5940 8672 5956 8736
rect 6020 8672 6036 8736
rect 6100 8672 6106 8736
rect 5790 8671 6106 8672
rect 36510 8736 36826 8737
rect 36510 8672 36516 8736
rect 36580 8672 36596 8736
rect 36660 8672 36676 8736
rect 36740 8672 36756 8736
rect 36820 8672 36826 8736
rect 36510 8671 36826 8672
rect 67230 8736 67546 8737
rect 67230 8672 67236 8736
rect 67300 8672 67316 8736
rect 67380 8672 67396 8736
rect 67460 8672 67476 8736
rect 67540 8672 67546 8736
rect 67230 8671 67546 8672
rect 11697 8666 11763 8669
rect 19885 8666 19951 8669
rect 11697 8664 19951 8666
rect 11697 8608 11702 8664
rect 11758 8608 19890 8664
rect 19946 8608 19951 8664
rect 11697 8606 19951 8608
rect 11697 8603 11763 8606
rect 19885 8603 19951 8606
rect 26233 8666 26299 8669
rect 32213 8666 32279 8669
rect 33133 8666 33199 8669
rect 26233 8664 32279 8666
rect 26233 8608 26238 8664
rect 26294 8608 32218 8664
rect 32274 8608 32279 8664
rect 26233 8606 32279 8608
rect 26233 8603 26299 8606
rect 32213 8603 32279 8606
rect 32446 8664 33199 8666
rect 32446 8608 33138 8664
rect 33194 8608 33199 8664
rect 32446 8606 33199 8608
rect 18270 8468 18276 8532
rect 18340 8530 18346 8532
rect 18597 8530 18663 8533
rect 18340 8528 18663 8530
rect 18340 8472 18602 8528
rect 18658 8472 18663 8528
rect 18340 8470 18663 8472
rect 18340 8468 18346 8470
rect 18597 8467 18663 8470
rect 19374 8468 19380 8532
rect 19444 8530 19450 8532
rect 19977 8530 20043 8533
rect 24301 8530 24367 8533
rect 19444 8528 20043 8530
rect 19444 8472 19982 8528
rect 20038 8472 20043 8528
rect 19444 8470 20043 8472
rect 19444 8468 19450 8470
rect 19977 8467 20043 8470
rect 20118 8528 24367 8530
rect 20118 8472 24306 8528
rect 24362 8472 24367 8528
rect 20118 8470 24367 8472
rect 15745 8394 15811 8397
rect 15745 8392 18338 8394
rect 15745 8336 15750 8392
rect 15806 8336 18338 8392
rect 15745 8334 18338 8336
rect 15745 8331 15811 8334
rect 18278 8258 18338 8334
rect 18454 8332 18460 8396
rect 18524 8394 18530 8396
rect 18689 8394 18755 8397
rect 20118 8394 20178 8470
rect 24301 8467 24367 8470
rect 25037 8530 25103 8533
rect 25262 8530 25268 8532
rect 25037 8528 25268 8530
rect 25037 8472 25042 8528
rect 25098 8472 25268 8528
rect 25037 8470 25268 8472
rect 25037 8467 25103 8470
rect 25262 8468 25268 8470
rect 25332 8468 25338 8532
rect 26325 8530 26391 8533
rect 26877 8530 26943 8533
rect 26325 8528 26943 8530
rect 26325 8472 26330 8528
rect 26386 8472 26882 8528
rect 26938 8472 26943 8528
rect 26325 8470 26943 8472
rect 26325 8467 26391 8470
rect 26877 8467 26943 8470
rect 27061 8530 27127 8533
rect 30189 8530 30255 8533
rect 27061 8528 30255 8530
rect 27061 8472 27066 8528
rect 27122 8472 30194 8528
rect 30250 8472 30255 8528
rect 27061 8470 30255 8472
rect 27061 8467 27127 8470
rect 30189 8467 30255 8470
rect 31150 8468 31156 8532
rect 31220 8530 31226 8532
rect 32446 8530 32506 8606
rect 33133 8603 33199 8606
rect 31220 8470 32506 8530
rect 31220 8468 31226 8470
rect 33358 8468 33364 8532
rect 33428 8530 33434 8532
rect 35249 8530 35315 8533
rect 33428 8528 35315 8530
rect 33428 8472 35254 8528
rect 35310 8472 35315 8528
rect 33428 8470 35315 8472
rect 33428 8468 33434 8470
rect 35249 8467 35315 8470
rect 37038 8468 37044 8532
rect 37108 8530 37114 8532
rect 37181 8530 37247 8533
rect 37108 8528 37247 8530
rect 37108 8472 37186 8528
rect 37242 8472 37247 8528
rect 37108 8470 37247 8472
rect 37108 8468 37114 8470
rect 37181 8467 37247 8470
rect 18524 8392 18755 8394
rect 18524 8336 18694 8392
rect 18750 8336 18755 8392
rect 18524 8334 18755 8336
rect 18524 8332 18530 8334
rect 18689 8331 18755 8334
rect 18830 8334 20178 8394
rect 18830 8258 18890 8334
rect 20662 8332 20668 8396
rect 20732 8394 20738 8396
rect 21173 8394 21239 8397
rect 20732 8392 21239 8394
rect 20732 8336 21178 8392
rect 21234 8336 21239 8392
rect 20732 8334 21239 8336
rect 20732 8332 20738 8334
rect 21173 8331 21239 8334
rect 25497 8394 25563 8397
rect 25814 8394 25820 8396
rect 25497 8392 25820 8394
rect 25497 8336 25502 8392
rect 25558 8336 25820 8392
rect 25497 8334 25820 8336
rect 25497 8331 25563 8334
rect 25814 8332 25820 8334
rect 25884 8332 25890 8396
rect 27153 8394 27219 8397
rect 27470 8394 27476 8396
rect 27153 8392 27476 8394
rect 27153 8336 27158 8392
rect 27214 8336 27476 8392
rect 27153 8334 27476 8336
rect 27153 8331 27219 8334
rect 27470 8332 27476 8334
rect 27540 8332 27546 8396
rect 27705 8394 27771 8397
rect 31385 8394 31451 8397
rect 27705 8392 31451 8394
rect 27705 8336 27710 8392
rect 27766 8336 31390 8392
rect 31446 8336 31451 8392
rect 27705 8334 31451 8336
rect 27705 8331 27771 8334
rect 31385 8331 31451 8334
rect 31753 8394 31819 8397
rect 31886 8394 31892 8396
rect 31753 8392 31892 8394
rect 31753 8336 31758 8392
rect 31814 8336 31892 8392
rect 31753 8334 31892 8336
rect 31753 8331 31819 8334
rect 31886 8332 31892 8334
rect 31956 8332 31962 8396
rect 33174 8332 33180 8396
rect 33244 8394 33250 8396
rect 33317 8394 33383 8397
rect 33244 8392 33383 8394
rect 33244 8336 33322 8392
rect 33378 8336 33383 8392
rect 33244 8334 33383 8336
rect 33244 8332 33250 8334
rect 33317 8331 33383 8334
rect 33726 8332 33732 8396
rect 33796 8394 33802 8396
rect 38653 8394 38719 8397
rect 33796 8392 38719 8394
rect 33796 8336 38658 8392
rect 38714 8336 38719 8392
rect 33796 8334 38719 8336
rect 33796 8332 33802 8334
rect 38653 8331 38719 8334
rect 18278 8198 18890 8258
rect 20897 8258 20963 8261
rect 27521 8258 27587 8261
rect 20897 8256 27587 8258
rect 20897 8200 20902 8256
rect 20958 8200 27526 8256
rect 27582 8200 27587 8256
rect 20897 8198 27587 8200
rect 20897 8195 20963 8198
rect 27521 8195 27587 8198
rect 32397 8258 32463 8261
rect 34697 8258 34763 8261
rect 32397 8256 34763 8258
rect 32397 8200 32402 8256
rect 32458 8200 34702 8256
rect 34758 8200 34763 8256
rect 32397 8198 34763 8200
rect 32397 8195 32463 8198
rect 34697 8195 34763 8198
rect 5130 8192 5446 8193
rect 5130 8128 5136 8192
rect 5200 8128 5216 8192
rect 5280 8128 5296 8192
rect 5360 8128 5376 8192
rect 5440 8128 5446 8192
rect 5130 8127 5446 8128
rect 35850 8192 36166 8193
rect 35850 8128 35856 8192
rect 35920 8128 35936 8192
rect 36000 8128 36016 8192
rect 36080 8128 36096 8192
rect 36160 8128 36166 8192
rect 35850 8127 36166 8128
rect 66570 8192 66886 8193
rect 66570 8128 66576 8192
rect 66640 8128 66656 8192
rect 66720 8128 66736 8192
rect 66800 8128 66816 8192
rect 66880 8128 66886 8192
rect 66570 8127 66886 8128
rect 17166 8060 17172 8124
rect 17236 8122 17242 8124
rect 24485 8122 24551 8125
rect 17236 8120 24551 8122
rect 17236 8064 24490 8120
rect 24546 8064 24551 8120
rect 17236 8062 24551 8064
rect 17236 8060 17242 8062
rect 24485 8059 24551 8062
rect 27153 8122 27219 8125
rect 30649 8122 30715 8125
rect 31385 8122 31451 8125
rect 27153 8120 31451 8122
rect 27153 8064 27158 8120
rect 27214 8064 30654 8120
rect 30710 8064 31390 8120
rect 31446 8064 31451 8120
rect 27153 8062 31451 8064
rect 27153 8059 27219 8062
rect 30649 8059 30715 8062
rect 31385 8059 31451 8062
rect 33133 8122 33199 8125
rect 33869 8122 33935 8125
rect 33133 8120 33935 8122
rect 33133 8064 33138 8120
rect 33194 8064 33874 8120
rect 33930 8064 33935 8120
rect 33133 8062 33935 8064
rect 33133 8059 33199 8062
rect 33869 8059 33935 8062
rect 20069 7986 20135 7989
rect 22553 7986 22619 7989
rect 24117 7986 24183 7989
rect 24894 7986 24900 7988
rect 20069 7984 24900 7986
rect 20069 7928 20074 7984
rect 20130 7928 22558 7984
rect 22614 7928 24122 7984
rect 24178 7928 24900 7984
rect 20069 7926 24900 7928
rect 20069 7923 20135 7926
rect 22553 7923 22619 7926
rect 24117 7923 24183 7926
rect 24894 7924 24900 7926
rect 24964 7924 24970 7988
rect 27613 7986 27679 7989
rect 28206 7986 28212 7988
rect 27613 7984 28212 7986
rect 27613 7928 27618 7984
rect 27674 7928 28212 7984
rect 27613 7926 28212 7928
rect 27613 7923 27679 7926
rect 28206 7924 28212 7926
rect 28276 7986 28282 7988
rect 28625 7986 28691 7989
rect 28276 7984 28691 7986
rect 28276 7928 28630 7984
rect 28686 7928 28691 7984
rect 28276 7926 28691 7928
rect 28276 7924 28282 7926
rect 28625 7923 28691 7926
rect 31477 7986 31543 7989
rect 31661 7986 31727 7989
rect 31477 7984 31727 7986
rect 31477 7928 31482 7984
rect 31538 7928 31666 7984
rect 31722 7928 31727 7984
rect 31477 7926 31727 7928
rect 31477 7923 31543 7926
rect 31661 7923 31727 7926
rect 33542 7924 33548 7988
rect 33612 7986 33618 7988
rect 38193 7986 38259 7989
rect 33612 7984 38259 7986
rect 33612 7928 38198 7984
rect 38254 7928 38259 7984
rect 33612 7926 38259 7928
rect 33612 7924 33618 7926
rect 38193 7923 38259 7926
rect 20110 7788 20116 7852
rect 20180 7850 20186 7852
rect 28165 7850 28231 7853
rect 30649 7852 30715 7853
rect 20180 7848 28231 7850
rect 20180 7792 28170 7848
rect 28226 7792 28231 7848
rect 20180 7790 28231 7792
rect 20180 7788 20186 7790
rect 28165 7787 28231 7790
rect 30598 7788 30604 7852
rect 30668 7850 30715 7852
rect 31753 7850 31819 7853
rect 32305 7852 32371 7853
rect 32254 7850 32260 7852
rect 30668 7848 31819 7850
rect 30710 7792 31758 7848
rect 31814 7792 31819 7848
rect 30668 7790 31819 7792
rect 32214 7790 32260 7850
rect 32324 7848 32371 7852
rect 32366 7792 32371 7848
rect 30668 7788 30715 7790
rect 30649 7787 30715 7788
rect 31753 7787 31819 7790
rect 32254 7788 32260 7790
rect 32324 7788 32371 7792
rect 32305 7787 32371 7788
rect 13670 7652 13676 7716
rect 13740 7714 13746 7716
rect 23473 7714 23539 7717
rect 13740 7712 23539 7714
rect 13740 7656 23478 7712
rect 23534 7656 23539 7712
rect 13740 7654 23539 7656
rect 13740 7652 13746 7654
rect 23473 7651 23539 7654
rect 23933 7714 23999 7717
rect 26969 7714 27035 7717
rect 23933 7712 27035 7714
rect 23933 7656 23938 7712
rect 23994 7656 26974 7712
rect 27030 7656 27035 7712
rect 23933 7654 27035 7656
rect 23933 7651 23999 7654
rect 26969 7651 27035 7654
rect 27102 7652 27108 7716
rect 27172 7714 27178 7716
rect 27429 7714 27495 7717
rect 27172 7712 27495 7714
rect 27172 7656 27434 7712
rect 27490 7656 27495 7712
rect 27172 7654 27495 7656
rect 27172 7652 27178 7654
rect 27429 7651 27495 7654
rect 31661 7714 31727 7717
rect 32305 7714 32371 7717
rect 31661 7712 32371 7714
rect 31661 7656 31666 7712
rect 31722 7656 32310 7712
rect 32366 7656 32371 7712
rect 31661 7654 32371 7656
rect 31661 7651 31727 7654
rect 32305 7651 32371 7654
rect 34462 7652 34468 7716
rect 34532 7714 34538 7716
rect 36261 7714 36327 7717
rect 34532 7712 36327 7714
rect 34532 7656 36266 7712
rect 36322 7656 36327 7712
rect 34532 7654 36327 7656
rect 34532 7652 34538 7654
rect 36261 7651 36327 7654
rect 5790 7648 6106 7649
rect 5790 7584 5796 7648
rect 5860 7584 5876 7648
rect 5940 7584 5956 7648
rect 6020 7584 6036 7648
rect 6100 7584 6106 7648
rect 5790 7583 6106 7584
rect 36510 7648 36826 7649
rect 36510 7584 36516 7648
rect 36580 7584 36596 7648
rect 36660 7584 36676 7648
rect 36740 7584 36756 7648
rect 36820 7584 36826 7648
rect 36510 7583 36826 7584
rect 67230 7648 67546 7649
rect 67230 7584 67236 7648
rect 67300 7584 67316 7648
rect 67380 7584 67396 7648
rect 67460 7584 67476 7648
rect 67540 7584 67546 7648
rect 67230 7583 67546 7584
rect 9673 7578 9739 7581
rect 21449 7578 21515 7581
rect 9673 7576 21515 7578
rect 9673 7520 9678 7576
rect 9734 7520 21454 7576
rect 21510 7520 21515 7576
rect 9673 7518 21515 7520
rect 9673 7515 9739 7518
rect 21449 7515 21515 7518
rect 21725 7578 21791 7581
rect 25037 7578 25103 7581
rect 21725 7576 25103 7578
rect 21725 7520 21730 7576
rect 21786 7520 25042 7576
rect 25098 7520 25103 7576
rect 21725 7518 25103 7520
rect 21725 7515 21791 7518
rect 25037 7515 25103 7518
rect 27286 7516 27292 7580
rect 27356 7578 27362 7580
rect 27521 7578 27587 7581
rect 33777 7578 33843 7581
rect 35985 7578 36051 7581
rect 27356 7576 36051 7578
rect 27356 7520 27526 7576
rect 27582 7520 33782 7576
rect 33838 7520 35990 7576
rect 36046 7520 36051 7576
rect 27356 7518 36051 7520
rect 27356 7516 27362 7518
rect 27521 7515 27587 7518
rect 33777 7515 33843 7518
rect 35985 7515 36051 7518
rect 22369 7442 22435 7445
rect 22829 7442 22895 7445
rect 22369 7440 22895 7442
rect 22369 7384 22374 7440
rect 22430 7384 22834 7440
rect 22890 7384 22895 7440
rect 22369 7382 22895 7384
rect 22369 7379 22435 7382
rect 22829 7379 22895 7382
rect 23422 7380 23428 7444
rect 23492 7442 23498 7444
rect 27153 7442 27219 7445
rect 23492 7440 27219 7442
rect 23492 7384 27158 7440
rect 27214 7384 27219 7440
rect 23492 7382 27219 7384
rect 23492 7380 23498 7382
rect 27153 7379 27219 7382
rect 29545 7442 29611 7445
rect 31937 7442 32003 7445
rect 29545 7440 32003 7442
rect 29545 7384 29550 7440
rect 29606 7384 31942 7440
rect 31998 7384 32003 7440
rect 29545 7382 32003 7384
rect 29545 7379 29611 7382
rect 31937 7379 32003 7382
rect 19425 7306 19491 7309
rect 21214 7306 21220 7308
rect 19425 7304 21220 7306
rect 19425 7248 19430 7304
rect 19486 7248 21220 7304
rect 19425 7246 21220 7248
rect 19425 7243 19491 7246
rect 21214 7244 21220 7246
rect 21284 7244 21290 7308
rect 22001 7306 22067 7309
rect 28073 7306 28139 7309
rect 22001 7304 28139 7306
rect 22001 7248 22006 7304
rect 22062 7248 28078 7304
rect 28134 7248 28139 7304
rect 22001 7246 28139 7248
rect 22001 7243 22067 7246
rect 28073 7243 28139 7246
rect 30097 7306 30163 7309
rect 32213 7306 32279 7309
rect 32806 7306 32812 7308
rect 30097 7304 32812 7306
rect 30097 7248 30102 7304
rect 30158 7248 32218 7304
rect 32274 7248 32812 7304
rect 30097 7246 32812 7248
rect 30097 7243 30163 7246
rect 32213 7243 32279 7246
rect 32806 7244 32812 7246
rect 32876 7244 32882 7308
rect 27153 7170 27219 7173
rect 27286 7170 27292 7172
rect 27153 7168 27292 7170
rect 27153 7112 27158 7168
rect 27214 7112 27292 7168
rect 27153 7110 27292 7112
rect 27153 7107 27219 7110
rect 27286 7108 27292 7110
rect 27356 7170 27362 7172
rect 27356 7110 29010 7170
rect 27356 7108 27362 7110
rect 5130 7104 5446 7105
rect 5130 7040 5136 7104
rect 5200 7040 5216 7104
rect 5280 7040 5296 7104
rect 5360 7040 5376 7104
rect 5440 7040 5446 7104
rect 5130 7039 5446 7040
rect 20897 7034 20963 7037
rect 16438 7032 20963 7034
rect 16438 6976 20902 7032
rect 20958 6976 20963 7032
rect 16438 6974 20963 6976
rect 15653 6898 15719 6901
rect 15837 6898 15903 6901
rect 15653 6896 15903 6898
rect 15653 6840 15658 6896
rect 15714 6840 15842 6896
rect 15898 6840 15903 6896
rect 15653 6838 15903 6840
rect 15653 6835 15719 6838
rect 15837 6835 15903 6838
rect 5790 6560 6106 6561
rect 5790 6496 5796 6560
rect 5860 6496 5876 6560
rect 5940 6496 5956 6560
rect 6020 6496 6036 6560
rect 6100 6496 6106 6560
rect 5790 6495 6106 6496
rect 12709 6354 12775 6357
rect 15561 6354 15627 6357
rect 12709 6352 15627 6354
rect 12709 6296 12714 6352
rect 12770 6296 15566 6352
rect 15622 6296 15627 6352
rect 12709 6294 15627 6296
rect 12709 6291 12775 6294
rect 15561 6291 15627 6294
rect 16113 6354 16179 6357
rect 16438 6354 16498 6974
rect 20897 6971 20963 6974
rect 22553 7034 22619 7037
rect 26785 7034 26851 7037
rect 22553 7032 26851 7034
rect 22553 6976 22558 7032
rect 22614 6976 26790 7032
rect 26846 6976 26851 7032
rect 22553 6974 26851 6976
rect 28950 7034 29010 7110
rect 35850 7104 36166 7105
rect 35850 7040 35856 7104
rect 35920 7040 35936 7104
rect 36000 7040 36016 7104
rect 36080 7040 36096 7104
rect 36160 7040 36166 7104
rect 35850 7039 36166 7040
rect 66570 7104 66886 7105
rect 66570 7040 66576 7104
rect 66640 7040 66656 7104
rect 66720 7040 66736 7104
rect 66800 7040 66816 7104
rect 66880 7040 66886 7104
rect 66570 7039 66886 7040
rect 30649 7034 30715 7037
rect 31845 7034 31911 7037
rect 32305 7034 32371 7037
rect 28950 7032 32371 7034
rect 28950 6976 30654 7032
rect 30710 6976 31850 7032
rect 31906 6976 32310 7032
rect 32366 6976 32371 7032
rect 28950 6974 32371 6976
rect 22553 6971 22619 6974
rect 26785 6971 26851 6974
rect 30649 6971 30715 6974
rect 31845 6971 31911 6974
rect 32305 6971 32371 6974
rect 20713 6898 20779 6901
rect 22369 6898 22435 6901
rect 20713 6896 22435 6898
rect 20713 6840 20718 6896
rect 20774 6840 22374 6896
rect 22430 6840 22435 6896
rect 20713 6838 22435 6840
rect 20713 6835 20779 6838
rect 22369 6835 22435 6838
rect 22737 6898 22803 6901
rect 25313 6898 25379 6901
rect 22737 6896 25379 6898
rect 22737 6840 22742 6896
rect 22798 6840 25318 6896
rect 25374 6840 25379 6896
rect 22737 6838 25379 6840
rect 22737 6835 22803 6838
rect 25313 6835 25379 6838
rect 30966 6836 30972 6900
rect 31036 6898 31042 6900
rect 31109 6898 31175 6901
rect 31036 6896 31175 6898
rect 31036 6840 31114 6896
rect 31170 6840 31175 6896
rect 31036 6838 31175 6840
rect 31036 6836 31042 6838
rect 31109 6835 31175 6838
rect 34881 6898 34947 6901
rect 35014 6898 35020 6900
rect 34881 6896 35020 6898
rect 34881 6840 34886 6896
rect 34942 6840 35020 6896
rect 34881 6838 35020 6840
rect 34881 6835 34947 6838
rect 35014 6836 35020 6838
rect 35084 6898 35090 6900
rect 39389 6898 39455 6901
rect 35084 6896 39455 6898
rect 35084 6840 39394 6896
rect 39450 6840 39455 6896
rect 35084 6838 39455 6840
rect 35084 6836 35090 6838
rect 39389 6835 39455 6838
rect 19609 6762 19675 6765
rect 22185 6762 22251 6765
rect 19609 6760 22251 6762
rect 19609 6704 19614 6760
rect 19670 6704 22190 6760
rect 22246 6704 22251 6760
rect 19609 6702 22251 6704
rect 19609 6699 19675 6702
rect 22185 6699 22251 6702
rect 22369 6762 22435 6765
rect 30097 6762 30163 6765
rect 22369 6760 30163 6762
rect 22369 6704 22374 6760
rect 22430 6704 30102 6760
rect 30158 6704 30163 6760
rect 22369 6702 30163 6704
rect 22369 6699 22435 6702
rect 30097 6699 30163 6702
rect 35157 6762 35223 6765
rect 35801 6762 35867 6765
rect 38101 6762 38167 6765
rect 35157 6760 38167 6762
rect 35157 6704 35162 6760
rect 35218 6704 35806 6760
rect 35862 6704 38106 6760
rect 38162 6704 38167 6760
rect 35157 6702 38167 6704
rect 35157 6699 35223 6702
rect 35801 6699 35867 6702
rect 38101 6699 38167 6702
rect 21817 6626 21883 6629
rect 27981 6626 28047 6629
rect 21817 6624 28047 6626
rect 21817 6568 21822 6624
rect 21878 6568 27986 6624
rect 28042 6568 28047 6624
rect 21817 6566 28047 6568
rect 21817 6563 21883 6566
rect 27981 6563 28047 6566
rect 30097 6626 30163 6629
rect 33317 6626 33383 6629
rect 30097 6624 33383 6626
rect 30097 6568 30102 6624
rect 30158 6568 33322 6624
rect 33378 6568 33383 6624
rect 30097 6566 33383 6568
rect 30097 6563 30163 6566
rect 33317 6563 33383 6566
rect 34329 6626 34395 6629
rect 35893 6626 35959 6629
rect 34329 6624 35959 6626
rect 34329 6568 34334 6624
rect 34390 6568 35898 6624
rect 35954 6568 35959 6624
rect 34329 6566 35959 6568
rect 34329 6563 34395 6566
rect 35893 6563 35959 6566
rect 38561 6626 38627 6629
rect 38561 6624 38670 6626
rect 38561 6568 38566 6624
rect 38622 6568 38670 6624
rect 38561 6563 38670 6568
rect 36510 6560 36826 6561
rect 36510 6496 36516 6560
rect 36580 6496 36596 6560
rect 36660 6496 36676 6560
rect 36740 6496 36756 6560
rect 36820 6496 36826 6560
rect 36510 6495 36826 6496
rect 22001 6490 22067 6493
rect 22134 6490 22140 6492
rect 22001 6488 22140 6490
rect 22001 6432 22006 6488
rect 22062 6432 22140 6488
rect 22001 6430 22140 6432
rect 22001 6427 22067 6430
rect 22134 6428 22140 6430
rect 22204 6428 22210 6492
rect 22277 6490 22343 6493
rect 26233 6490 26299 6493
rect 28625 6490 28691 6493
rect 22277 6488 28691 6490
rect 22277 6432 22282 6488
rect 22338 6432 26238 6488
rect 26294 6432 28630 6488
rect 28686 6432 28691 6488
rect 22277 6430 28691 6432
rect 22277 6427 22343 6430
rect 26233 6427 26299 6430
rect 28625 6427 28691 6430
rect 30925 6488 30991 6493
rect 30925 6432 30930 6488
rect 30986 6432 30991 6488
rect 30925 6427 30991 6432
rect 32397 6490 32463 6493
rect 33777 6490 33843 6493
rect 32397 6488 33843 6490
rect 32397 6432 32402 6488
rect 32458 6432 33782 6488
rect 33838 6432 33843 6488
rect 32397 6430 33843 6432
rect 32397 6427 32463 6430
rect 33777 6427 33843 6430
rect 37825 6490 37891 6493
rect 38469 6490 38535 6493
rect 37825 6488 38535 6490
rect 37825 6432 37830 6488
rect 37886 6432 38474 6488
rect 38530 6432 38535 6488
rect 37825 6430 38535 6432
rect 37825 6427 37891 6430
rect 38469 6427 38535 6430
rect 16113 6352 16498 6354
rect 16113 6296 16118 6352
rect 16174 6296 16498 6352
rect 16113 6294 16498 6296
rect 19241 6354 19307 6357
rect 26509 6354 26575 6357
rect 19241 6352 26575 6354
rect 19241 6296 19246 6352
rect 19302 6296 26514 6352
rect 26570 6296 26575 6352
rect 19241 6294 26575 6296
rect 16113 6291 16179 6294
rect 19241 6291 19307 6294
rect 26509 6291 26575 6294
rect 30928 6221 30988 6427
rect 10133 6218 10199 6221
rect 17166 6218 17172 6220
rect 10133 6216 17172 6218
rect 10133 6160 10138 6216
rect 10194 6160 17172 6216
rect 10133 6158 17172 6160
rect 10133 6155 10199 6158
rect 17166 6156 17172 6158
rect 17236 6156 17242 6220
rect 19333 6218 19399 6221
rect 28441 6218 28507 6221
rect 19333 6216 28507 6218
rect 19333 6160 19338 6216
rect 19394 6160 28446 6216
rect 28502 6160 28507 6216
rect 19333 6158 28507 6160
rect 19333 6155 19399 6158
rect 28441 6155 28507 6158
rect 30925 6216 30991 6221
rect 30925 6160 30930 6216
rect 30986 6160 30991 6216
rect 30925 6155 30991 6160
rect 31201 6218 31267 6221
rect 31661 6218 31727 6221
rect 33041 6218 33107 6221
rect 31201 6216 33107 6218
rect 31201 6160 31206 6216
rect 31262 6160 31666 6216
rect 31722 6160 33046 6216
rect 33102 6160 33107 6216
rect 31201 6158 33107 6160
rect 31201 6155 31267 6158
rect 31661 6155 31727 6158
rect 33041 6155 33107 6158
rect 35157 6218 35223 6221
rect 37825 6218 37891 6221
rect 35157 6216 37891 6218
rect 35157 6160 35162 6216
rect 35218 6160 37830 6216
rect 37886 6160 37891 6216
rect 35157 6158 37891 6160
rect 35157 6155 35223 6158
rect 37825 6155 37891 6158
rect 38469 6218 38535 6221
rect 38610 6218 38670 6563
rect 67230 6560 67546 6561
rect 67230 6496 67236 6560
rect 67300 6496 67316 6560
rect 67380 6496 67396 6560
rect 67460 6496 67476 6560
rect 67540 6496 67546 6560
rect 67230 6495 67546 6496
rect 38929 6354 38995 6357
rect 39481 6354 39547 6357
rect 38929 6352 39547 6354
rect 38929 6296 38934 6352
rect 38990 6296 39486 6352
rect 39542 6296 39547 6352
rect 38929 6294 39547 6296
rect 38929 6291 38995 6294
rect 39481 6291 39547 6294
rect 38469 6216 38670 6218
rect 38469 6160 38474 6216
rect 38530 6160 38670 6216
rect 38469 6158 38670 6160
rect 38469 6155 38535 6158
rect 12709 6082 12775 6085
rect 16389 6084 16455 6085
rect 18597 6084 18663 6085
rect 16062 6082 16068 6084
rect 12709 6080 16068 6082
rect 12709 6024 12714 6080
rect 12770 6024 16068 6080
rect 12709 6022 16068 6024
rect 12709 6019 12775 6022
rect 16062 6020 16068 6022
rect 16132 6020 16138 6084
rect 16389 6082 16436 6084
rect 16344 6080 16436 6082
rect 16344 6024 16394 6080
rect 16344 6022 16436 6024
rect 16389 6020 16436 6022
rect 16500 6020 16506 6084
rect 16982 6020 16988 6084
rect 17052 6082 17058 6084
rect 18086 6082 18092 6084
rect 17052 6022 18092 6082
rect 17052 6020 17058 6022
rect 18086 6020 18092 6022
rect 18156 6020 18162 6084
rect 18597 6082 18644 6084
rect 18552 6080 18644 6082
rect 18552 6024 18602 6080
rect 18552 6022 18644 6024
rect 18597 6020 18644 6022
rect 18708 6020 18714 6084
rect 28574 6020 28580 6084
rect 28644 6082 28650 6084
rect 32121 6082 32187 6085
rect 35709 6082 35775 6085
rect 28644 6022 31954 6082
rect 28644 6020 28650 6022
rect 16389 6019 16455 6020
rect 18597 6019 18663 6020
rect 5130 6016 5446 6017
rect 5130 5952 5136 6016
rect 5200 5952 5216 6016
rect 5280 5952 5296 6016
rect 5360 5952 5376 6016
rect 5440 5952 5446 6016
rect 5130 5951 5446 5952
rect 14089 5946 14155 5949
rect 23749 5948 23815 5949
rect 20662 5946 20668 5948
rect 14089 5944 20668 5946
rect 14089 5888 14094 5944
rect 14150 5888 20668 5944
rect 14089 5886 20668 5888
rect 14089 5883 14155 5886
rect 20662 5884 20668 5886
rect 20732 5884 20738 5948
rect 23749 5946 23796 5948
rect 23704 5944 23796 5946
rect 23704 5888 23754 5944
rect 23704 5886 23796 5888
rect 23749 5884 23796 5886
rect 23860 5884 23866 5948
rect 28257 5946 28323 5949
rect 28390 5946 28396 5948
rect 28257 5944 28396 5946
rect 28257 5888 28262 5944
rect 28318 5888 28396 5944
rect 28257 5886 28396 5888
rect 23749 5883 23815 5884
rect 28257 5883 28323 5886
rect 28390 5884 28396 5886
rect 28460 5946 28466 5948
rect 31894 5946 31954 6022
rect 32121 6080 35775 6082
rect 32121 6024 32126 6080
rect 32182 6024 35714 6080
rect 35770 6024 35775 6080
rect 32121 6022 35775 6024
rect 32121 6019 32187 6022
rect 35709 6019 35775 6022
rect 35850 6016 36166 6017
rect 35850 5952 35856 6016
rect 35920 5952 35936 6016
rect 36000 5952 36016 6016
rect 36080 5952 36096 6016
rect 36160 5952 36166 6016
rect 35850 5951 36166 5952
rect 66570 6016 66886 6017
rect 66570 5952 66576 6016
rect 66640 5952 66656 6016
rect 66720 5952 66736 6016
rect 66800 5952 66816 6016
rect 66880 5952 66886 6016
rect 66570 5951 66886 5952
rect 32213 5946 32279 5949
rect 28460 5886 31770 5946
rect 31894 5944 32279 5946
rect 31894 5888 32218 5944
rect 32274 5888 32279 5944
rect 31894 5886 32279 5888
rect 28460 5884 28466 5886
rect 31710 5813 31770 5886
rect 32213 5883 32279 5886
rect 36445 5946 36511 5949
rect 38561 5946 38627 5949
rect 36445 5944 38627 5946
rect 36445 5888 36450 5944
rect 36506 5888 38566 5944
rect 38622 5888 38627 5944
rect 36445 5886 38627 5888
rect 36445 5883 36511 5886
rect 38561 5883 38627 5886
rect 16297 5810 16363 5813
rect 19190 5810 19196 5812
rect 16297 5808 19196 5810
rect 16297 5752 16302 5808
rect 16358 5752 19196 5808
rect 16297 5750 19196 5752
rect 16297 5747 16363 5750
rect 19190 5748 19196 5750
rect 19260 5748 19266 5812
rect 19425 5810 19491 5813
rect 19926 5810 19932 5812
rect 19425 5808 19932 5810
rect 19425 5752 19430 5808
rect 19486 5752 19932 5808
rect 19425 5750 19932 5752
rect 19425 5747 19491 5750
rect 19926 5748 19932 5750
rect 19996 5748 20002 5812
rect 21214 5748 21220 5812
rect 21284 5810 21290 5812
rect 21357 5810 21423 5813
rect 21284 5808 21423 5810
rect 21284 5752 21362 5808
rect 21418 5752 21423 5808
rect 21284 5750 21423 5752
rect 21284 5748 21290 5750
rect 21357 5747 21423 5750
rect 25681 5810 25747 5813
rect 29085 5810 29151 5813
rect 25681 5808 29151 5810
rect 25681 5752 25686 5808
rect 25742 5752 29090 5808
rect 29146 5752 29151 5808
rect 25681 5750 29151 5752
rect 25681 5747 25747 5750
rect 29085 5747 29151 5750
rect 31661 5810 31770 5813
rect 40217 5810 40283 5813
rect 31661 5808 40283 5810
rect 31661 5752 31666 5808
rect 31722 5752 40222 5808
rect 40278 5752 40283 5808
rect 31661 5750 40283 5752
rect 31661 5747 31727 5750
rect 40217 5747 40283 5750
rect 12157 5674 12223 5677
rect 15101 5674 15167 5677
rect 12157 5672 15167 5674
rect 12157 5616 12162 5672
rect 12218 5616 15106 5672
rect 15162 5616 15167 5672
rect 12157 5614 15167 5616
rect 12157 5611 12223 5614
rect 15101 5611 15167 5614
rect 15285 5674 15351 5677
rect 22686 5674 22692 5676
rect 15285 5672 22692 5674
rect 15285 5616 15290 5672
rect 15346 5616 22692 5672
rect 15285 5614 22692 5616
rect 15285 5611 15351 5614
rect 22686 5612 22692 5614
rect 22756 5612 22762 5676
rect 23749 5674 23815 5677
rect 30557 5674 30623 5677
rect 32121 5674 32187 5677
rect 33961 5674 34027 5677
rect 23749 5672 29010 5674
rect 23749 5616 23754 5672
rect 23810 5616 29010 5672
rect 23749 5614 29010 5616
rect 23749 5611 23815 5614
rect 18597 5538 18663 5541
rect 24158 5538 24164 5540
rect 18597 5536 24164 5538
rect 18597 5480 18602 5536
rect 18658 5480 24164 5536
rect 18597 5478 24164 5480
rect 18597 5475 18663 5478
rect 24158 5476 24164 5478
rect 24228 5476 24234 5540
rect 27470 5476 27476 5540
rect 27540 5538 27546 5540
rect 27705 5538 27771 5541
rect 27540 5536 27771 5538
rect 27540 5480 27710 5536
rect 27766 5480 27771 5536
rect 27540 5478 27771 5480
rect 28950 5538 29010 5614
rect 30557 5672 32187 5674
rect 30557 5616 30562 5672
rect 30618 5616 32126 5672
rect 32182 5616 32187 5672
rect 30557 5614 32187 5616
rect 30557 5611 30623 5614
rect 32121 5611 32187 5614
rect 32446 5672 34027 5674
rect 32446 5616 33966 5672
rect 34022 5616 34027 5672
rect 32446 5614 34027 5616
rect 29637 5538 29703 5541
rect 28950 5536 29703 5538
rect 28950 5480 29642 5536
rect 29698 5480 29703 5536
rect 28950 5478 29703 5480
rect 27540 5476 27546 5478
rect 27705 5475 27771 5478
rect 29637 5475 29703 5478
rect 31845 5538 31911 5541
rect 32446 5538 32506 5614
rect 33961 5611 34027 5614
rect 34145 5674 34211 5677
rect 37273 5674 37339 5677
rect 34145 5672 37339 5674
rect 34145 5616 34150 5672
rect 34206 5616 37278 5672
rect 37334 5616 37339 5672
rect 34145 5614 37339 5616
rect 34145 5611 34211 5614
rect 37273 5611 37339 5614
rect 31845 5536 32506 5538
rect 31845 5480 31850 5536
rect 31906 5480 32506 5536
rect 31845 5478 32506 5480
rect 31845 5475 31911 5478
rect 5790 5472 6106 5473
rect 5790 5408 5796 5472
rect 5860 5408 5876 5472
rect 5940 5408 5956 5472
rect 6020 5408 6036 5472
rect 6100 5408 6106 5472
rect 5790 5407 6106 5408
rect 36510 5472 36826 5473
rect 36510 5408 36516 5472
rect 36580 5408 36596 5472
rect 36660 5408 36676 5472
rect 36740 5408 36756 5472
rect 36820 5408 36826 5472
rect 36510 5407 36826 5408
rect 67230 5472 67546 5473
rect 67230 5408 67236 5472
rect 67300 5408 67316 5472
rect 67380 5408 67396 5472
rect 67460 5408 67476 5472
rect 67540 5408 67546 5472
rect 67230 5407 67546 5408
rect 15193 5402 15259 5405
rect 15326 5402 15332 5404
rect 15193 5400 15332 5402
rect 15193 5344 15198 5400
rect 15254 5344 15332 5400
rect 15193 5342 15332 5344
rect 15193 5339 15259 5342
rect 15326 5340 15332 5342
rect 15396 5340 15402 5404
rect 19517 5402 19583 5405
rect 21449 5402 21515 5405
rect 22093 5402 22159 5405
rect 19517 5400 21515 5402
rect 19517 5344 19522 5400
rect 19578 5344 21454 5400
rect 21510 5344 21515 5400
rect 19517 5342 21515 5344
rect 19517 5339 19583 5342
rect 21449 5339 21515 5342
rect 21774 5400 22159 5402
rect 21774 5344 22098 5400
rect 22154 5344 22159 5400
rect 21774 5342 22159 5344
rect 13169 5266 13235 5269
rect 13302 5266 13308 5268
rect 13169 5264 13308 5266
rect 13169 5208 13174 5264
rect 13230 5208 13308 5264
rect 13169 5206 13308 5208
rect 13169 5203 13235 5206
rect 13302 5204 13308 5206
rect 13372 5204 13378 5268
rect 17677 5266 17743 5269
rect 20069 5266 20135 5269
rect 17677 5264 20135 5266
rect 17677 5208 17682 5264
rect 17738 5208 20074 5264
rect 20130 5208 20135 5264
rect 17677 5206 20135 5208
rect 17677 5203 17743 5206
rect 20069 5203 20135 5206
rect 20345 5266 20411 5269
rect 21774 5266 21834 5342
rect 22093 5339 22159 5342
rect 22277 5402 22343 5405
rect 26325 5402 26391 5405
rect 22277 5400 26391 5402
rect 22277 5344 22282 5400
rect 22338 5344 26330 5400
rect 26386 5344 26391 5400
rect 22277 5342 26391 5344
rect 22277 5339 22343 5342
rect 26325 5339 26391 5342
rect 29126 5340 29132 5404
rect 29196 5402 29202 5404
rect 29269 5402 29335 5405
rect 29196 5400 29335 5402
rect 29196 5344 29274 5400
rect 29330 5344 29335 5400
rect 29196 5342 29335 5344
rect 29196 5340 29202 5342
rect 29269 5339 29335 5342
rect 31201 5402 31267 5405
rect 34237 5402 34303 5405
rect 31201 5400 34303 5402
rect 31201 5344 31206 5400
rect 31262 5344 34242 5400
rect 34298 5344 34303 5400
rect 31201 5342 34303 5344
rect 31201 5339 31267 5342
rect 34237 5339 34303 5342
rect 20345 5264 21834 5266
rect 20345 5208 20350 5264
rect 20406 5208 21834 5264
rect 20345 5206 21834 5208
rect 20345 5203 20411 5206
rect 22134 5204 22140 5268
rect 22204 5266 22210 5268
rect 25405 5266 25471 5269
rect 27153 5266 27219 5269
rect 27429 5266 27495 5269
rect 22204 5264 27495 5266
rect 22204 5208 25410 5264
rect 25466 5208 27158 5264
rect 27214 5208 27434 5264
rect 27490 5208 27495 5264
rect 22204 5206 27495 5208
rect 22204 5204 22210 5206
rect 25405 5203 25471 5206
rect 27153 5203 27219 5206
rect 27429 5203 27495 5206
rect 27981 5266 28047 5269
rect 31569 5266 31635 5269
rect 32213 5268 32279 5269
rect 32213 5266 32260 5268
rect 27981 5264 31635 5266
rect 27981 5208 27986 5264
rect 28042 5208 31574 5264
rect 31630 5208 31635 5264
rect 27981 5206 31635 5208
rect 32168 5264 32260 5266
rect 32168 5208 32218 5264
rect 32168 5206 32260 5208
rect 27981 5203 28047 5206
rect 31569 5203 31635 5206
rect 32213 5204 32260 5206
rect 32324 5204 32330 5268
rect 34605 5266 34671 5269
rect 44909 5266 44975 5269
rect 34605 5264 44975 5266
rect 34605 5208 34610 5264
rect 34666 5208 44914 5264
rect 44970 5208 44975 5264
rect 34605 5206 44975 5208
rect 32213 5203 32279 5204
rect 34605 5203 34671 5206
rect 44909 5203 44975 5206
rect 18689 5130 18755 5133
rect 25037 5130 25103 5133
rect 29545 5130 29611 5133
rect 37917 5130 37983 5133
rect 18689 5128 24962 5130
rect 18689 5072 18694 5128
rect 18750 5072 24962 5128
rect 18689 5070 24962 5072
rect 18689 5067 18755 5070
rect 14089 4994 14155 4997
rect 23841 4994 23907 4997
rect 14089 4992 23907 4994
rect 14089 4936 14094 4992
rect 14150 4936 23846 4992
rect 23902 4936 23907 4992
rect 14089 4934 23907 4936
rect 24902 4994 24962 5070
rect 25037 5128 29194 5130
rect 25037 5072 25042 5128
rect 25098 5072 29194 5128
rect 25037 5070 29194 5072
rect 25037 5067 25103 5070
rect 25405 4994 25471 4997
rect 28993 4996 29059 4997
rect 28942 4994 28948 4996
rect 24902 4992 25471 4994
rect 24902 4936 25410 4992
rect 25466 4936 25471 4992
rect 24902 4934 25471 4936
rect 28902 4934 28948 4994
rect 29012 4992 29059 4996
rect 29054 4936 29059 4992
rect 14089 4931 14155 4934
rect 23841 4931 23907 4934
rect 25405 4931 25471 4934
rect 28942 4932 28948 4934
rect 29012 4932 29059 4936
rect 29134 4994 29194 5070
rect 29545 5128 37983 5130
rect 29545 5072 29550 5128
rect 29606 5072 37922 5128
rect 37978 5072 37983 5128
rect 29545 5070 37983 5072
rect 29545 5067 29611 5070
rect 37917 5067 37983 5070
rect 32397 4994 32463 4997
rect 29134 4992 32463 4994
rect 29134 4936 32402 4992
rect 32458 4936 32463 4992
rect 29134 4934 32463 4936
rect 28993 4931 29059 4932
rect 32397 4931 32463 4934
rect 36813 4994 36879 4997
rect 37549 4994 37615 4997
rect 36813 4992 37615 4994
rect 36813 4936 36818 4992
rect 36874 4936 37554 4992
rect 37610 4936 37615 4992
rect 36813 4934 37615 4936
rect 36813 4931 36879 4934
rect 37549 4931 37615 4934
rect 5130 4928 5446 4929
rect 5130 4864 5136 4928
rect 5200 4864 5216 4928
rect 5280 4864 5296 4928
rect 5360 4864 5376 4928
rect 5440 4864 5446 4928
rect 5130 4863 5446 4864
rect 35850 4928 36166 4929
rect 35850 4864 35856 4928
rect 35920 4864 35936 4928
rect 36000 4864 36016 4928
rect 36080 4864 36096 4928
rect 36160 4864 36166 4928
rect 35850 4863 36166 4864
rect 66570 4928 66886 4929
rect 66570 4864 66576 4928
rect 66640 4864 66656 4928
rect 66720 4864 66736 4928
rect 66800 4864 66816 4928
rect 66880 4864 66886 4928
rect 66570 4863 66886 4864
rect 12617 4858 12683 4861
rect 12750 4858 12756 4860
rect 12617 4856 12756 4858
rect 12617 4800 12622 4856
rect 12678 4800 12756 4856
rect 12617 4798 12756 4800
rect 12617 4795 12683 4798
rect 12750 4796 12756 4798
rect 12820 4796 12826 4860
rect 17033 4858 17099 4861
rect 17677 4860 17743 4861
rect 17350 4858 17356 4860
rect 17033 4856 17356 4858
rect 17033 4800 17038 4856
rect 17094 4800 17356 4856
rect 17033 4798 17356 4800
rect 17033 4795 17099 4798
rect 17350 4796 17356 4798
rect 17420 4796 17426 4860
rect 17677 4858 17724 4860
rect 17632 4856 17724 4858
rect 17632 4800 17682 4856
rect 17632 4798 17724 4800
rect 17677 4796 17724 4798
rect 17788 4796 17794 4860
rect 19425 4858 19491 4861
rect 19742 4858 19748 4860
rect 19425 4856 19748 4858
rect 19425 4800 19430 4856
rect 19486 4800 19748 4856
rect 19425 4798 19748 4800
rect 17677 4795 17743 4796
rect 19425 4795 19491 4798
rect 19742 4796 19748 4798
rect 19812 4796 19818 4860
rect 21173 4858 21239 4861
rect 21173 4856 24824 4858
rect 21173 4800 21178 4856
rect 21234 4800 24824 4856
rect 21173 4798 24824 4800
rect 21173 4795 21239 4798
rect 12617 4722 12683 4725
rect 20897 4722 20963 4725
rect 12617 4720 20963 4722
rect 12617 4664 12622 4720
rect 12678 4664 20902 4720
rect 20958 4664 20963 4720
rect 12617 4662 20963 4664
rect 12617 4659 12683 4662
rect 20897 4659 20963 4662
rect 23197 4722 23263 4725
rect 23657 4722 23723 4725
rect 23197 4720 23723 4722
rect 23197 4664 23202 4720
rect 23258 4664 23662 4720
rect 23718 4664 23723 4720
rect 23197 4662 23723 4664
rect 24764 4722 24824 4798
rect 28758 4796 28764 4860
rect 28828 4858 28834 4860
rect 28901 4858 28967 4861
rect 28828 4856 28967 4858
rect 28828 4800 28906 4856
rect 28962 4800 28967 4856
rect 28828 4798 28967 4800
rect 28828 4796 28834 4798
rect 28901 4795 28967 4798
rect 30833 4858 30899 4861
rect 32121 4858 32187 4861
rect 30833 4856 32187 4858
rect 30833 4800 30838 4856
rect 30894 4800 32126 4856
rect 32182 4800 32187 4856
rect 30833 4798 32187 4800
rect 30833 4795 30899 4798
rect 32121 4795 32187 4798
rect 37733 4722 37799 4725
rect 51073 4722 51139 4725
rect 24764 4720 51139 4722
rect 24764 4664 37738 4720
rect 37794 4664 51078 4720
rect 51134 4664 51139 4720
rect 24764 4662 51139 4664
rect 23197 4659 23263 4662
rect 23657 4659 23723 4662
rect 37733 4659 37799 4662
rect 51073 4659 51139 4662
rect 16849 4586 16915 4589
rect 19149 4586 19215 4589
rect 16849 4584 19215 4586
rect 16849 4528 16854 4584
rect 16910 4528 19154 4584
rect 19210 4528 19215 4584
rect 16849 4526 19215 4528
rect 16849 4523 16915 4526
rect 19149 4523 19215 4526
rect 19701 4586 19767 4589
rect 21817 4586 21883 4589
rect 19701 4584 21883 4586
rect 19701 4528 19706 4584
rect 19762 4528 21822 4584
rect 21878 4528 21883 4584
rect 19701 4526 21883 4528
rect 19701 4523 19767 4526
rect 21817 4523 21883 4526
rect 22277 4586 22343 4589
rect 33317 4586 33383 4589
rect 22277 4584 33383 4586
rect 22277 4528 22282 4584
rect 22338 4528 33322 4584
rect 33378 4528 33383 4584
rect 22277 4526 33383 4528
rect 22277 4523 22343 4526
rect 33317 4523 33383 4526
rect 15009 4450 15075 4453
rect 15142 4450 15148 4452
rect 15009 4448 15148 4450
rect 15009 4392 15014 4448
rect 15070 4392 15148 4448
rect 15009 4390 15148 4392
rect 15009 4387 15075 4390
rect 15142 4388 15148 4390
rect 15212 4388 15218 4452
rect 19977 4450 20043 4453
rect 20110 4450 20116 4452
rect 19977 4448 20116 4450
rect 19977 4392 19982 4448
rect 20038 4392 20116 4448
rect 19977 4390 20116 4392
rect 19977 4387 20043 4390
rect 20110 4388 20116 4390
rect 20180 4388 20186 4452
rect 22093 4450 22159 4453
rect 33501 4450 33567 4453
rect 22093 4448 33567 4450
rect 22093 4392 22098 4448
rect 22154 4392 33506 4448
rect 33562 4392 33567 4448
rect 22093 4390 33567 4392
rect 22093 4387 22159 4390
rect 33501 4387 33567 4390
rect 5790 4384 6106 4385
rect 5790 4320 5796 4384
rect 5860 4320 5876 4384
rect 5940 4320 5956 4384
rect 6020 4320 6036 4384
rect 6100 4320 6106 4384
rect 5790 4319 6106 4320
rect 36510 4384 36826 4385
rect 36510 4320 36516 4384
rect 36580 4320 36596 4384
rect 36660 4320 36676 4384
rect 36740 4320 36756 4384
rect 36820 4320 36826 4384
rect 36510 4319 36826 4320
rect 67230 4384 67546 4385
rect 67230 4320 67236 4384
rect 67300 4320 67316 4384
rect 67380 4320 67396 4384
rect 67460 4320 67476 4384
rect 67540 4320 67546 4384
rect 67230 4319 67546 4320
rect 18505 4314 18571 4317
rect 28441 4314 28507 4317
rect 18505 4312 28507 4314
rect 18505 4256 18510 4312
rect 18566 4256 28446 4312
rect 28502 4256 28507 4312
rect 18505 4254 28507 4256
rect 18505 4251 18571 4254
rect 28441 4251 28507 4254
rect 30833 4314 30899 4317
rect 35249 4314 35315 4317
rect 30833 4312 35315 4314
rect 30833 4256 30838 4312
rect 30894 4256 35254 4312
rect 35310 4256 35315 4312
rect 30833 4254 35315 4256
rect 30833 4251 30899 4254
rect 35249 4251 35315 4254
rect 15101 4178 15167 4181
rect 19057 4178 19123 4181
rect 15101 4176 19123 4178
rect 15101 4120 15106 4176
rect 15162 4120 19062 4176
rect 19118 4120 19123 4176
rect 15101 4118 19123 4120
rect 15101 4115 15167 4118
rect 19057 4115 19123 4118
rect 19333 4178 19399 4181
rect 19609 4178 19675 4181
rect 19333 4176 19675 4178
rect 19333 4120 19338 4176
rect 19394 4120 19614 4176
rect 19670 4120 19675 4176
rect 19333 4118 19675 4120
rect 19333 4115 19399 4118
rect 19609 4115 19675 4118
rect 20529 4178 20595 4181
rect 24710 4178 24716 4180
rect 20529 4176 24716 4178
rect 20529 4120 20534 4176
rect 20590 4120 24716 4176
rect 20529 4118 24716 4120
rect 20529 4115 20595 4118
rect 24710 4116 24716 4118
rect 24780 4116 24786 4180
rect 25497 4178 25563 4181
rect 29310 4178 29316 4180
rect 25497 4176 29316 4178
rect 25497 4120 25502 4176
rect 25558 4120 29316 4176
rect 25497 4118 29316 4120
rect 25497 4115 25563 4118
rect 29310 4116 29316 4118
rect 29380 4116 29386 4180
rect 35709 4178 35775 4181
rect 52637 4178 52703 4181
rect 35709 4176 52703 4178
rect 35709 4120 35714 4176
rect 35770 4120 52642 4176
rect 52698 4120 52703 4176
rect 35709 4118 52703 4120
rect 35709 4115 35775 4118
rect 52637 4115 52703 4118
rect 10869 4044 10935 4045
rect 10869 4040 10916 4044
rect 10980 4042 10986 4044
rect 11697 4042 11763 4045
rect 21541 4042 21607 4045
rect 10869 3984 10874 4040
rect 10869 3980 10916 3984
rect 10980 3982 11026 4042
rect 11697 4040 21607 4042
rect 11697 3984 11702 4040
rect 11758 3984 21546 4040
rect 21602 3984 21607 4040
rect 11697 3982 21607 3984
rect 10980 3980 10986 3982
rect 10869 3979 10935 3980
rect 11697 3979 11763 3982
rect 21541 3979 21607 3982
rect 21766 3980 21772 4044
rect 21836 4042 21842 4044
rect 22093 4042 22159 4045
rect 21836 4040 22159 4042
rect 21836 3984 22098 4040
rect 22154 3984 22159 4040
rect 21836 3982 22159 3984
rect 21836 3980 21842 3982
rect 22093 3979 22159 3982
rect 22645 4042 22711 4045
rect 23054 4042 23060 4044
rect 22645 4040 23060 4042
rect 22645 3984 22650 4040
rect 22706 3984 23060 4040
rect 22645 3982 23060 3984
rect 22645 3979 22711 3982
rect 23054 3980 23060 3982
rect 23124 3980 23130 4044
rect 25814 3980 25820 4044
rect 25884 4042 25890 4044
rect 25957 4042 26023 4045
rect 25884 4040 26023 4042
rect 25884 3984 25962 4040
rect 26018 3984 26023 4040
rect 25884 3982 26023 3984
rect 25884 3980 25890 3982
rect 25957 3979 26023 3982
rect 26550 3980 26556 4044
rect 26620 4042 26626 4044
rect 26693 4042 26759 4045
rect 26620 4040 26759 4042
rect 26620 3984 26698 4040
rect 26754 3984 26759 4040
rect 26620 3982 26759 3984
rect 26620 3980 26626 3982
rect 26693 3979 26759 3982
rect 11697 3906 11763 3909
rect 11830 3906 11836 3908
rect 11697 3904 11836 3906
rect 11697 3848 11702 3904
rect 11758 3848 11836 3904
rect 11697 3846 11836 3848
rect 11697 3843 11763 3846
rect 11830 3844 11836 3846
rect 11900 3844 11906 3908
rect 12985 3906 13051 3909
rect 16941 3908 17007 3909
rect 13670 3906 13676 3908
rect 12985 3904 13676 3906
rect 12985 3848 12990 3904
rect 13046 3848 13676 3904
rect 12985 3846 13676 3848
rect 12985 3843 13051 3846
rect 13670 3844 13676 3846
rect 13740 3844 13746 3908
rect 16941 3906 16988 3908
rect 16896 3904 16988 3906
rect 16896 3848 16946 3904
rect 16896 3846 16988 3848
rect 16941 3844 16988 3846
rect 17052 3844 17058 3908
rect 21357 3906 21423 3909
rect 33041 3906 33107 3909
rect 21357 3904 33107 3906
rect 21357 3848 21362 3904
rect 21418 3848 33046 3904
rect 33102 3848 33107 3904
rect 21357 3846 33107 3848
rect 16941 3843 17007 3844
rect 21357 3843 21423 3846
rect 33041 3843 33107 3846
rect 5130 3840 5446 3841
rect 5130 3776 5136 3840
rect 5200 3776 5216 3840
rect 5280 3776 5296 3840
rect 5360 3776 5376 3840
rect 5440 3776 5446 3840
rect 5130 3775 5446 3776
rect 35850 3840 36166 3841
rect 35850 3776 35856 3840
rect 35920 3776 35936 3840
rect 36000 3776 36016 3840
rect 36080 3776 36096 3840
rect 36160 3776 36166 3840
rect 35850 3775 36166 3776
rect 66570 3840 66886 3841
rect 66570 3776 66576 3840
rect 66640 3776 66656 3840
rect 66720 3776 66736 3840
rect 66800 3776 66816 3840
rect 66880 3776 66886 3840
rect 66570 3775 66886 3776
rect 14273 3770 14339 3773
rect 23749 3770 23815 3773
rect 25313 3770 25379 3773
rect 74073 3772 74139 3773
rect 14273 3768 23815 3770
rect 14273 3712 14278 3768
rect 14334 3712 23754 3768
rect 23810 3712 23815 3768
rect 14273 3710 23815 3712
rect 14273 3707 14339 3710
rect 23749 3707 23815 3710
rect 23982 3768 25379 3770
rect 23982 3712 25318 3768
rect 25374 3712 25379 3768
rect 23982 3710 25379 3712
rect 4838 3572 4844 3636
rect 4908 3634 4914 3636
rect 5073 3634 5139 3637
rect 4908 3632 5139 3634
rect 4908 3576 5078 3632
rect 5134 3576 5139 3632
rect 4908 3574 5139 3576
rect 4908 3572 4914 3574
rect 5073 3571 5139 3574
rect 7465 3634 7531 3637
rect 13537 3634 13603 3637
rect 7465 3632 13603 3634
rect 7465 3576 7470 3632
rect 7526 3576 13542 3632
rect 13598 3576 13603 3632
rect 7465 3574 13603 3576
rect 7465 3571 7531 3574
rect 13537 3571 13603 3574
rect 13997 3634 14063 3637
rect 23982 3634 24042 3710
rect 25313 3707 25379 3710
rect 74022 3708 74028 3772
rect 74092 3770 74139 3772
rect 74092 3768 74184 3770
rect 74134 3712 74184 3768
rect 74092 3710 74184 3712
rect 74092 3708 74139 3710
rect 74073 3707 74139 3708
rect 13997 3632 24042 3634
rect 13997 3576 14002 3632
rect 14058 3576 24042 3632
rect 13997 3574 24042 3576
rect 24853 3634 24919 3637
rect 27061 3634 27127 3637
rect 24853 3632 27127 3634
rect 24853 3576 24858 3632
rect 24914 3576 27066 3632
rect 27122 3576 27127 3632
rect 24853 3574 27127 3576
rect 13997 3571 14063 3574
rect 24853 3571 24919 3574
rect 27061 3571 27127 3574
rect 28073 3634 28139 3637
rect 28574 3634 28580 3636
rect 28073 3632 28580 3634
rect 28073 3576 28078 3632
rect 28134 3576 28580 3632
rect 28073 3574 28580 3576
rect 28073 3571 28139 3574
rect 28574 3572 28580 3574
rect 28644 3572 28650 3636
rect 34053 3634 34119 3637
rect 34329 3634 34395 3637
rect 37917 3634 37983 3637
rect 34053 3632 37983 3634
rect 34053 3576 34058 3632
rect 34114 3576 34334 3632
rect 34390 3576 37922 3632
rect 37978 3576 37983 3632
rect 34053 3574 37983 3576
rect 34053 3571 34119 3574
rect 34329 3571 34395 3574
rect 37917 3571 37983 3574
rect 10225 3498 10291 3501
rect 20897 3498 20963 3501
rect 10225 3496 20963 3498
rect 10225 3440 10230 3496
rect 10286 3440 20902 3496
rect 20958 3440 20963 3496
rect 10225 3438 20963 3440
rect 10225 3435 10291 3438
rect 20897 3435 20963 3438
rect 25037 3498 25103 3501
rect 32857 3498 32923 3501
rect 25037 3496 32923 3498
rect 25037 3440 25042 3496
rect 25098 3440 32862 3496
rect 32918 3440 32923 3496
rect 25037 3438 32923 3440
rect 25037 3435 25103 3438
rect 32857 3435 32923 3438
rect 33777 3498 33843 3501
rect 38653 3498 38719 3501
rect 33777 3496 38719 3498
rect 33777 3440 33782 3496
rect 33838 3440 38658 3496
rect 38714 3440 38719 3496
rect 33777 3438 38719 3440
rect 33777 3435 33843 3438
rect 38653 3435 38719 3438
rect 11329 3362 11395 3365
rect 12709 3362 12775 3365
rect 13629 3362 13695 3365
rect 15653 3362 15719 3365
rect 11329 3360 15719 3362
rect 11329 3304 11334 3360
rect 11390 3304 12714 3360
rect 12770 3304 13634 3360
rect 13690 3304 15658 3360
rect 15714 3304 15719 3360
rect 11329 3302 15719 3304
rect 11329 3299 11395 3302
rect 12709 3299 12775 3302
rect 13629 3299 13695 3302
rect 15653 3299 15719 3302
rect 15929 3362 15995 3365
rect 16062 3362 16068 3364
rect 15929 3360 16068 3362
rect 15929 3304 15934 3360
rect 15990 3304 16068 3360
rect 15929 3302 16068 3304
rect 15929 3299 15995 3302
rect 16062 3300 16068 3302
rect 16132 3300 16138 3364
rect 22001 3362 22067 3365
rect 25405 3362 25471 3365
rect 22001 3360 25471 3362
rect 22001 3304 22006 3360
rect 22062 3304 25410 3360
rect 25466 3304 25471 3360
rect 22001 3302 25471 3304
rect 22001 3299 22067 3302
rect 25405 3299 25471 3302
rect 26693 3362 26759 3365
rect 31886 3362 31892 3364
rect 26693 3360 31892 3362
rect 26693 3304 26698 3360
rect 26754 3304 31892 3360
rect 26693 3302 31892 3304
rect 26693 3299 26759 3302
rect 31886 3300 31892 3302
rect 31956 3300 31962 3364
rect 33777 3362 33843 3365
rect 35157 3362 35223 3365
rect 33777 3360 35223 3362
rect 33777 3304 33782 3360
rect 33838 3304 35162 3360
rect 35218 3304 35223 3360
rect 33777 3302 35223 3304
rect 33777 3299 33843 3302
rect 35157 3299 35223 3302
rect 5790 3296 6106 3297
rect 5790 3232 5796 3296
rect 5860 3232 5876 3296
rect 5940 3232 5956 3296
rect 6020 3232 6036 3296
rect 6100 3232 6106 3296
rect 5790 3231 6106 3232
rect 7649 3226 7715 3229
rect 15469 3226 15535 3229
rect 7649 3224 15535 3226
rect 7649 3168 7654 3224
rect 7710 3168 15474 3224
rect 15530 3168 15535 3224
rect 7649 3166 15535 3168
rect 15656 3226 15716 3299
rect 36510 3296 36826 3297
rect 36510 3232 36516 3296
rect 36580 3232 36596 3296
rect 36660 3232 36676 3296
rect 36740 3232 36756 3296
rect 36820 3232 36826 3296
rect 36510 3231 36826 3232
rect 67230 3296 67546 3297
rect 67230 3232 67236 3296
rect 67300 3232 67316 3296
rect 67380 3232 67396 3296
rect 67460 3232 67476 3296
rect 67540 3232 67546 3296
rect 67230 3231 67546 3232
rect 16849 3226 16915 3229
rect 15656 3224 16915 3226
rect 15656 3168 16854 3224
rect 16910 3168 16915 3224
rect 15656 3166 16915 3168
rect 7649 3163 7715 3166
rect 15469 3163 15535 3166
rect 16849 3163 16915 3166
rect 22277 3226 22343 3229
rect 23422 3226 23428 3228
rect 22277 3224 23428 3226
rect 22277 3168 22282 3224
rect 22338 3168 23428 3224
rect 22277 3166 23428 3168
rect 22277 3163 22343 3166
rect 23422 3164 23428 3166
rect 23492 3164 23498 3228
rect 25262 3164 25268 3228
rect 25332 3226 25338 3228
rect 28717 3226 28783 3229
rect 31753 3226 31819 3229
rect 33869 3226 33935 3229
rect 25332 3166 28642 3226
rect 25332 3164 25338 3166
rect 8385 3090 8451 3093
rect 19517 3090 19583 3093
rect 8385 3088 19583 3090
rect 8385 3032 8390 3088
rect 8446 3032 19522 3088
rect 19578 3032 19583 3088
rect 8385 3030 19583 3032
rect 8385 3027 8451 3030
rect 19517 3027 19583 3030
rect 19885 3090 19951 3093
rect 21725 3090 21791 3093
rect 24577 3090 24643 3093
rect 19885 3088 24643 3090
rect 19885 3032 19890 3088
rect 19946 3032 21730 3088
rect 21786 3032 24582 3088
rect 24638 3032 24643 3088
rect 19885 3030 24643 3032
rect 19885 3027 19951 3030
rect 21725 3027 21791 3030
rect 24577 3027 24643 3030
rect 25129 3090 25195 3093
rect 25405 3090 25471 3093
rect 27337 3092 27403 3093
rect 27286 3090 27292 3092
rect 25129 3088 25471 3090
rect 25129 3032 25134 3088
rect 25190 3032 25410 3088
rect 25466 3032 25471 3088
rect 25129 3030 25471 3032
rect 27246 3030 27292 3090
rect 27356 3088 27403 3092
rect 27398 3032 27403 3088
rect 25129 3027 25195 3030
rect 25405 3027 25471 3030
rect 27286 3028 27292 3030
rect 27356 3028 27403 3032
rect 28582 3090 28642 3166
rect 28717 3224 33935 3226
rect 28717 3168 28722 3224
rect 28778 3168 31758 3224
rect 31814 3168 33874 3224
rect 33930 3168 33935 3224
rect 28717 3166 33935 3168
rect 28717 3163 28783 3166
rect 31753 3163 31819 3166
rect 33869 3163 33935 3166
rect 42977 3090 43043 3093
rect 28582 3088 43043 3090
rect 28582 3032 42982 3088
rect 43038 3032 43043 3088
rect 28582 3030 43043 3032
rect 27337 3027 27403 3028
rect 42977 3027 43043 3030
rect 10501 2954 10567 2957
rect 13905 2954 13971 2957
rect 10501 2952 13971 2954
rect 10501 2896 10506 2952
rect 10562 2896 13910 2952
rect 13966 2896 13971 2952
rect 10501 2894 13971 2896
rect 10501 2891 10567 2894
rect 13905 2891 13971 2894
rect 23289 2954 23355 2957
rect 33041 2954 33107 2957
rect 23289 2952 33107 2954
rect 23289 2896 23294 2952
rect 23350 2896 33046 2952
rect 33102 2896 33107 2952
rect 23289 2894 33107 2896
rect 23289 2891 23355 2894
rect 33041 2891 33107 2894
rect 36905 2954 36971 2957
rect 37038 2954 37044 2956
rect 36905 2952 37044 2954
rect 36905 2896 36910 2952
rect 36966 2896 37044 2952
rect 36905 2894 37044 2896
rect 36905 2891 36971 2894
rect 37038 2892 37044 2894
rect 37108 2892 37114 2956
rect 9949 2818 10015 2821
rect 17953 2818 18019 2821
rect 9949 2816 18019 2818
rect 9949 2760 9954 2816
rect 10010 2760 17958 2816
rect 18014 2760 18019 2816
rect 9949 2758 18019 2760
rect 9949 2755 10015 2758
rect 17953 2755 18019 2758
rect 25221 2818 25287 2821
rect 31150 2818 31156 2820
rect 25221 2816 31156 2818
rect 25221 2760 25226 2816
rect 25282 2760 31156 2816
rect 25221 2758 31156 2760
rect 25221 2755 25287 2758
rect 31150 2756 31156 2758
rect 31220 2756 31226 2820
rect 36261 2818 36327 2821
rect 37549 2818 37615 2821
rect 36261 2816 37615 2818
rect 36261 2760 36266 2816
rect 36322 2760 37554 2816
rect 37610 2760 37615 2816
rect 36261 2758 37615 2760
rect 36261 2755 36327 2758
rect 37549 2755 37615 2758
rect 5130 2752 5446 2753
rect 5130 2688 5136 2752
rect 5200 2688 5216 2752
rect 5280 2688 5296 2752
rect 5360 2688 5376 2752
rect 5440 2688 5446 2752
rect 5130 2687 5446 2688
rect 35850 2752 36166 2753
rect 35850 2688 35856 2752
rect 35920 2688 35936 2752
rect 36000 2688 36016 2752
rect 36080 2688 36096 2752
rect 36160 2688 36166 2752
rect 35850 2687 36166 2688
rect 66570 2752 66886 2753
rect 66570 2688 66576 2752
rect 66640 2688 66656 2752
rect 66720 2688 66736 2752
rect 66800 2688 66816 2752
rect 66880 2688 66886 2752
rect 66570 2687 66886 2688
rect 10409 2682 10475 2685
rect 10726 2682 10732 2684
rect 10409 2680 10732 2682
rect 10409 2624 10414 2680
rect 10470 2624 10732 2680
rect 10409 2622 10732 2624
rect 10409 2619 10475 2622
rect 10726 2620 10732 2622
rect 10796 2620 10802 2684
rect 18270 2682 18276 2684
rect 12390 2622 18276 2682
rect 5809 2546 5875 2549
rect 12390 2546 12450 2622
rect 18270 2620 18276 2622
rect 18340 2620 18346 2684
rect 24393 2682 24459 2685
rect 33542 2682 33548 2684
rect 24393 2680 33548 2682
rect 24393 2624 24398 2680
rect 24454 2624 33548 2680
rect 24393 2622 33548 2624
rect 24393 2619 24459 2622
rect 33542 2620 33548 2622
rect 33612 2620 33618 2684
rect 5809 2544 12450 2546
rect 5809 2488 5814 2544
rect 5870 2488 12450 2544
rect 5809 2486 12450 2488
rect 5809 2483 5875 2486
rect 17902 2484 17908 2548
rect 17972 2546 17978 2548
rect 19333 2546 19399 2549
rect 17972 2544 19399 2546
rect 17972 2488 19338 2544
rect 19394 2488 19399 2544
rect 17972 2486 19399 2488
rect 17972 2484 17978 2486
rect 19333 2483 19399 2486
rect 25313 2546 25379 2549
rect 33358 2546 33364 2548
rect 25313 2544 33364 2546
rect 25313 2488 25318 2544
rect 25374 2488 33364 2544
rect 25313 2486 33364 2488
rect 25313 2483 25379 2486
rect 33358 2484 33364 2486
rect 33428 2484 33434 2548
rect 5625 2410 5691 2413
rect 18454 2410 18460 2412
rect 5625 2408 18460 2410
rect 5625 2352 5630 2408
rect 5686 2352 18460 2408
rect 5625 2350 18460 2352
rect 5625 2347 5691 2350
rect 18454 2348 18460 2350
rect 18524 2348 18530 2412
rect 24577 2410 24643 2413
rect 24710 2410 24716 2412
rect 24577 2408 24716 2410
rect 24577 2352 24582 2408
rect 24638 2352 24716 2408
rect 24577 2350 24716 2352
rect 24577 2347 24643 2350
rect 24710 2348 24716 2350
rect 24780 2348 24786 2412
rect 28809 2410 28875 2413
rect 41781 2410 41847 2413
rect 28809 2408 41847 2410
rect 28809 2352 28814 2408
rect 28870 2352 41786 2408
rect 41842 2352 41847 2408
rect 28809 2350 41847 2352
rect 28809 2347 28875 2350
rect 41781 2347 41847 2350
rect 20713 2274 20779 2277
rect 26233 2274 26299 2277
rect 34462 2274 34468 2276
rect 20713 2272 22110 2274
rect 20713 2216 20718 2272
rect 20774 2216 22110 2272
rect 20713 2214 22110 2216
rect 20713 2211 20779 2214
rect 5790 2208 6106 2209
rect 5790 2144 5796 2208
rect 5860 2144 5876 2208
rect 5940 2144 5956 2208
rect 6020 2144 6036 2208
rect 6100 2144 6106 2208
rect 5790 2143 6106 2144
rect 22050 2138 22110 2214
rect 26233 2272 34468 2274
rect 26233 2216 26238 2272
rect 26294 2216 34468 2272
rect 26233 2214 34468 2216
rect 26233 2211 26299 2214
rect 34462 2212 34468 2214
rect 34532 2212 34538 2276
rect 36510 2208 36826 2209
rect 36510 2144 36516 2208
rect 36580 2144 36596 2208
rect 36660 2144 36676 2208
rect 36740 2144 36756 2208
rect 36820 2144 36826 2208
rect 36510 2143 36826 2144
rect 67230 2208 67546 2209
rect 67230 2144 67236 2208
rect 67300 2144 67316 2208
rect 67380 2144 67396 2208
rect 67460 2144 67476 2208
rect 67540 2144 67546 2208
rect 67230 2143 67546 2144
rect 33174 2138 33180 2140
rect 22050 2078 33180 2138
rect 33174 2076 33180 2078
rect 33244 2076 33250 2140
rect 28073 1866 28139 1869
rect 38285 1866 38351 1869
rect 28073 1864 38351 1866
rect 28073 1808 28078 1864
rect 28134 1808 38290 1864
rect 38346 1808 38351 1864
rect 28073 1806 38351 1808
rect 28073 1803 28139 1806
rect 38285 1803 38351 1806
rect 21541 1730 21607 1733
rect 30230 1730 30236 1732
rect 21541 1728 30236 1730
rect 21541 1672 21546 1728
rect 21602 1672 30236 1728
rect 21541 1670 30236 1672
rect 21541 1667 21607 1670
rect 30230 1668 30236 1670
rect 30300 1668 30306 1732
rect 19977 1458 20043 1461
rect 20805 1458 20871 1461
rect 19977 1456 20871 1458
rect 19977 1400 19982 1456
rect 20038 1400 20810 1456
rect 20866 1400 20871 1456
rect 19977 1398 20871 1400
rect 19977 1395 20043 1398
rect 20805 1395 20871 1398
rect 22553 1458 22619 1461
rect 23657 1458 23723 1461
rect 22553 1456 23723 1458
rect 22553 1400 22558 1456
rect 22614 1400 23662 1456
rect 23718 1400 23723 1456
rect 22553 1398 23723 1400
rect 22553 1395 22619 1398
rect 23657 1395 23723 1398
rect 36077 1458 36143 1461
rect 37273 1458 37339 1461
rect 36077 1456 37339 1458
rect 36077 1400 36082 1456
rect 36138 1400 37278 1456
rect 37334 1400 37339 1456
rect 36077 1398 37339 1400
rect 36077 1395 36143 1398
rect 37273 1395 37339 1398
rect 17401 1322 17467 1325
rect 19333 1322 19399 1325
rect 17401 1320 19399 1322
rect 17401 1264 17406 1320
rect 17462 1264 19338 1320
rect 19394 1264 19399 1320
rect 17401 1262 19399 1264
rect 17401 1259 17467 1262
rect 19333 1259 19399 1262
rect 18597 1186 18663 1189
rect 23841 1186 23907 1189
rect 18597 1184 23907 1186
rect 18597 1128 18602 1184
rect 18658 1128 23846 1184
rect 23902 1128 23907 1184
rect 18597 1126 23907 1128
rect 18597 1123 18663 1126
rect 23841 1123 23907 1126
rect 19190 988 19196 1052
rect 19260 1050 19266 1052
rect 25773 1050 25839 1053
rect 19260 1048 25839 1050
rect 19260 992 25778 1048
rect 25834 992 25839 1048
rect 19260 990 25839 992
rect 19260 988 19266 990
rect 25773 987 25839 990
<< via3 >>
rect 5136 37564 5200 37568
rect 5136 37508 5140 37564
rect 5140 37508 5196 37564
rect 5196 37508 5200 37564
rect 5136 37504 5200 37508
rect 5216 37564 5280 37568
rect 5216 37508 5220 37564
rect 5220 37508 5276 37564
rect 5276 37508 5280 37564
rect 5216 37504 5280 37508
rect 5296 37564 5360 37568
rect 5296 37508 5300 37564
rect 5300 37508 5356 37564
rect 5356 37508 5360 37564
rect 5296 37504 5360 37508
rect 5376 37564 5440 37568
rect 5376 37508 5380 37564
rect 5380 37508 5436 37564
rect 5436 37508 5440 37564
rect 5376 37504 5440 37508
rect 35856 37564 35920 37568
rect 35856 37508 35860 37564
rect 35860 37508 35916 37564
rect 35916 37508 35920 37564
rect 35856 37504 35920 37508
rect 35936 37564 36000 37568
rect 35936 37508 35940 37564
rect 35940 37508 35996 37564
rect 35996 37508 36000 37564
rect 35936 37504 36000 37508
rect 36016 37564 36080 37568
rect 36016 37508 36020 37564
rect 36020 37508 36076 37564
rect 36076 37508 36080 37564
rect 36016 37504 36080 37508
rect 36096 37564 36160 37568
rect 36096 37508 36100 37564
rect 36100 37508 36156 37564
rect 36156 37508 36160 37564
rect 36096 37504 36160 37508
rect 66576 37564 66640 37568
rect 66576 37508 66580 37564
rect 66580 37508 66636 37564
rect 66636 37508 66640 37564
rect 66576 37504 66640 37508
rect 66656 37564 66720 37568
rect 66656 37508 66660 37564
rect 66660 37508 66716 37564
rect 66716 37508 66720 37564
rect 66656 37504 66720 37508
rect 66736 37564 66800 37568
rect 66736 37508 66740 37564
rect 66740 37508 66796 37564
rect 66796 37508 66800 37564
rect 66736 37504 66800 37508
rect 66816 37564 66880 37568
rect 66816 37508 66820 37564
rect 66820 37508 66876 37564
rect 66876 37508 66880 37564
rect 66816 37504 66880 37508
rect 5796 37020 5860 37024
rect 5796 36964 5800 37020
rect 5800 36964 5856 37020
rect 5856 36964 5860 37020
rect 5796 36960 5860 36964
rect 5876 37020 5940 37024
rect 5876 36964 5880 37020
rect 5880 36964 5936 37020
rect 5936 36964 5940 37020
rect 5876 36960 5940 36964
rect 5956 37020 6020 37024
rect 5956 36964 5960 37020
rect 5960 36964 6016 37020
rect 6016 36964 6020 37020
rect 5956 36960 6020 36964
rect 6036 37020 6100 37024
rect 6036 36964 6040 37020
rect 6040 36964 6096 37020
rect 6096 36964 6100 37020
rect 6036 36960 6100 36964
rect 36516 37020 36580 37024
rect 36516 36964 36520 37020
rect 36520 36964 36576 37020
rect 36576 36964 36580 37020
rect 36516 36960 36580 36964
rect 36596 37020 36660 37024
rect 36596 36964 36600 37020
rect 36600 36964 36656 37020
rect 36656 36964 36660 37020
rect 36596 36960 36660 36964
rect 36676 37020 36740 37024
rect 36676 36964 36680 37020
rect 36680 36964 36736 37020
rect 36736 36964 36740 37020
rect 36676 36960 36740 36964
rect 36756 37020 36820 37024
rect 36756 36964 36760 37020
rect 36760 36964 36816 37020
rect 36816 36964 36820 37020
rect 36756 36960 36820 36964
rect 67236 37020 67300 37024
rect 67236 36964 67240 37020
rect 67240 36964 67296 37020
rect 67296 36964 67300 37020
rect 67236 36960 67300 36964
rect 67316 37020 67380 37024
rect 67316 36964 67320 37020
rect 67320 36964 67376 37020
rect 67376 36964 67380 37020
rect 67316 36960 67380 36964
rect 67396 37020 67460 37024
rect 67396 36964 67400 37020
rect 67400 36964 67456 37020
rect 67456 36964 67460 37020
rect 67396 36960 67460 36964
rect 67476 37020 67540 37024
rect 67476 36964 67480 37020
rect 67480 36964 67536 37020
rect 67536 36964 67540 37020
rect 67476 36960 67540 36964
rect 7052 36544 7116 36548
rect 7052 36488 7066 36544
rect 7066 36488 7116 36544
rect 7052 36484 7116 36488
rect 32812 36544 32876 36548
rect 32812 36488 32826 36544
rect 32826 36488 32876 36544
rect 32812 36484 32876 36488
rect 5136 36476 5200 36480
rect 5136 36420 5140 36476
rect 5140 36420 5196 36476
rect 5196 36420 5200 36476
rect 5136 36416 5200 36420
rect 5216 36476 5280 36480
rect 5216 36420 5220 36476
rect 5220 36420 5276 36476
rect 5276 36420 5280 36476
rect 5216 36416 5280 36420
rect 5296 36476 5360 36480
rect 5296 36420 5300 36476
rect 5300 36420 5356 36476
rect 5356 36420 5360 36476
rect 5296 36416 5360 36420
rect 5376 36476 5440 36480
rect 5376 36420 5380 36476
rect 5380 36420 5436 36476
rect 5436 36420 5440 36476
rect 5376 36416 5440 36420
rect 35856 36476 35920 36480
rect 35856 36420 35860 36476
rect 35860 36420 35916 36476
rect 35916 36420 35920 36476
rect 35856 36416 35920 36420
rect 35936 36476 36000 36480
rect 35936 36420 35940 36476
rect 35940 36420 35996 36476
rect 35996 36420 36000 36476
rect 35936 36416 36000 36420
rect 36016 36476 36080 36480
rect 36016 36420 36020 36476
rect 36020 36420 36076 36476
rect 36076 36420 36080 36476
rect 36016 36416 36080 36420
rect 36096 36476 36160 36480
rect 36096 36420 36100 36476
rect 36100 36420 36156 36476
rect 36156 36420 36160 36476
rect 36096 36416 36160 36420
rect 66576 36476 66640 36480
rect 66576 36420 66580 36476
rect 66580 36420 66636 36476
rect 66636 36420 66640 36476
rect 66576 36416 66640 36420
rect 66656 36476 66720 36480
rect 66656 36420 66660 36476
rect 66660 36420 66716 36476
rect 66716 36420 66720 36476
rect 66656 36416 66720 36420
rect 66736 36476 66800 36480
rect 66736 36420 66740 36476
rect 66740 36420 66796 36476
rect 66796 36420 66800 36476
rect 66736 36416 66800 36420
rect 66816 36476 66880 36480
rect 66816 36420 66820 36476
rect 66820 36420 66876 36476
rect 66876 36420 66880 36476
rect 66816 36416 66880 36420
rect 5796 35932 5860 35936
rect 5796 35876 5800 35932
rect 5800 35876 5856 35932
rect 5856 35876 5860 35932
rect 5796 35872 5860 35876
rect 5876 35932 5940 35936
rect 5876 35876 5880 35932
rect 5880 35876 5936 35932
rect 5936 35876 5940 35932
rect 5876 35872 5940 35876
rect 5956 35932 6020 35936
rect 5956 35876 5960 35932
rect 5960 35876 6016 35932
rect 6016 35876 6020 35932
rect 5956 35872 6020 35876
rect 6036 35932 6100 35936
rect 6036 35876 6040 35932
rect 6040 35876 6096 35932
rect 6096 35876 6100 35932
rect 6036 35872 6100 35876
rect 36516 35932 36580 35936
rect 36516 35876 36520 35932
rect 36520 35876 36576 35932
rect 36576 35876 36580 35932
rect 36516 35872 36580 35876
rect 36596 35932 36660 35936
rect 36596 35876 36600 35932
rect 36600 35876 36656 35932
rect 36656 35876 36660 35932
rect 36596 35872 36660 35876
rect 36676 35932 36740 35936
rect 36676 35876 36680 35932
rect 36680 35876 36736 35932
rect 36736 35876 36740 35932
rect 36676 35872 36740 35876
rect 36756 35932 36820 35936
rect 36756 35876 36760 35932
rect 36760 35876 36816 35932
rect 36816 35876 36820 35932
rect 36756 35872 36820 35876
rect 67236 35932 67300 35936
rect 67236 35876 67240 35932
rect 67240 35876 67296 35932
rect 67296 35876 67300 35932
rect 67236 35872 67300 35876
rect 67316 35932 67380 35936
rect 67316 35876 67320 35932
rect 67320 35876 67376 35932
rect 67376 35876 67380 35932
rect 67316 35872 67380 35876
rect 67396 35932 67460 35936
rect 67396 35876 67400 35932
rect 67400 35876 67456 35932
rect 67456 35876 67460 35932
rect 67396 35872 67460 35876
rect 67476 35932 67540 35936
rect 67476 35876 67480 35932
rect 67480 35876 67536 35932
rect 67536 35876 67540 35932
rect 67476 35872 67540 35876
rect 5136 35388 5200 35392
rect 5136 35332 5140 35388
rect 5140 35332 5196 35388
rect 5196 35332 5200 35388
rect 5136 35328 5200 35332
rect 5216 35388 5280 35392
rect 5216 35332 5220 35388
rect 5220 35332 5276 35388
rect 5276 35332 5280 35388
rect 5216 35328 5280 35332
rect 5296 35388 5360 35392
rect 5296 35332 5300 35388
rect 5300 35332 5356 35388
rect 5356 35332 5360 35388
rect 5296 35328 5360 35332
rect 5376 35388 5440 35392
rect 5376 35332 5380 35388
rect 5380 35332 5436 35388
rect 5436 35332 5440 35388
rect 5376 35328 5440 35332
rect 35856 35388 35920 35392
rect 35856 35332 35860 35388
rect 35860 35332 35916 35388
rect 35916 35332 35920 35388
rect 35856 35328 35920 35332
rect 35936 35388 36000 35392
rect 35936 35332 35940 35388
rect 35940 35332 35996 35388
rect 35996 35332 36000 35388
rect 35936 35328 36000 35332
rect 36016 35388 36080 35392
rect 36016 35332 36020 35388
rect 36020 35332 36076 35388
rect 36076 35332 36080 35388
rect 36016 35328 36080 35332
rect 36096 35388 36160 35392
rect 36096 35332 36100 35388
rect 36100 35332 36156 35388
rect 36156 35332 36160 35388
rect 36096 35328 36160 35332
rect 66576 35388 66640 35392
rect 66576 35332 66580 35388
rect 66580 35332 66636 35388
rect 66636 35332 66640 35388
rect 66576 35328 66640 35332
rect 66656 35388 66720 35392
rect 66656 35332 66660 35388
rect 66660 35332 66716 35388
rect 66716 35332 66720 35388
rect 66656 35328 66720 35332
rect 66736 35388 66800 35392
rect 66736 35332 66740 35388
rect 66740 35332 66796 35388
rect 66796 35332 66800 35388
rect 66736 35328 66800 35332
rect 66816 35388 66880 35392
rect 66816 35332 66820 35388
rect 66820 35332 66876 35388
rect 66876 35332 66880 35388
rect 66816 35328 66880 35332
rect 5796 34844 5860 34848
rect 5796 34788 5800 34844
rect 5800 34788 5856 34844
rect 5856 34788 5860 34844
rect 5796 34784 5860 34788
rect 5876 34844 5940 34848
rect 5876 34788 5880 34844
rect 5880 34788 5936 34844
rect 5936 34788 5940 34844
rect 5876 34784 5940 34788
rect 5956 34844 6020 34848
rect 5956 34788 5960 34844
rect 5960 34788 6016 34844
rect 6016 34788 6020 34844
rect 5956 34784 6020 34788
rect 6036 34844 6100 34848
rect 6036 34788 6040 34844
rect 6040 34788 6096 34844
rect 6096 34788 6100 34844
rect 6036 34784 6100 34788
rect 36516 34844 36580 34848
rect 36516 34788 36520 34844
rect 36520 34788 36576 34844
rect 36576 34788 36580 34844
rect 36516 34784 36580 34788
rect 36596 34844 36660 34848
rect 36596 34788 36600 34844
rect 36600 34788 36656 34844
rect 36656 34788 36660 34844
rect 36596 34784 36660 34788
rect 36676 34844 36740 34848
rect 36676 34788 36680 34844
rect 36680 34788 36736 34844
rect 36736 34788 36740 34844
rect 36676 34784 36740 34788
rect 36756 34844 36820 34848
rect 36756 34788 36760 34844
rect 36760 34788 36816 34844
rect 36816 34788 36820 34844
rect 36756 34784 36820 34788
rect 67236 34844 67300 34848
rect 67236 34788 67240 34844
rect 67240 34788 67296 34844
rect 67296 34788 67300 34844
rect 67236 34784 67300 34788
rect 67316 34844 67380 34848
rect 67316 34788 67320 34844
rect 67320 34788 67376 34844
rect 67376 34788 67380 34844
rect 67316 34784 67380 34788
rect 67396 34844 67460 34848
rect 67396 34788 67400 34844
rect 67400 34788 67456 34844
rect 67456 34788 67460 34844
rect 67396 34784 67460 34788
rect 67476 34844 67540 34848
rect 67476 34788 67480 34844
rect 67480 34788 67536 34844
rect 67536 34788 67540 34844
rect 67476 34784 67540 34788
rect 5136 34300 5200 34304
rect 5136 34244 5140 34300
rect 5140 34244 5196 34300
rect 5196 34244 5200 34300
rect 5136 34240 5200 34244
rect 5216 34300 5280 34304
rect 5216 34244 5220 34300
rect 5220 34244 5276 34300
rect 5276 34244 5280 34300
rect 5216 34240 5280 34244
rect 5296 34300 5360 34304
rect 5296 34244 5300 34300
rect 5300 34244 5356 34300
rect 5356 34244 5360 34300
rect 5296 34240 5360 34244
rect 5376 34300 5440 34304
rect 5376 34244 5380 34300
rect 5380 34244 5436 34300
rect 5436 34244 5440 34300
rect 5376 34240 5440 34244
rect 35856 34300 35920 34304
rect 35856 34244 35860 34300
rect 35860 34244 35916 34300
rect 35916 34244 35920 34300
rect 35856 34240 35920 34244
rect 35936 34300 36000 34304
rect 35936 34244 35940 34300
rect 35940 34244 35996 34300
rect 35996 34244 36000 34300
rect 35936 34240 36000 34244
rect 36016 34300 36080 34304
rect 36016 34244 36020 34300
rect 36020 34244 36076 34300
rect 36076 34244 36080 34300
rect 36016 34240 36080 34244
rect 36096 34300 36160 34304
rect 36096 34244 36100 34300
rect 36100 34244 36156 34300
rect 36156 34244 36160 34300
rect 36096 34240 36160 34244
rect 66576 34300 66640 34304
rect 66576 34244 66580 34300
rect 66580 34244 66636 34300
rect 66636 34244 66640 34300
rect 66576 34240 66640 34244
rect 66656 34300 66720 34304
rect 66656 34244 66660 34300
rect 66660 34244 66716 34300
rect 66716 34244 66720 34300
rect 66656 34240 66720 34244
rect 66736 34300 66800 34304
rect 66736 34244 66740 34300
rect 66740 34244 66796 34300
rect 66796 34244 66800 34300
rect 66736 34240 66800 34244
rect 66816 34300 66880 34304
rect 66816 34244 66820 34300
rect 66820 34244 66876 34300
rect 66876 34244 66880 34300
rect 66816 34240 66880 34244
rect 5796 33756 5860 33760
rect 5796 33700 5800 33756
rect 5800 33700 5856 33756
rect 5856 33700 5860 33756
rect 5796 33696 5860 33700
rect 5876 33756 5940 33760
rect 5876 33700 5880 33756
rect 5880 33700 5936 33756
rect 5936 33700 5940 33756
rect 5876 33696 5940 33700
rect 5956 33756 6020 33760
rect 5956 33700 5960 33756
rect 5960 33700 6016 33756
rect 6016 33700 6020 33756
rect 5956 33696 6020 33700
rect 6036 33756 6100 33760
rect 6036 33700 6040 33756
rect 6040 33700 6096 33756
rect 6096 33700 6100 33756
rect 6036 33696 6100 33700
rect 36516 33756 36580 33760
rect 36516 33700 36520 33756
rect 36520 33700 36576 33756
rect 36576 33700 36580 33756
rect 36516 33696 36580 33700
rect 36596 33756 36660 33760
rect 36596 33700 36600 33756
rect 36600 33700 36656 33756
rect 36656 33700 36660 33756
rect 36596 33696 36660 33700
rect 36676 33756 36740 33760
rect 36676 33700 36680 33756
rect 36680 33700 36736 33756
rect 36736 33700 36740 33756
rect 36676 33696 36740 33700
rect 36756 33756 36820 33760
rect 36756 33700 36760 33756
rect 36760 33700 36816 33756
rect 36816 33700 36820 33756
rect 36756 33696 36820 33700
rect 67236 33756 67300 33760
rect 67236 33700 67240 33756
rect 67240 33700 67296 33756
rect 67296 33700 67300 33756
rect 67236 33696 67300 33700
rect 67316 33756 67380 33760
rect 67316 33700 67320 33756
rect 67320 33700 67376 33756
rect 67376 33700 67380 33756
rect 67316 33696 67380 33700
rect 67396 33756 67460 33760
rect 67396 33700 67400 33756
rect 67400 33700 67456 33756
rect 67456 33700 67460 33756
rect 67396 33696 67460 33700
rect 67476 33756 67540 33760
rect 67476 33700 67480 33756
rect 67480 33700 67536 33756
rect 67536 33700 67540 33756
rect 67476 33696 67540 33700
rect 5136 33212 5200 33216
rect 5136 33156 5140 33212
rect 5140 33156 5196 33212
rect 5196 33156 5200 33212
rect 5136 33152 5200 33156
rect 5216 33212 5280 33216
rect 5216 33156 5220 33212
rect 5220 33156 5276 33212
rect 5276 33156 5280 33212
rect 5216 33152 5280 33156
rect 5296 33212 5360 33216
rect 5296 33156 5300 33212
rect 5300 33156 5356 33212
rect 5356 33156 5360 33212
rect 5296 33152 5360 33156
rect 5376 33212 5440 33216
rect 5376 33156 5380 33212
rect 5380 33156 5436 33212
rect 5436 33156 5440 33212
rect 5376 33152 5440 33156
rect 35856 33212 35920 33216
rect 35856 33156 35860 33212
rect 35860 33156 35916 33212
rect 35916 33156 35920 33212
rect 35856 33152 35920 33156
rect 35936 33212 36000 33216
rect 35936 33156 35940 33212
rect 35940 33156 35996 33212
rect 35996 33156 36000 33212
rect 35936 33152 36000 33156
rect 36016 33212 36080 33216
rect 36016 33156 36020 33212
rect 36020 33156 36076 33212
rect 36076 33156 36080 33212
rect 36016 33152 36080 33156
rect 36096 33212 36160 33216
rect 36096 33156 36100 33212
rect 36100 33156 36156 33212
rect 36156 33156 36160 33212
rect 36096 33152 36160 33156
rect 66576 33212 66640 33216
rect 66576 33156 66580 33212
rect 66580 33156 66636 33212
rect 66636 33156 66640 33212
rect 66576 33152 66640 33156
rect 66656 33212 66720 33216
rect 66656 33156 66660 33212
rect 66660 33156 66716 33212
rect 66716 33156 66720 33212
rect 66656 33152 66720 33156
rect 66736 33212 66800 33216
rect 66736 33156 66740 33212
rect 66740 33156 66796 33212
rect 66796 33156 66800 33212
rect 66736 33152 66800 33156
rect 66816 33212 66880 33216
rect 66816 33156 66820 33212
rect 66820 33156 66876 33212
rect 66876 33156 66880 33212
rect 66816 33152 66880 33156
rect 5796 32668 5860 32672
rect 5796 32612 5800 32668
rect 5800 32612 5856 32668
rect 5856 32612 5860 32668
rect 5796 32608 5860 32612
rect 5876 32668 5940 32672
rect 5876 32612 5880 32668
rect 5880 32612 5936 32668
rect 5936 32612 5940 32668
rect 5876 32608 5940 32612
rect 5956 32668 6020 32672
rect 5956 32612 5960 32668
rect 5960 32612 6016 32668
rect 6016 32612 6020 32668
rect 5956 32608 6020 32612
rect 6036 32668 6100 32672
rect 6036 32612 6040 32668
rect 6040 32612 6096 32668
rect 6096 32612 6100 32668
rect 6036 32608 6100 32612
rect 36516 32668 36580 32672
rect 36516 32612 36520 32668
rect 36520 32612 36576 32668
rect 36576 32612 36580 32668
rect 36516 32608 36580 32612
rect 36596 32668 36660 32672
rect 36596 32612 36600 32668
rect 36600 32612 36656 32668
rect 36656 32612 36660 32668
rect 36596 32608 36660 32612
rect 36676 32668 36740 32672
rect 36676 32612 36680 32668
rect 36680 32612 36736 32668
rect 36736 32612 36740 32668
rect 36676 32608 36740 32612
rect 36756 32668 36820 32672
rect 36756 32612 36760 32668
rect 36760 32612 36816 32668
rect 36816 32612 36820 32668
rect 36756 32608 36820 32612
rect 67236 32668 67300 32672
rect 67236 32612 67240 32668
rect 67240 32612 67296 32668
rect 67296 32612 67300 32668
rect 67236 32608 67300 32612
rect 67316 32668 67380 32672
rect 67316 32612 67320 32668
rect 67320 32612 67376 32668
rect 67376 32612 67380 32668
rect 67316 32608 67380 32612
rect 67396 32668 67460 32672
rect 67396 32612 67400 32668
rect 67400 32612 67456 32668
rect 67456 32612 67460 32668
rect 67396 32608 67460 32612
rect 67476 32668 67540 32672
rect 67476 32612 67480 32668
rect 67480 32612 67536 32668
rect 67536 32612 67540 32668
rect 67476 32608 67540 32612
rect 5136 32124 5200 32128
rect 5136 32068 5140 32124
rect 5140 32068 5196 32124
rect 5196 32068 5200 32124
rect 5136 32064 5200 32068
rect 5216 32124 5280 32128
rect 5216 32068 5220 32124
rect 5220 32068 5276 32124
rect 5276 32068 5280 32124
rect 5216 32064 5280 32068
rect 5296 32124 5360 32128
rect 5296 32068 5300 32124
rect 5300 32068 5356 32124
rect 5356 32068 5360 32124
rect 5296 32064 5360 32068
rect 5376 32124 5440 32128
rect 5376 32068 5380 32124
rect 5380 32068 5436 32124
rect 5436 32068 5440 32124
rect 5376 32064 5440 32068
rect 35856 32124 35920 32128
rect 35856 32068 35860 32124
rect 35860 32068 35916 32124
rect 35916 32068 35920 32124
rect 35856 32064 35920 32068
rect 35936 32124 36000 32128
rect 35936 32068 35940 32124
rect 35940 32068 35996 32124
rect 35996 32068 36000 32124
rect 35936 32064 36000 32068
rect 36016 32124 36080 32128
rect 36016 32068 36020 32124
rect 36020 32068 36076 32124
rect 36076 32068 36080 32124
rect 36016 32064 36080 32068
rect 36096 32124 36160 32128
rect 36096 32068 36100 32124
rect 36100 32068 36156 32124
rect 36156 32068 36160 32124
rect 36096 32064 36160 32068
rect 66576 32124 66640 32128
rect 66576 32068 66580 32124
rect 66580 32068 66636 32124
rect 66636 32068 66640 32124
rect 66576 32064 66640 32068
rect 66656 32124 66720 32128
rect 66656 32068 66660 32124
rect 66660 32068 66716 32124
rect 66716 32068 66720 32124
rect 66656 32064 66720 32068
rect 66736 32124 66800 32128
rect 66736 32068 66740 32124
rect 66740 32068 66796 32124
rect 66796 32068 66800 32124
rect 66736 32064 66800 32068
rect 66816 32124 66880 32128
rect 66816 32068 66820 32124
rect 66820 32068 66876 32124
rect 66876 32068 66880 32124
rect 66816 32064 66880 32068
rect 5796 31580 5860 31584
rect 5796 31524 5800 31580
rect 5800 31524 5856 31580
rect 5856 31524 5860 31580
rect 5796 31520 5860 31524
rect 5876 31580 5940 31584
rect 5876 31524 5880 31580
rect 5880 31524 5936 31580
rect 5936 31524 5940 31580
rect 5876 31520 5940 31524
rect 5956 31580 6020 31584
rect 5956 31524 5960 31580
rect 5960 31524 6016 31580
rect 6016 31524 6020 31580
rect 5956 31520 6020 31524
rect 6036 31580 6100 31584
rect 6036 31524 6040 31580
rect 6040 31524 6096 31580
rect 6096 31524 6100 31580
rect 6036 31520 6100 31524
rect 36516 31580 36580 31584
rect 36516 31524 36520 31580
rect 36520 31524 36576 31580
rect 36576 31524 36580 31580
rect 36516 31520 36580 31524
rect 36596 31580 36660 31584
rect 36596 31524 36600 31580
rect 36600 31524 36656 31580
rect 36656 31524 36660 31580
rect 36596 31520 36660 31524
rect 36676 31580 36740 31584
rect 36676 31524 36680 31580
rect 36680 31524 36736 31580
rect 36736 31524 36740 31580
rect 36676 31520 36740 31524
rect 36756 31580 36820 31584
rect 36756 31524 36760 31580
rect 36760 31524 36816 31580
rect 36816 31524 36820 31580
rect 36756 31520 36820 31524
rect 67236 31580 67300 31584
rect 67236 31524 67240 31580
rect 67240 31524 67296 31580
rect 67296 31524 67300 31580
rect 67236 31520 67300 31524
rect 67316 31580 67380 31584
rect 67316 31524 67320 31580
rect 67320 31524 67376 31580
rect 67376 31524 67380 31580
rect 67316 31520 67380 31524
rect 67396 31580 67460 31584
rect 67396 31524 67400 31580
rect 67400 31524 67456 31580
rect 67456 31524 67460 31580
rect 67396 31520 67460 31524
rect 67476 31580 67540 31584
rect 67476 31524 67480 31580
rect 67480 31524 67536 31580
rect 67536 31524 67540 31580
rect 67476 31520 67540 31524
rect 5136 31036 5200 31040
rect 5136 30980 5140 31036
rect 5140 30980 5196 31036
rect 5196 30980 5200 31036
rect 5136 30976 5200 30980
rect 5216 31036 5280 31040
rect 5216 30980 5220 31036
rect 5220 30980 5276 31036
rect 5276 30980 5280 31036
rect 5216 30976 5280 30980
rect 5296 31036 5360 31040
rect 5296 30980 5300 31036
rect 5300 30980 5356 31036
rect 5356 30980 5360 31036
rect 5296 30976 5360 30980
rect 5376 31036 5440 31040
rect 5376 30980 5380 31036
rect 5380 30980 5436 31036
rect 5436 30980 5440 31036
rect 5376 30976 5440 30980
rect 35856 31036 35920 31040
rect 35856 30980 35860 31036
rect 35860 30980 35916 31036
rect 35916 30980 35920 31036
rect 35856 30976 35920 30980
rect 35936 31036 36000 31040
rect 35936 30980 35940 31036
rect 35940 30980 35996 31036
rect 35996 30980 36000 31036
rect 35936 30976 36000 30980
rect 36016 31036 36080 31040
rect 36016 30980 36020 31036
rect 36020 30980 36076 31036
rect 36076 30980 36080 31036
rect 36016 30976 36080 30980
rect 36096 31036 36160 31040
rect 36096 30980 36100 31036
rect 36100 30980 36156 31036
rect 36156 30980 36160 31036
rect 36096 30976 36160 30980
rect 66576 31036 66640 31040
rect 66576 30980 66580 31036
rect 66580 30980 66636 31036
rect 66636 30980 66640 31036
rect 66576 30976 66640 30980
rect 66656 31036 66720 31040
rect 66656 30980 66660 31036
rect 66660 30980 66716 31036
rect 66716 30980 66720 31036
rect 66656 30976 66720 30980
rect 66736 31036 66800 31040
rect 66736 30980 66740 31036
rect 66740 30980 66796 31036
rect 66796 30980 66800 31036
rect 66736 30976 66800 30980
rect 66816 31036 66880 31040
rect 66816 30980 66820 31036
rect 66820 30980 66876 31036
rect 66876 30980 66880 31036
rect 66816 30976 66880 30980
rect 5796 30492 5860 30496
rect 5796 30436 5800 30492
rect 5800 30436 5856 30492
rect 5856 30436 5860 30492
rect 5796 30432 5860 30436
rect 5876 30492 5940 30496
rect 5876 30436 5880 30492
rect 5880 30436 5936 30492
rect 5936 30436 5940 30492
rect 5876 30432 5940 30436
rect 5956 30492 6020 30496
rect 5956 30436 5960 30492
rect 5960 30436 6016 30492
rect 6016 30436 6020 30492
rect 5956 30432 6020 30436
rect 6036 30492 6100 30496
rect 6036 30436 6040 30492
rect 6040 30436 6096 30492
rect 6096 30436 6100 30492
rect 6036 30432 6100 30436
rect 36516 30492 36580 30496
rect 36516 30436 36520 30492
rect 36520 30436 36576 30492
rect 36576 30436 36580 30492
rect 36516 30432 36580 30436
rect 36596 30492 36660 30496
rect 36596 30436 36600 30492
rect 36600 30436 36656 30492
rect 36656 30436 36660 30492
rect 36596 30432 36660 30436
rect 36676 30492 36740 30496
rect 36676 30436 36680 30492
rect 36680 30436 36736 30492
rect 36736 30436 36740 30492
rect 36676 30432 36740 30436
rect 36756 30492 36820 30496
rect 36756 30436 36760 30492
rect 36760 30436 36816 30492
rect 36816 30436 36820 30492
rect 36756 30432 36820 30436
rect 67236 30492 67300 30496
rect 67236 30436 67240 30492
rect 67240 30436 67296 30492
rect 67296 30436 67300 30492
rect 67236 30432 67300 30436
rect 67316 30492 67380 30496
rect 67316 30436 67320 30492
rect 67320 30436 67376 30492
rect 67376 30436 67380 30492
rect 67316 30432 67380 30436
rect 67396 30492 67460 30496
rect 67396 30436 67400 30492
rect 67400 30436 67456 30492
rect 67456 30436 67460 30492
rect 67396 30432 67460 30436
rect 67476 30492 67540 30496
rect 67476 30436 67480 30492
rect 67480 30436 67536 30492
rect 67536 30436 67540 30492
rect 67476 30432 67540 30436
rect 5136 29948 5200 29952
rect 5136 29892 5140 29948
rect 5140 29892 5196 29948
rect 5196 29892 5200 29948
rect 5136 29888 5200 29892
rect 5216 29948 5280 29952
rect 5216 29892 5220 29948
rect 5220 29892 5276 29948
rect 5276 29892 5280 29948
rect 5216 29888 5280 29892
rect 5296 29948 5360 29952
rect 5296 29892 5300 29948
rect 5300 29892 5356 29948
rect 5356 29892 5360 29948
rect 5296 29888 5360 29892
rect 5376 29948 5440 29952
rect 5376 29892 5380 29948
rect 5380 29892 5436 29948
rect 5436 29892 5440 29948
rect 5376 29888 5440 29892
rect 35856 29948 35920 29952
rect 35856 29892 35860 29948
rect 35860 29892 35916 29948
rect 35916 29892 35920 29948
rect 35856 29888 35920 29892
rect 35936 29948 36000 29952
rect 35936 29892 35940 29948
rect 35940 29892 35996 29948
rect 35996 29892 36000 29948
rect 35936 29888 36000 29892
rect 36016 29948 36080 29952
rect 36016 29892 36020 29948
rect 36020 29892 36076 29948
rect 36076 29892 36080 29948
rect 36016 29888 36080 29892
rect 36096 29948 36160 29952
rect 36096 29892 36100 29948
rect 36100 29892 36156 29948
rect 36156 29892 36160 29948
rect 36096 29888 36160 29892
rect 66576 29948 66640 29952
rect 66576 29892 66580 29948
rect 66580 29892 66636 29948
rect 66636 29892 66640 29948
rect 66576 29888 66640 29892
rect 66656 29948 66720 29952
rect 66656 29892 66660 29948
rect 66660 29892 66716 29948
rect 66716 29892 66720 29948
rect 66656 29888 66720 29892
rect 66736 29948 66800 29952
rect 66736 29892 66740 29948
rect 66740 29892 66796 29948
rect 66796 29892 66800 29948
rect 66736 29888 66800 29892
rect 66816 29948 66880 29952
rect 66816 29892 66820 29948
rect 66820 29892 66876 29948
rect 66876 29892 66880 29948
rect 66816 29888 66880 29892
rect 27476 29548 27540 29612
rect 5796 29404 5860 29408
rect 5796 29348 5800 29404
rect 5800 29348 5856 29404
rect 5856 29348 5860 29404
rect 5796 29344 5860 29348
rect 5876 29404 5940 29408
rect 5876 29348 5880 29404
rect 5880 29348 5936 29404
rect 5936 29348 5940 29404
rect 5876 29344 5940 29348
rect 5956 29404 6020 29408
rect 5956 29348 5960 29404
rect 5960 29348 6016 29404
rect 6016 29348 6020 29404
rect 5956 29344 6020 29348
rect 6036 29404 6100 29408
rect 6036 29348 6040 29404
rect 6040 29348 6096 29404
rect 6096 29348 6100 29404
rect 6036 29344 6100 29348
rect 36516 29404 36580 29408
rect 36516 29348 36520 29404
rect 36520 29348 36576 29404
rect 36576 29348 36580 29404
rect 36516 29344 36580 29348
rect 36596 29404 36660 29408
rect 36596 29348 36600 29404
rect 36600 29348 36656 29404
rect 36656 29348 36660 29404
rect 36596 29344 36660 29348
rect 36676 29404 36740 29408
rect 36676 29348 36680 29404
rect 36680 29348 36736 29404
rect 36736 29348 36740 29404
rect 36676 29344 36740 29348
rect 36756 29404 36820 29408
rect 36756 29348 36760 29404
rect 36760 29348 36816 29404
rect 36816 29348 36820 29404
rect 36756 29344 36820 29348
rect 67236 29404 67300 29408
rect 67236 29348 67240 29404
rect 67240 29348 67296 29404
rect 67296 29348 67300 29404
rect 67236 29344 67300 29348
rect 67316 29404 67380 29408
rect 67316 29348 67320 29404
rect 67320 29348 67376 29404
rect 67376 29348 67380 29404
rect 67316 29344 67380 29348
rect 67396 29404 67460 29408
rect 67396 29348 67400 29404
rect 67400 29348 67456 29404
rect 67456 29348 67460 29404
rect 67396 29344 67460 29348
rect 67476 29404 67540 29408
rect 67476 29348 67480 29404
rect 67480 29348 67536 29404
rect 67536 29348 67540 29404
rect 67476 29344 67540 29348
rect 5136 28860 5200 28864
rect 5136 28804 5140 28860
rect 5140 28804 5196 28860
rect 5196 28804 5200 28860
rect 5136 28800 5200 28804
rect 5216 28860 5280 28864
rect 5216 28804 5220 28860
rect 5220 28804 5276 28860
rect 5276 28804 5280 28860
rect 5216 28800 5280 28804
rect 5296 28860 5360 28864
rect 5296 28804 5300 28860
rect 5300 28804 5356 28860
rect 5356 28804 5360 28860
rect 5296 28800 5360 28804
rect 5376 28860 5440 28864
rect 5376 28804 5380 28860
rect 5380 28804 5436 28860
rect 5436 28804 5440 28860
rect 5376 28800 5440 28804
rect 35856 28860 35920 28864
rect 35856 28804 35860 28860
rect 35860 28804 35916 28860
rect 35916 28804 35920 28860
rect 35856 28800 35920 28804
rect 35936 28860 36000 28864
rect 35936 28804 35940 28860
rect 35940 28804 35996 28860
rect 35996 28804 36000 28860
rect 35936 28800 36000 28804
rect 36016 28860 36080 28864
rect 36016 28804 36020 28860
rect 36020 28804 36076 28860
rect 36076 28804 36080 28860
rect 36016 28800 36080 28804
rect 36096 28860 36160 28864
rect 36096 28804 36100 28860
rect 36100 28804 36156 28860
rect 36156 28804 36160 28860
rect 36096 28800 36160 28804
rect 66576 28860 66640 28864
rect 66576 28804 66580 28860
rect 66580 28804 66636 28860
rect 66636 28804 66640 28860
rect 66576 28800 66640 28804
rect 66656 28860 66720 28864
rect 66656 28804 66660 28860
rect 66660 28804 66716 28860
rect 66716 28804 66720 28860
rect 66656 28800 66720 28804
rect 66736 28860 66800 28864
rect 66736 28804 66740 28860
rect 66740 28804 66796 28860
rect 66796 28804 66800 28860
rect 66736 28800 66800 28804
rect 66816 28860 66880 28864
rect 66816 28804 66820 28860
rect 66820 28804 66876 28860
rect 66876 28804 66880 28860
rect 66816 28800 66880 28804
rect 5796 28316 5860 28320
rect 5796 28260 5800 28316
rect 5800 28260 5856 28316
rect 5856 28260 5860 28316
rect 5796 28256 5860 28260
rect 5876 28316 5940 28320
rect 5876 28260 5880 28316
rect 5880 28260 5936 28316
rect 5936 28260 5940 28316
rect 5876 28256 5940 28260
rect 5956 28316 6020 28320
rect 5956 28260 5960 28316
rect 5960 28260 6016 28316
rect 6016 28260 6020 28316
rect 5956 28256 6020 28260
rect 6036 28316 6100 28320
rect 6036 28260 6040 28316
rect 6040 28260 6096 28316
rect 6096 28260 6100 28316
rect 6036 28256 6100 28260
rect 36516 28316 36580 28320
rect 36516 28260 36520 28316
rect 36520 28260 36576 28316
rect 36576 28260 36580 28316
rect 36516 28256 36580 28260
rect 36596 28316 36660 28320
rect 36596 28260 36600 28316
rect 36600 28260 36656 28316
rect 36656 28260 36660 28316
rect 36596 28256 36660 28260
rect 36676 28316 36740 28320
rect 36676 28260 36680 28316
rect 36680 28260 36736 28316
rect 36736 28260 36740 28316
rect 36676 28256 36740 28260
rect 36756 28316 36820 28320
rect 36756 28260 36760 28316
rect 36760 28260 36816 28316
rect 36816 28260 36820 28316
rect 36756 28256 36820 28260
rect 67236 28316 67300 28320
rect 67236 28260 67240 28316
rect 67240 28260 67296 28316
rect 67296 28260 67300 28316
rect 67236 28256 67300 28260
rect 67316 28316 67380 28320
rect 67316 28260 67320 28316
rect 67320 28260 67376 28316
rect 67376 28260 67380 28316
rect 67316 28256 67380 28260
rect 67396 28316 67460 28320
rect 67396 28260 67400 28316
rect 67400 28260 67456 28316
rect 67456 28260 67460 28316
rect 67396 28256 67460 28260
rect 67476 28316 67540 28320
rect 67476 28260 67480 28316
rect 67480 28260 67536 28316
rect 67536 28260 67540 28316
rect 67476 28256 67540 28260
rect 5136 27772 5200 27776
rect 5136 27716 5140 27772
rect 5140 27716 5196 27772
rect 5196 27716 5200 27772
rect 5136 27712 5200 27716
rect 5216 27772 5280 27776
rect 5216 27716 5220 27772
rect 5220 27716 5276 27772
rect 5276 27716 5280 27772
rect 5216 27712 5280 27716
rect 5296 27772 5360 27776
rect 5296 27716 5300 27772
rect 5300 27716 5356 27772
rect 5356 27716 5360 27772
rect 5296 27712 5360 27716
rect 5376 27772 5440 27776
rect 5376 27716 5380 27772
rect 5380 27716 5436 27772
rect 5436 27716 5440 27772
rect 5376 27712 5440 27716
rect 35856 27772 35920 27776
rect 35856 27716 35860 27772
rect 35860 27716 35916 27772
rect 35916 27716 35920 27772
rect 35856 27712 35920 27716
rect 35936 27772 36000 27776
rect 35936 27716 35940 27772
rect 35940 27716 35996 27772
rect 35996 27716 36000 27772
rect 35936 27712 36000 27716
rect 36016 27772 36080 27776
rect 36016 27716 36020 27772
rect 36020 27716 36076 27772
rect 36076 27716 36080 27772
rect 36016 27712 36080 27716
rect 36096 27772 36160 27776
rect 36096 27716 36100 27772
rect 36100 27716 36156 27772
rect 36156 27716 36160 27772
rect 36096 27712 36160 27716
rect 66576 27772 66640 27776
rect 66576 27716 66580 27772
rect 66580 27716 66636 27772
rect 66636 27716 66640 27772
rect 66576 27712 66640 27716
rect 66656 27772 66720 27776
rect 66656 27716 66660 27772
rect 66660 27716 66716 27772
rect 66716 27716 66720 27772
rect 66656 27712 66720 27716
rect 66736 27772 66800 27776
rect 66736 27716 66740 27772
rect 66740 27716 66796 27772
rect 66796 27716 66800 27772
rect 66736 27712 66800 27716
rect 66816 27772 66880 27776
rect 66816 27716 66820 27772
rect 66820 27716 66876 27772
rect 66876 27716 66880 27772
rect 66816 27712 66880 27716
rect 5796 27228 5860 27232
rect 5796 27172 5800 27228
rect 5800 27172 5856 27228
rect 5856 27172 5860 27228
rect 5796 27168 5860 27172
rect 5876 27228 5940 27232
rect 5876 27172 5880 27228
rect 5880 27172 5936 27228
rect 5936 27172 5940 27228
rect 5876 27168 5940 27172
rect 5956 27228 6020 27232
rect 5956 27172 5960 27228
rect 5960 27172 6016 27228
rect 6016 27172 6020 27228
rect 5956 27168 6020 27172
rect 6036 27228 6100 27232
rect 6036 27172 6040 27228
rect 6040 27172 6096 27228
rect 6096 27172 6100 27228
rect 6036 27168 6100 27172
rect 36516 27228 36580 27232
rect 36516 27172 36520 27228
rect 36520 27172 36576 27228
rect 36576 27172 36580 27228
rect 36516 27168 36580 27172
rect 36596 27228 36660 27232
rect 36596 27172 36600 27228
rect 36600 27172 36656 27228
rect 36656 27172 36660 27228
rect 36596 27168 36660 27172
rect 36676 27228 36740 27232
rect 36676 27172 36680 27228
rect 36680 27172 36736 27228
rect 36736 27172 36740 27228
rect 36676 27168 36740 27172
rect 36756 27228 36820 27232
rect 36756 27172 36760 27228
rect 36760 27172 36816 27228
rect 36816 27172 36820 27228
rect 36756 27168 36820 27172
rect 67236 27228 67300 27232
rect 67236 27172 67240 27228
rect 67240 27172 67296 27228
rect 67296 27172 67300 27228
rect 67236 27168 67300 27172
rect 67316 27228 67380 27232
rect 67316 27172 67320 27228
rect 67320 27172 67376 27228
rect 67376 27172 67380 27228
rect 67316 27168 67380 27172
rect 67396 27228 67460 27232
rect 67396 27172 67400 27228
rect 67400 27172 67456 27228
rect 67456 27172 67460 27228
rect 67396 27168 67460 27172
rect 67476 27228 67540 27232
rect 67476 27172 67480 27228
rect 67480 27172 67536 27228
rect 67536 27172 67540 27228
rect 67476 27168 67540 27172
rect 28396 26828 28460 26892
rect 5136 26684 5200 26688
rect 5136 26628 5140 26684
rect 5140 26628 5196 26684
rect 5196 26628 5200 26684
rect 5136 26624 5200 26628
rect 5216 26684 5280 26688
rect 5216 26628 5220 26684
rect 5220 26628 5276 26684
rect 5276 26628 5280 26684
rect 5216 26624 5280 26628
rect 5296 26684 5360 26688
rect 5296 26628 5300 26684
rect 5300 26628 5356 26684
rect 5356 26628 5360 26684
rect 5296 26624 5360 26628
rect 5376 26684 5440 26688
rect 5376 26628 5380 26684
rect 5380 26628 5436 26684
rect 5436 26628 5440 26684
rect 5376 26624 5440 26628
rect 35856 26684 35920 26688
rect 35856 26628 35860 26684
rect 35860 26628 35916 26684
rect 35916 26628 35920 26684
rect 35856 26624 35920 26628
rect 35936 26684 36000 26688
rect 35936 26628 35940 26684
rect 35940 26628 35996 26684
rect 35996 26628 36000 26684
rect 35936 26624 36000 26628
rect 36016 26684 36080 26688
rect 36016 26628 36020 26684
rect 36020 26628 36076 26684
rect 36076 26628 36080 26684
rect 36016 26624 36080 26628
rect 36096 26684 36160 26688
rect 36096 26628 36100 26684
rect 36100 26628 36156 26684
rect 36156 26628 36160 26684
rect 36096 26624 36160 26628
rect 66576 26684 66640 26688
rect 66576 26628 66580 26684
rect 66580 26628 66636 26684
rect 66636 26628 66640 26684
rect 66576 26624 66640 26628
rect 66656 26684 66720 26688
rect 66656 26628 66660 26684
rect 66660 26628 66716 26684
rect 66716 26628 66720 26684
rect 66656 26624 66720 26628
rect 66736 26684 66800 26688
rect 66736 26628 66740 26684
rect 66740 26628 66796 26684
rect 66796 26628 66800 26684
rect 66736 26624 66800 26628
rect 66816 26684 66880 26688
rect 66816 26628 66820 26684
rect 66820 26628 66876 26684
rect 66876 26628 66880 26684
rect 66816 26624 66880 26628
rect 5796 26140 5860 26144
rect 5796 26084 5800 26140
rect 5800 26084 5856 26140
rect 5856 26084 5860 26140
rect 5796 26080 5860 26084
rect 5876 26140 5940 26144
rect 5876 26084 5880 26140
rect 5880 26084 5936 26140
rect 5936 26084 5940 26140
rect 5876 26080 5940 26084
rect 5956 26140 6020 26144
rect 5956 26084 5960 26140
rect 5960 26084 6016 26140
rect 6016 26084 6020 26140
rect 5956 26080 6020 26084
rect 6036 26140 6100 26144
rect 6036 26084 6040 26140
rect 6040 26084 6096 26140
rect 6096 26084 6100 26140
rect 6036 26080 6100 26084
rect 36516 26140 36580 26144
rect 36516 26084 36520 26140
rect 36520 26084 36576 26140
rect 36576 26084 36580 26140
rect 36516 26080 36580 26084
rect 36596 26140 36660 26144
rect 36596 26084 36600 26140
rect 36600 26084 36656 26140
rect 36656 26084 36660 26140
rect 36596 26080 36660 26084
rect 36676 26140 36740 26144
rect 36676 26084 36680 26140
rect 36680 26084 36736 26140
rect 36736 26084 36740 26140
rect 36676 26080 36740 26084
rect 36756 26140 36820 26144
rect 36756 26084 36760 26140
rect 36760 26084 36816 26140
rect 36816 26084 36820 26140
rect 36756 26080 36820 26084
rect 67236 26140 67300 26144
rect 67236 26084 67240 26140
rect 67240 26084 67296 26140
rect 67296 26084 67300 26140
rect 67236 26080 67300 26084
rect 67316 26140 67380 26144
rect 67316 26084 67320 26140
rect 67320 26084 67376 26140
rect 67376 26084 67380 26140
rect 67316 26080 67380 26084
rect 67396 26140 67460 26144
rect 67396 26084 67400 26140
rect 67400 26084 67456 26140
rect 67456 26084 67460 26140
rect 67396 26080 67460 26084
rect 67476 26140 67540 26144
rect 67476 26084 67480 26140
rect 67480 26084 67536 26140
rect 67536 26084 67540 26140
rect 67476 26080 67540 26084
rect 5136 25596 5200 25600
rect 5136 25540 5140 25596
rect 5140 25540 5196 25596
rect 5196 25540 5200 25596
rect 5136 25536 5200 25540
rect 5216 25596 5280 25600
rect 5216 25540 5220 25596
rect 5220 25540 5276 25596
rect 5276 25540 5280 25596
rect 5216 25536 5280 25540
rect 5296 25596 5360 25600
rect 5296 25540 5300 25596
rect 5300 25540 5356 25596
rect 5356 25540 5360 25596
rect 5296 25536 5360 25540
rect 5376 25596 5440 25600
rect 5376 25540 5380 25596
rect 5380 25540 5436 25596
rect 5436 25540 5440 25596
rect 5376 25536 5440 25540
rect 35856 25596 35920 25600
rect 35856 25540 35860 25596
rect 35860 25540 35916 25596
rect 35916 25540 35920 25596
rect 35856 25536 35920 25540
rect 35936 25596 36000 25600
rect 35936 25540 35940 25596
rect 35940 25540 35996 25596
rect 35996 25540 36000 25596
rect 35936 25536 36000 25540
rect 36016 25596 36080 25600
rect 36016 25540 36020 25596
rect 36020 25540 36076 25596
rect 36076 25540 36080 25596
rect 36016 25536 36080 25540
rect 36096 25596 36160 25600
rect 36096 25540 36100 25596
rect 36100 25540 36156 25596
rect 36156 25540 36160 25596
rect 36096 25536 36160 25540
rect 66576 25596 66640 25600
rect 66576 25540 66580 25596
rect 66580 25540 66636 25596
rect 66636 25540 66640 25596
rect 66576 25536 66640 25540
rect 66656 25596 66720 25600
rect 66656 25540 66660 25596
rect 66660 25540 66716 25596
rect 66716 25540 66720 25596
rect 66656 25536 66720 25540
rect 66736 25596 66800 25600
rect 66736 25540 66740 25596
rect 66740 25540 66796 25596
rect 66796 25540 66800 25596
rect 66736 25536 66800 25540
rect 66816 25596 66880 25600
rect 66816 25540 66820 25596
rect 66820 25540 66876 25596
rect 66876 25540 66880 25596
rect 66816 25536 66880 25540
rect 5796 25052 5860 25056
rect 5796 24996 5800 25052
rect 5800 24996 5856 25052
rect 5856 24996 5860 25052
rect 5796 24992 5860 24996
rect 5876 25052 5940 25056
rect 5876 24996 5880 25052
rect 5880 24996 5936 25052
rect 5936 24996 5940 25052
rect 5876 24992 5940 24996
rect 5956 25052 6020 25056
rect 5956 24996 5960 25052
rect 5960 24996 6016 25052
rect 6016 24996 6020 25052
rect 5956 24992 6020 24996
rect 6036 25052 6100 25056
rect 6036 24996 6040 25052
rect 6040 24996 6096 25052
rect 6096 24996 6100 25052
rect 6036 24992 6100 24996
rect 36516 25052 36580 25056
rect 36516 24996 36520 25052
rect 36520 24996 36576 25052
rect 36576 24996 36580 25052
rect 36516 24992 36580 24996
rect 36596 25052 36660 25056
rect 36596 24996 36600 25052
rect 36600 24996 36656 25052
rect 36656 24996 36660 25052
rect 36596 24992 36660 24996
rect 36676 25052 36740 25056
rect 36676 24996 36680 25052
rect 36680 24996 36736 25052
rect 36736 24996 36740 25052
rect 36676 24992 36740 24996
rect 36756 25052 36820 25056
rect 36756 24996 36760 25052
rect 36760 24996 36816 25052
rect 36816 24996 36820 25052
rect 36756 24992 36820 24996
rect 67236 25052 67300 25056
rect 67236 24996 67240 25052
rect 67240 24996 67296 25052
rect 67296 24996 67300 25052
rect 67236 24992 67300 24996
rect 67316 25052 67380 25056
rect 67316 24996 67320 25052
rect 67320 24996 67376 25052
rect 67376 24996 67380 25052
rect 67316 24992 67380 24996
rect 67396 25052 67460 25056
rect 67396 24996 67400 25052
rect 67400 24996 67456 25052
rect 67456 24996 67460 25052
rect 67396 24992 67460 24996
rect 67476 25052 67540 25056
rect 67476 24996 67480 25052
rect 67480 24996 67536 25052
rect 67536 24996 67540 25052
rect 67476 24992 67540 24996
rect 5136 24508 5200 24512
rect 5136 24452 5140 24508
rect 5140 24452 5196 24508
rect 5196 24452 5200 24508
rect 5136 24448 5200 24452
rect 5216 24508 5280 24512
rect 5216 24452 5220 24508
rect 5220 24452 5276 24508
rect 5276 24452 5280 24508
rect 5216 24448 5280 24452
rect 5296 24508 5360 24512
rect 5296 24452 5300 24508
rect 5300 24452 5356 24508
rect 5356 24452 5360 24508
rect 5296 24448 5360 24452
rect 5376 24508 5440 24512
rect 5376 24452 5380 24508
rect 5380 24452 5436 24508
rect 5436 24452 5440 24508
rect 5376 24448 5440 24452
rect 35856 24508 35920 24512
rect 35856 24452 35860 24508
rect 35860 24452 35916 24508
rect 35916 24452 35920 24508
rect 35856 24448 35920 24452
rect 35936 24508 36000 24512
rect 35936 24452 35940 24508
rect 35940 24452 35996 24508
rect 35996 24452 36000 24508
rect 35936 24448 36000 24452
rect 36016 24508 36080 24512
rect 36016 24452 36020 24508
rect 36020 24452 36076 24508
rect 36076 24452 36080 24508
rect 36016 24448 36080 24452
rect 36096 24508 36160 24512
rect 36096 24452 36100 24508
rect 36100 24452 36156 24508
rect 36156 24452 36160 24508
rect 36096 24448 36160 24452
rect 66576 24508 66640 24512
rect 66576 24452 66580 24508
rect 66580 24452 66636 24508
rect 66636 24452 66640 24508
rect 66576 24448 66640 24452
rect 66656 24508 66720 24512
rect 66656 24452 66660 24508
rect 66660 24452 66716 24508
rect 66716 24452 66720 24508
rect 66656 24448 66720 24452
rect 66736 24508 66800 24512
rect 66736 24452 66740 24508
rect 66740 24452 66796 24508
rect 66796 24452 66800 24508
rect 66736 24448 66800 24452
rect 66816 24508 66880 24512
rect 66816 24452 66820 24508
rect 66820 24452 66876 24508
rect 66876 24452 66880 24508
rect 66816 24448 66880 24452
rect 35020 24108 35084 24172
rect 5796 23964 5860 23968
rect 5796 23908 5800 23964
rect 5800 23908 5856 23964
rect 5856 23908 5860 23964
rect 5796 23904 5860 23908
rect 5876 23964 5940 23968
rect 5876 23908 5880 23964
rect 5880 23908 5936 23964
rect 5936 23908 5940 23964
rect 5876 23904 5940 23908
rect 5956 23964 6020 23968
rect 5956 23908 5960 23964
rect 5960 23908 6016 23964
rect 6016 23908 6020 23964
rect 5956 23904 6020 23908
rect 6036 23964 6100 23968
rect 6036 23908 6040 23964
rect 6040 23908 6096 23964
rect 6096 23908 6100 23964
rect 6036 23904 6100 23908
rect 36516 23964 36580 23968
rect 36516 23908 36520 23964
rect 36520 23908 36576 23964
rect 36576 23908 36580 23964
rect 36516 23904 36580 23908
rect 36596 23964 36660 23968
rect 36596 23908 36600 23964
rect 36600 23908 36656 23964
rect 36656 23908 36660 23964
rect 36596 23904 36660 23908
rect 36676 23964 36740 23968
rect 36676 23908 36680 23964
rect 36680 23908 36736 23964
rect 36736 23908 36740 23964
rect 36676 23904 36740 23908
rect 36756 23964 36820 23968
rect 36756 23908 36760 23964
rect 36760 23908 36816 23964
rect 36816 23908 36820 23964
rect 36756 23904 36820 23908
rect 67236 23964 67300 23968
rect 67236 23908 67240 23964
rect 67240 23908 67296 23964
rect 67296 23908 67300 23964
rect 67236 23904 67300 23908
rect 67316 23964 67380 23968
rect 67316 23908 67320 23964
rect 67320 23908 67376 23964
rect 67376 23908 67380 23964
rect 67316 23904 67380 23908
rect 67396 23964 67460 23968
rect 67396 23908 67400 23964
rect 67400 23908 67456 23964
rect 67456 23908 67460 23964
rect 67396 23904 67460 23908
rect 67476 23964 67540 23968
rect 67476 23908 67480 23964
rect 67480 23908 67536 23964
rect 67536 23908 67540 23964
rect 67476 23904 67540 23908
rect 5136 23420 5200 23424
rect 5136 23364 5140 23420
rect 5140 23364 5196 23420
rect 5196 23364 5200 23420
rect 5136 23360 5200 23364
rect 5216 23420 5280 23424
rect 5216 23364 5220 23420
rect 5220 23364 5276 23420
rect 5276 23364 5280 23420
rect 5216 23360 5280 23364
rect 5296 23420 5360 23424
rect 5296 23364 5300 23420
rect 5300 23364 5356 23420
rect 5356 23364 5360 23420
rect 5296 23360 5360 23364
rect 5376 23420 5440 23424
rect 5376 23364 5380 23420
rect 5380 23364 5436 23420
rect 5436 23364 5440 23420
rect 5376 23360 5440 23364
rect 35856 23420 35920 23424
rect 35856 23364 35860 23420
rect 35860 23364 35916 23420
rect 35916 23364 35920 23420
rect 35856 23360 35920 23364
rect 35936 23420 36000 23424
rect 35936 23364 35940 23420
rect 35940 23364 35996 23420
rect 35996 23364 36000 23420
rect 35936 23360 36000 23364
rect 36016 23420 36080 23424
rect 36016 23364 36020 23420
rect 36020 23364 36076 23420
rect 36076 23364 36080 23420
rect 36016 23360 36080 23364
rect 36096 23420 36160 23424
rect 36096 23364 36100 23420
rect 36100 23364 36156 23420
rect 36156 23364 36160 23420
rect 36096 23360 36160 23364
rect 66576 23420 66640 23424
rect 66576 23364 66580 23420
rect 66580 23364 66636 23420
rect 66636 23364 66640 23420
rect 66576 23360 66640 23364
rect 66656 23420 66720 23424
rect 66656 23364 66660 23420
rect 66660 23364 66716 23420
rect 66716 23364 66720 23420
rect 66656 23360 66720 23364
rect 66736 23420 66800 23424
rect 66736 23364 66740 23420
rect 66740 23364 66796 23420
rect 66796 23364 66800 23420
rect 66736 23360 66800 23364
rect 66816 23420 66880 23424
rect 66816 23364 66820 23420
rect 66820 23364 66876 23420
rect 66876 23364 66880 23420
rect 66816 23360 66880 23364
rect 5796 22876 5860 22880
rect 5796 22820 5800 22876
rect 5800 22820 5856 22876
rect 5856 22820 5860 22876
rect 5796 22816 5860 22820
rect 5876 22876 5940 22880
rect 5876 22820 5880 22876
rect 5880 22820 5936 22876
rect 5936 22820 5940 22876
rect 5876 22816 5940 22820
rect 5956 22876 6020 22880
rect 5956 22820 5960 22876
rect 5960 22820 6016 22876
rect 6016 22820 6020 22876
rect 5956 22816 6020 22820
rect 6036 22876 6100 22880
rect 6036 22820 6040 22876
rect 6040 22820 6096 22876
rect 6096 22820 6100 22876
rect 6036 22816 6100 22820
rect 36516 22876 36580 22880
rect 36516 22820 36520 22876
rect 36520 22820 36576 22876
rect 36576 22820 36580 22876
rect 36516 22816 36580 22820
rect 36596 22876 36660 22880
rect 36596 22820 36600 22876
rect 36600 22820 36656 22876
rect 36656 22820 36660 22876
rect 36596 22816 36660 22820
rect 36676 22876 36740 22880
rect 36676 22820 36680 22876
rect 36680 22820 36736 22876
rect 36736 22820 36740 22876
rect 36676 22816 36740 22820
rect 36756 22876 36820 22880
rect 36756 22820 36760 22876
rect 36760 22820 36816 22876
rect 36816 22820 36820 22876
rect 36756 22816 36820 22820
rect 67236 22876 67300 22880
rect 67236 22820 67240 22876
rect 67240 22820 67296 22876
rect 67296 22820 67300 22876
rect 67236 22816 67300 22820
rect 67316 22876 67380 22880
rect 67316 22820 67320 22876
rect 67320 22820 67376 22876
rect 67376 22820 67380 22876
rect 67316 22816 67380 22820
rect 67396 22876 67460 22880
rect 67396 22820 67400 22876
rect 67400 22820 67456 22876
rect 67456 22820 67460 22876
rect 67396 22816 67460 22820
rect 67476 22876 67540 22880
rect 67476 22820 67480 22876
rect 67480 22820 67536 22876
rect 67536 22820 67540 22876
rect 67476 22816 67540 22820
rect 5136 22332 5200 22336
rect 5136 22276 5140 22332
rect 5140 22276 5196 22332
rect 5196 22276 5200 22332
rect 5136 22272 5200 22276
rect 5216 22332 5280 22336
rect 5216 22276 5220 22332
rect 5220 22276 5276 22332
rect 5276 22276 5280 22332
rect 5216 22272 5280 22276
rect 5296 22332 5360 22336
rect 5296 22276 5300 22332
rect 5300 22276 5356 22332
rect 5356 22276 5360 22332
rect 5296 22272 5360 22276
rect 5376 22332 5440 22336
rect 5376 22276 5380 22332
rect 5380 22276 5436 22332
rect 5436 22276 5440 22332
rect 5376 22272 5440 22276
rect 35856 22332 35920 22336
rect 35856 22276 35860 22332
rect 35860 22276 35916 22332
rect 35916 22276 35920 22332
rect 35856 22272 35920 22276
rect 35936 22332 36000 22336
rect 35936 22276 35940 22332
rect 35940 22276 35996 22332
rect 35996 22276 36000 22332
rect 35936 22272 36000 22276
rect 36016 22332 36080 22336
rect 36016 22276 36020 22332
rect 36020 22276 36076 22332
rect 36076 22276 36080 22332
rect 36016 22272 36080 22276
rect 36096 22332 36160 22336
rect 36096 22276 36100 22332
rect 36100 22276 36156 22332
rect 36156 22276 36160 22332
rect 36096 22272 36160 22276
rect 66576 22332 66640 22336
rect 66576 22276 66580 22332
rect 66580 22276 66636 22332
rect 66636 22276 66640 22332
rect 66576 22272 66640 22276
rect 66656 22332 66720 22336
rect 66656 22276 66660 22332
rect 66660 22276 66716 22332
rect 66716 22276 66720 22332
rect 66656 22272 66720 22276
rect 66736 22332 66800 22336
rect 66736 22276 66740 22332
rect 66740 22276 66796 22332
rect 66796 22276 66800 22332
rect 66736 22272 66800 22276
rect 66816 22332 66880 22336
rect 66816 22276 66820 22332
rect 66820 22276 66876 22332
rect 66876 22276 66880 22332
rect 66816 22272 66880 22276
rect 5796 21788 5860 21792
rect 5796 21732 5800 21788
rect 5800 21732 5856 21788
rect 5856 21732 5860 21788
rect 5796 21728 5860 21732
rect 5876 21788 5940 21792
rect 5876 21732 5880 21788
rect 5880 21732 5936 21788
rect 5936 21732 5940 21788
rect 5876 21728 5940 21732
rect 5956 21788 6020 21792
rect 5956 21732 5960 21788
rect 5960 21732 6016 21788
rect 6016 21732 6020 21788
rect 5956 21728 6020 21732
rect 6036 21788 6100 21792
rect 6036 21732 6040 21788
rect 6040 21732 6096 21788
rect 6096 21732 6100 21788
rect 6036 21728 6100 21732
rect 36516 21788 36580 21792
rect 36516 21732 36520 21788
rect 36520 21732 36576 21788
rect 36576 21732 36580 21788
rect 36516 21728 36580 21732
rect 36596 21788 36660 21792
rect 36596 21732 36600 21788
rect 36600 21732 36656 21788
rect 36656 21732 36660 21788
rect 36596 21728 36660 21732
rect 36676 21788 36740 21792
rect 36676 21732 36680 21788
rect 36680 21732 36736 21788
rect 36736 21732 36740 21788
rect 36676 21728 36740 21732
rect 36756 21788 36820 21792
rect 36756 21732 36760 21788
rect 36760 21732 36816 21788
rect 36816 21732 36820 21788
rect 36756 21728 36820 21732
rect 67236 21788 67300 21792
rect 67236 21732 67240 21788
rect 67240 21732 67296 21788
rect 67296 21732 67300 21788
rect 67236 21728 67300 21732
rect 67316 21788 67380 21792
rect 67316 21732 67320 21788
rect 67320 21732 67376 21788
rect 67376 21732 67380 21788
rect 67316 21728 67380 21732
rect 67396 21788 67460 21792
rect 67396 21732 67400 21788
rect 67400 21732 67456 21788
rect 67456 21732 67460 21788
rect 67396 21728 67460 21732
rect 67476 21788 67540 21792
rect 67476 21732 67480 21788
rect 67480 21732 67536 21788
rect 67536 21732 67540 21788
rect 67476 21728 67540 21732
rect 5136 21244 5200 21248
rect 5136 21188 5140 21244
rect 5140 21188 5196 21244
rect 5196 21188 5200 21244
rect 5136 21184 5200 21188
rect 5216 21244 5280 21248
rect 5216 21188 5220 21244
rect 5220 21188 5276 21244
rect 5276 21188 5280 21244
rect 5216 21184 5280 21188
rect 5296 21244 5360 21248
rect 5296 21188 5300 21244
rect 5300 21188 5356 21244
rect 5356 21188 5360 21244
rect 5296 21184 5360 21188
rect 5376 21244 5440 21248
rect 5376 21188 5380 21244
rect 5380 21188 5436 21244
rect 5436 21188 5440 21244
rect 5376 21184 5440 21188
rect 35856 21244 35920 21248
rect 35856 21188 35860 21244
rect 35860 21188 35916 21244
rect 35916 21188 35920 21244
rect 35856 21184 35920 21188
rect 35936 21244 36000 21248
rect 35936 21188 35940 21244
rect 35940 21188 35996 21244
rect 35996 21188 36000 21244
rect 35936 21184 36000 21188
rect 36016 21244 36080 21248
rect 36016 21188 36020 21244
rect 36020 21188 36076 21244
rect 36076 21188 36080 21244
rect 36016 21184 36080 21188
rect 36096 21244 36160 21248
rect 36096 21188 36100 21244
rect 36100 21188 36156 21244
rect 36156 21188 36160 21244
rect 36096 21184 36160 21188
rect 66576 21244 66640 21248
rect 66576 21188 66580 21244
rect 66580 21188 66636 21244
rect 66636 21188 66640 21244
rect 66576 21184 66640 21188
rect 66656 21244 66720 21248
rect 66656 21188 66660 21244
rect 66660 21188 66716 21244
rect 66716 21188 66720 21244
rect 66656 21184 66720 21188
rect 66736 21244 66800 21248
rect 66736 21188 66740 21244
rect 66740 21188 66796 21244
rect 66796 21188 66800 21244
rect 66736 21184 66800 21188
rect 66816 21244 66880 21248
rect 66816 21188 66820 21244
rect 66820 21188 66876 21244
rect 66876 21188 66880 21244
rect 66816 21184 66880 21188
rect 5796 20700 5860 20704
rect 5796 20644 5800 20700
rect 5800 20644 5856 20700
rect 5856 20644 5860 20700
rect 5796 20640 5860 20644
rect 5876 20700 5940 20704
rect 5876 20644 5880 20700
rect 5880 20644 5936 20700
rect 5936 20644 5940 20700
rect 5876 20640 5940 20644
rect 5956 20700 6020 20704
rect 5956 20644 5960 20700
rect 5960 20644 6016 20700
rect 6016 20644 6020 20700
rect 5956 20640 6020 20644
rect 6036 20700 6100 20704
rect 6036 20644 6040 20700
rect 6040 20644 6096 20700
rect 6096 20644 6100 20700
rect 6036 20640 6100 20644
rect 36516 20700 36580 20704
rect 36516 20644 36520 20700
rect 36520 20644 36576 20700
rect 36576 20644 36580 20700
rect 36516 20640 36580 20644
rect 36596 20700 36660 20704
rect 36596 20644 36600 20700
rect 36600 20644 36656 20700
rect 36656 20644 36660 20700
rect 36596 20640 36660 20644
rect 36676 20700 36740 20704
rect 36676 20644 36680 20700
rect 36680 20644 36736 20700
rect 36736 20644 36740 20700
rect 36676 20640 36740 20644
rect 36756 20700 36820 20704
rect 36756 20644 36760 20700
rect 36760 20644 36816 20700
rect 36816 20644 36820 20700
rect 36756 20640 36820 20644
rect 67236 20700 67300 20704
rect 67236 20644 67240 20700
rect 67240 20644 67296 20700
rect 67296 20644 67300 20700
rect 67236 20640 67300 20644
rect 67316 20700 67380 20704
rect 67316 20644 67320 20700
rect 67320 20644 67376 20700
rect 67376 20644 67380 20700
rect 67316 20640 67380 20644
rect 67396 20700 67460 20704
rect 67396 20644 67400 20700
rect 67400 20644 67456 20700
rect 67456 20644 67460 20700
rect 67396 20640 67460 20644
rect 67476 20700 67540 20704
rect 67476 20644 67480 20700
rect 67480 20644 67536 20700
rect 67536 20644 67540 20700
rect 67476 20640 67540 20644
rect 5136 20156 5200 20160
rect 5136 20100 5140 20156
rect 5140 20100 5196 20156
rect 5196 20100 5200 20156
rect 5136 20096 5200 20100
rect 5216 20156 5280 20160
rect 5216 20100 5220 20156
rect 5220 20100 5276 20156
rect 5276 20100 5280 20156
rect 5216 20096 5280 20100
rect 5296 20156 5360 20160
rect 5296 20100 5300 20156
rect 5300 20100 5356 20156
rect 5356 20100 5360 20156
rect 5296 20096 5360 20100
rect 5376 20156 5440 20160
rect 5376 20100 5380 20156
rect 5380 20100 5436 20156
rect 5436 20100 5440 20156
rect 5376 20096 5440 20100
rect 35856 20156 35920 20160
rect 35856 20100 35860 20156
rect 35860 20100 35916 20156
rect 35916 20100 35920 20156
rect 35856 20096 35920 20100
rect 35936 20156 36000 20160
rect 35936 20100 35940 20156
rect 35940 20100 35996 20156
rect 35996 20100 36000 20156
rect 35936 20096 36000 20100
rect 36016 20156 36080 20160
rect 36016 20100 36020 20156
rect 36020 20100 36076 20156
rect 36076 20100 36080 20156
rect 36016 20096 36080 20100
rect 36096 20156 36160 20160
rect 36096 20100 36100 20156
rect 36100 20100 36156 20156
rect 36156 20100 36160 20156
rect 36096 20096 36160 20100
rect 66576 20156 66640 20160
rect 66576 20100 66580 20156
rect 66580 20100 66636 20156
rect 66636 20100 66640 20156
rect 66576 20096 66640 20100
rect 66656 20156 66720 20160
rect 66656 20100 66660 20156
rect 66660 20100 66716 20156
rect 66716 20100 66720 20156
rect 66656 20096 66720 20100
rect 66736 20156 66800 20160
rect 66736 20100 66740 20156
rect 66740 20100 66796 20156
rect 66796 20100 66800 20156
rect 66736 20096 66800 20100
rect 66816 20156 66880 20160
rect 66816 20100 66820 20156
rect 66820 20100 66876 20156
rect 66876 20100 66880 20156
rect 66816 20096 66880 20100
rect 5796 19612 5860 19616
rect 5796 19556 5800 19612
rect 5800 19556 5856 19612
rect 5856 19556 5860 19612
rect 5796 19552 5860 19556
rect 5876 19612 5940 19616
rect 5876 19556 5880 19612
rect 5880 19556 5936 19612
rect 5936 19556 5940 19612
rect 5876 19552 5940 19556
rect 5956 19612 6020 19616
rect 5956 19556 5960 19612
rect 5960 19556 6016 19612
rect 6016 19556 6020 19612
rect 5956 19552 6020 19556
rect 6036 19612 6100 19616
rect 6036 19556 6040 19612
rect 6040 19556 6096 19612
rect 6096 19556 6100 19612
rect 6036 19552 6100 19556
rect 36516 19612 36580 19616
rect 36516 19556 36520 19612
rect 36520 19556 36576 19612
rect 36576 19556 36580 19612
rect 36516 19552 36580 19556
rect 36596 19612 36660 19616
rect 36596 19556 36600 19612
rect 36600 19556 36656 19612
rect 36656 19556 36660 19612
rect 36596 19552 36660 19556
rect 36676 19612 36740 19616
rect 36676 19556 36680 19612
rect 36680 19556 36736 19612
rect 36736 19556 36740 19612
rect 36676 19552 36740 19556
rect 36756 19612 36820 19616
rect 36756 19556 36760 19612
rect 36760 19556 36816 19612
rect 36816 19556 36820 19612
rect 36756 19552 36820 19556
rect 67236 19612 67300 19616
rect 67236 19556 67240 19612
rect 67240 19556 67296 19612
rect 67296 19556 67300 19612
rect 67236 19552 67300 19556
rect 67316 19612 67380 19616
rect 67316 19556 67320 19612
rect 67320 19556 67376 19612
rect 67376 19556 67380 19612
rect 67316 19552 67380 19556
rect 67396 19612 67460 19616
rect 67396 19556 67400 19612
rect 67400 19556 67456 19612
rect 67456 19556 67460 19612
rect 67396 19552 67460 19556
rect 67476 19612 67540 19616
rect 67476 19556 67480 19612
rect 67480 19556 67536 19612
rect 67536 19556 67540 19612
rect 67476 19552 67540 19556
rect 5136 19068 5200 19072
rect 5136 19012 5140 19068
rect 5140 19012 5196 19068
rect 5196 19012 5200 19068
rect 5136 19008 5200 19012
rect 5216 19068 5280 19072
rect 5216 19012 5220 19068
rect 5220 19012 5276 19068
rect 5276 19012 5280 19068
rect 5216 19008 5280 19012
rect 5296 19068 5360 19072
rect 5296 19012 5300 19068
rect 5300 19012 5356 19068
rect 5356 19012 5360 19068
rect 5296 19008 5360 19012
rect 5376 19068 5440 19072
rect 5376 19012 5380 19068
rect 5380 19012 5436 19068
rect 5436 19012 5440 19068
rect 5376 19008 5440 19012
rect 35856 19068 35920 19072
rect 35856 19012 35860 19068
rect 35860 19012 35916 19068
rect 35916 19012 35920 19068
rect 35856 19008 35920 19012
rect 35936 19068 36000 19072
rect 35936 19012 35940 19068
rect 35940 19012 35996 19068
rect 35996 19012 36000 19068
rect 35936 19008 36000 19012
rect 36016 19068 36080 19072
rect 36016 19012 36020 19068
rect 36020 19012 36076 19068
rect 36076 19012 36080 19068
rect 36016 19008 36080 19012
rect 36096 19068 36160 19072
rect 36096 19012 36100 19068
rect 36100 19012 36156 19068
rect 36156 19012 36160 19068
rect 36096 19008 36160 19012
rect 66576 19068 66640 19072
rect 66576 19012 66580 19068
rect 66580 19012 66636 19068
rect 66636 19012 66640 19068
rect 66576 19008 66640 19012
rect 66656 19068 66720 19072
rect 66656 19012 66660 19068
rect 66660 19012 66716 19068
rect 66716 19012 66720 19068
rect 66656 19008 66720 19012
rect 66736 19068 66800 19072
rect 66736 19012 66740 19068
rect 66740 19012 66796 19068
rect 66796 19012 66800 19068
rect 66736 19008 66800 19012
rect 66816 19068 66880 19072
rect 66816 19012 66820 19068
rect 66820 19012 66876 19068
rect 66876 19012 66880 19068
rect 66816 19008 66880 19012
rect 5796 18524 5860 18528
rect 5796 18468 5800 18524
rect 5800 18468 5856 18524
rect 5856 18468 5860 18524
rect 5796 18464 5860 18468
rect 5876 18524 5940 18528
rect 5876 18468 5880 18524
rect 5880 18468 5936 18524
rect 5936 18468 5940 18524
rect 5876 18464 5940 18468
rect 5956 18524 6020 18528
rect 5956 18468 5960 18524
rect 5960 18468 6016 18524
rect 6016 18468 6020 18524
rect 5956 18464 6020 18468
rect 6036 18524 6100 18528
rect 6036 18468 6040 18524
rect 6040 18468 6096 18524
rect 6096 18468 6100 18524
rect 6036 18464 6100 18468
rect 36516 18524 36580 18528
rect 36516 18468 36520 18524
rect 36520 18468 36576 18524
rect 36576 18468 36580 18524
rect 36516 18464 36580 18468
rect 36596 18524 36660 18528
rect 36596 18468 36600 18524
rect 36600 18468 36656 18524
rect 36656 18468 36660 18524
rect 36596 18464 36660 18468
rect 36676 18524 36740 18528
rect 36676 18468 36680 18524
rect 36680 18468 36736 18524
rect 36736 18468 36740 18524
rect 36676 18464 36740 18468
rect 36756 18524 36820 18528
rect 36756 18468 36760 18524
rect 36760 18468 36816 18524
rect 36816 18468 36820 18524
rect 36756 18464 36820 18468
rect 67236 18524 67300 18528
rect 67236 18468 67240 18524
rect 67240 18468 67296 18524
rect 67296 18468 67300 18524
rect 67236 18464 67300 18468
rect 67316 18524 67380 18528
rect 67316 18468 67320 18524
rect 67320 18468 67376 18524
rect 67376 18468 67380 18524
rect 67316 18464 67380 18468
rect 67396 18524 67460 18528
rect 67396 18468 67400 18524
rect 67400 18468 67456 18524
rect 67456 18468 67460 18524
rect 67396 18464 67460 18468
rect 67476 18524 67540 18528
rect 67476 18468 67480 18524
rect 67480 18468 67536 18524
rect 67536 18468 67540 18524
rect 67476 18464 67540 18468
rect 27292 17988 27356 18052
rect 5136 17980 5200 17984
rect 5136 17924 5140 17980
rect 5140 17924 5196 17980
rect 5196 17924 5200 17980
rect 5136 17920 5200 17924
rect 5216 17980 5280 17984
rect 5216 17924 5220 17980
rect 5220 17924 5276 17980
rect 5276 17924 5280 17980
rect 5216 17920 5280 17924
rect 5296 17980 5360 17984
rect 5296 17924 5300 17980
rect 5300 17924 5356 17980
rect 5356 17924 5360 17980
rect 5296 17920 5360 17924
rect 5376 17980 5440 17984
rect 5376 17924 5380 17980
rect 5380 17924 5436 17980
rect 5436 17924 5440 17980
rect 5376 17920 5440 17924
rect 35856 17980 35920 17984
rect 35856 17924 35860 17980
rect 35860 17924 35916 17980
rect 35916 17924 35920 17980
rect 35856 17920 35920 17924
rect 35936 17980 36000 17984
rect 35936 17924 35940 17980
rect 35940 17924 35996 17980
rect 35996 17924 36000 17980
rect 35936 17920 36000 17924
rect 36016 17980 36080 17984
rect 36016 17924 36020 17980
rect 36020 17924 36076 17980
rect 36076 17924 36080 17980
rect 36016 17920 36080 17924
rect 36096 17980 36160 17984
rect 36096 17924 36100 17980
rect 36100 17924 36156 17980
rect 36156 17924 36160 17980
rect 36096 17920 36160 17924
rect 66576 17980 66640 17984
rect 66576 17924 66580 17980
rect 66580 17924 66636 17980
rect 66636 17924 66640 17980
rect 66576 17920 66640 17924
rect 66656 17980 66720 17984
rect 66656 17924 66660 17980
rect 66660 17924 66716 17980
rect 66716 17924 66720 17980
rect 66656 17920 66720 17924
rect 66736 17980 66800 17984
rect 66736 17924 66740 17980
rect 66740 17924 66796 17980
rect 66796 17924 66800 17980
rect 66736 17920 66800 17924
rect 66816 17980 66880 17984
rect 66816 17924 66820 17980
rect 66820 17924 66876 17980
rect 66876 17924 66880 17980
rect 66816 17920 66880 17924
rect 5796 17436 5860 17440
rect 5796 17380 5800 17436
rect 5800 17380 5856 17436
rect 5856 17380 5860 17436
rect 5796 17376 5860 17380
rect 5876 17436 5940 17440
rect 5876 17380 5880 17436
rect 5880 17380 5936 17436
rect 5936 17380 5940 17436
rect 5876 17376 5940 17380
rect 5956 17436 6020 17440
rect 5956 17380 5960 17436
rect 5960 17380 6016 17436
rect 6016 17380 6020 17436
rect 5956 17376 6020 17380
rect 6036 17436 6100 17440
rect 6036 17380 6040 17436
rect 6040 17380 6096 17436
rect 6096 17380 6100 17436
rect 6036 17376 6100 17380
rect 36516 17436 36580 17440
rect 36516 17380 36520 17436
rect 36520 17380 36576 17436
rect 36576 17380 36580 17436
rect 36516 17376 36580 17380
rect 36596 17436 36660 17440
rect 36596 17380 36600 17436
rect 36600 17380 36656 17436
rect 36656 17380 36660 17436
rect 36596 17376 36660 17380
rect 36676 17436 36740 17440
rect 36676 17380 36680 17436
rect 36680 17380 36736 17436
rect 36736 17380 36740 17436
rect 36676 17376 36740 17380
rect 36756 17436 36820 17440
rect 36756 17380 36760 17436
rect 36760 17380 36816 17436
rect 36816 17380 36820 17436
rect 36756 17376 36820 17380
rect 67236 17436 67300 17440
rect 67236 17380 67240 17436
rect 67240 17380 67296 17436
rect 67296 17380 67300 17436
rect 67236 17376 67300 17380
rect 67316 17436 67380 17440
rect 67316 17380 67320 17436
rect 67320 17380 67376 17436
rect 67376 17380 67380 17436
rect 67316 17376 67380 17380
rect 67396 17436 67460 17440
rect 67396 17380 67400 17436
rect 67400 17380 67456 17436
rect 67456 17380 67460 17436
rect 67396 17376 67460 17380
rect 67476 17436 67540 17440
rect 67476 17380 67480 17436
rect 67480 17380 67536 17436
rect 67536 17380 67540 17436
rect 67476 17376 67540 17380
rect 5136 16892 5200 16896
rect 5136 16836 5140 16892
rect 5140 16836 5196 16892
rect 5196 16836 5200 16892
rect 5136 16832 5200 16836
rect 5216 16892 5280 16896
rect 5216 16836 5220 16892
rect 5220 16836 5276 16892
rect 5276 16836 5280 16892
rect 5216 16832 5280 16836
rect 5296 16892 5360 16896
rect 5296 16836 5300 16892
rect 5300 16836 5356 16892
rect 5356 16836 5360 16892
rect 5296 16832 5360 16836
rect 5376 16892 5440 16896
rect 5376 16836 5380 16892
rect 5380 16836 5436 16892
rect 5436 16836 5440 16892
rect 5376 16832 5440 16836
rect 35856 16892 35920 16896
rect 35856 16836 35860 16892
rect 35860 16836 35916 16892
rect 35916 16836 35920 16892
rect 35856 16832 35920 16836
rect 35936 16892 36000 16896
rect 35936 16836 35940 16892
rect 35940 16836 35996 16892
rect 35996 16836 36000 16892
rect 35936 16832 36000 16836
rect 36016 16892 36080 16896
rect 36016 16836 36020 16892
rect 36020 16836 36076 16892
rect 36076 16836 36080 16892
rect 36016 16832 36080 16836
rect 36096 16892 36160 16896
rect 36096 16836 36100 16892
rect 36100 16836 36156 16892
rect 36156 16836 36160 16892
rect 36096 16832 36160 16836
rect 66576 16892 66640 16896
rect 66576 16836 66580 16892
rect 66580 16836 66636 16892
rect 66636 16836 66640 16892
rect 66576 16832 66640 16836
rect 66656 16892 66720 16896
rect 66656 16836 66660 16892
rect 66660 16836 66716 16892
rect 66716 16836 66720 16892
rect 66656 16832 66720 16836
rect 66736 16892 66800 16896
rect 66736 16836 66740 16892
rect 66740 16836 66796 16892
rect 66796 16836 66800 16892
rect 66736 16832 66800 16836
rect 66816 16892 66880 16896
rect 66816 16836 66820 16892
rect 66820 16836 66876 16892
rect 66876 16836 66880 16892
rect 66816 16832 66880 16836
rect 5796 16348 5860 16352
rect 5796 16292 5800 16348
rect 5800 16292 5856 16348
rect 5856 16292 5860 16348
rect 5796 16288 5860 16292
rect 5876 16348 5940 16352
rect 5876 16292 5880 16348
rect 5880 16292 5936 16348
rect 5936 16292 5940 16348
rect 5876 16288 5940 16292
rect 5956 16348 6020 16352
rect 5956 16292 5960 16348
rect 5960 16292 6016 16348
rect 6016 16292 6020 16348
rect 5956 16288 6020 16292
rect 6036 16348 6100 16352
rect 6036 16292 6040 16348
rect 6040 16292 6096 16348
rect 6096 16292 6100 16348
rect 6036 16288 6100 16292
rect 36516 16348 36580 16352
rect 36516 16292 36520 16348
rect 36520 16292 36576 16348
rect 36576 16292 36580 16348
rect 36516 16288 36580 16292
rect 36596 16348 36660 16352
rect 36596 16292 36600 16348
rect 36600 16292 36656 16348
rect 36656 16292 36660 16348
rect 36596 16288 36660 16292
rect 36676 16348 36740 16352
rect 36676 16292 36680 16348
rect 36680 16292 36736 16348
rect 36736 16292 36740 16348
rect 36676 16288 36740 16292
rect 36756 16348 36820 16352
rect 36756 16292 36760 16348
rect 36760 16292 36816 16348
rect 36816 16292 36820 16348
rect 36756 16288 36820 16292
rect 67236 16348 67300 16352
rect 67236 16292 67240 16348
rect 67240 16292 67296 16348
rect 67296 16292 67300 16348
rect 67236 16288 67300 16292
rect 67316 16348 67380 16352
rect 67316 16292 67320 16348
rect 67320 16292 67376 16348
rect 67376 16292 67380 16348
rect 67316 16288 67380 16292
rect 67396 16348 67460 16352
rect 67396 16292 67400 16348
rect 67400 16292 67456 16348
rect 67456 16292 67460 16348
rect 67396 16288 67460 16292
rect 67476 16348 67540 16352
rect 67476 16292 67480 16348
rect 67480 16292 67536 16348
rect 67536 16292 67540 16348
rect 67476 16288 67540 16292
rect 5136 15804 5200 15808
rect 5136 15748 5140 15804
rect 5140 15748 5196 15804
rect 5196 15748 5200 15804
rect 5136 15744 5200 15748
rect 5216 15804 5280 15808
rect 5216 15748 5220 15804
rect 5220 15748 5276 15804
rect 5276 15748 5280 15804
rect 5216 15744 5280 15748
rect 5296 15804 5360 15808
rect 5296 15748 5300 15804
rect 5300 15748 5356 15804
rect 5356 15748 5360 15804
rect 5296 15744 5360 15748
rect 5376 15804 5440 15808
rect 5376 15748 5380 15804
rect 5380 15748 5436 15804
rect 5436 15748 5440 15804
rect 5376 15744 5440 15748
rect 35856 15804 35920 15808
rect 35856 15748 35860 15804
rect 35860 15748 35916 15804
rect 35916 15748 35920 15804
rect 35856 15744 35920 15748
rect 35936 15804 36000 15808
rect 35936 15748 35940 15804
rect 35940 15748 35996 15804
rect 35996 15748 36000 15804
rect 35936 15744 36000 15748
rect 36016 15804 36080 15808
rect 36016 15748 36020 15804
rect 36020 15748 36076 15804
rect 36076 15748 36080 15804
rect 36016 15744 36080 15748
rect 36096 15804 36160 15808
rect 36096 15748 36100 15804
rect 36100 15748 36156 15804
rect 36156 15748 36160 15804
rect 36096 15744 36160 15748
rect 66576 15804 66640 15808
rect 66576 15748 66580 15804
rect 66580 15748 66636 15804
rect 66636 15748 66640 15804
rect 66576 15744 66640 15748
rect 66656 15804 66720 15808
rect 66656 15748 66660 15804
rect 66660 15748 66716 15804
rect 66716 15748 66720 15804
rect 66656 15744 66720 15748
rect 66736 15804 66800 15808
rect 66736 15748 66740 15804
rect 66740 15748 66796 15804
rect 66796 15748 66800 15804
rect 66736 15744 66800 15748
rect 66816 15804 66880 15808
rect 66816 15748 66820 15804
rect 66820 15748 66876 15804
rect 66876 15748 66880 15804
rect 66816 15744 66880 15748
rect 5796 15260 5860 15264
rect 5796 15204 5800 15260
rect 5800 15204 5856 15260
rect 5856 15204 5860 15260
rect 5796 15200 5860 15204
rect 5876 15260 5940 15264
rect 5876 15204 5880 15260
rect 5880 15204 5936 15260
rect 5936 15204 5940 15260
rect 5876 15200 5940 15204
rect 5956 15260 6020 15264
rect 5956 15204 5960 15260
rect 5960 15204 6016 15260
rect 6016 15204 6020 15260
rect 5956 15200 6020 15204
rect 6036 15260 6100 15264
rect 6036 15204 6040 15260
rect 6040 15204 6096 15260
rect 6096 15204 6100 15260
rect 6036 15200 6100 15204
rect 36516 15260 36580 15264
rect 36516 15204 36520 15260
rect 36520 15204 36576 15260
rect 36576 15204 36580 15260
rect 36516 15200 36580 15204
rect 36596 15260 36660 15264
rect 36596 15204 36600 15260
rect 36600 15204 36656 15260
rect 36656 15204 36660 15260
rect 36596 15200 36660 15204
rect 36676 15260 36740 15264
rect 36676 15204 36680 15260
rect 36680 15204 36736 15260
rect 36736 15204 36740 15260
rect 36676 15200 36740 15204
rect 36756 15260 36820 15264
rect 36756 15204 36760 15260
rect 36760 15204 36816 15260
rect 36816 15204 36820 15260
rect 36756 15200 36820 15204
rect 67236 15260 67300 15264
rect 67236 15204 67240 15260
rect 67240 15204 67296 15260
rect 67296 15204 67300 15260
rect 67236 15200 67300 15204
rect 67316 15260 67380 15264
rect 67316 15204 67320 15260
rect 67320 15204 67376 15260
rect 67376 15204 67380 15260
rect 67316 15200 67380 15204
rect 67396 15260 67460 15264
rect 67396 15204 67400 15260
rect 67400 15204 67456 15260
rect 67456 15204 67460 15260
rect 67396 15200 67460 15204
rect 67476 15260 67540 15264
rect 67476 15204 67480 15260
rect 67480 15204 67536 15260
rect 67536 15204 67540 15260
rect 67476 15200 67540 15204
rect 5136 14716 5200 14720
rect 5136 14660 5140 14716
rect 5140 14660 5196 14716
rect 5196 14660 5200 14716
rect 5136 14656 5200 14660
rect 5216 14716 5280 14720
rect 5216 14660 5220 14716
rect 5220 14660 5276 14716
rect 5276 14660 5280 14716
rect 5216 14656 5280 14660
rect 5296 14716 5360 14720
rect 5296 14660 5300 14716
rect 5300 14660 5356 14716
rect 5356 14660 5360 14716
rect 5296 14656 5360 14660
rect 5376 14716 5440 14720
rect 5376 14660 5380 14716
rect 5380 14660 5436 14716
rect 5436 14660 5440 14716
rect 5376 14656 5440 14660
rect 35856 14716 35920 14720
rect 35856 14660 35860 14716
rect 35860 14660 35916 14716
rect 35916 14660 35920 14716
rect 35856 14656 35920 14660
rect 35936 14716 36000 14720
rect 35936 14660 35940 14716
rect 35940 14660 35996 14716
rect 35996 14660 36000 14716
rect 35936 14656 36000 14660
rect 36016 14716 36080 14720
rect 36016 14660 36020 14716
rect 36020 14660 36076 14716
rect 36076 14660 36080 14716
rect 36016 14656 36080 14660
rect 36096 14716 36160 14720
rect 36096 14660 36100 14716
rect 36100 14660 36156 14716
rect 36156 14660 36160 14716
rect 36096 14656 36160 14660
rect 66576 14716 66640 14720
rect 66576 14660 66580 14716
rect 66580 14660 66636 14716
rect 66636 14660 66640 14716
rect 66576 14656 66640 14660
rect 66656 14716 66720 14720
rect 66656 14660 66660 14716
rect 66660 14660 66716 14716
rect 66716 14660 66720 14716
rect 66656 14656 66720 14660
rect 66736 14716 66800 14720
rect 66736 14660 66740 14716
rect 66740 14660 66796 14716
rect 66796 14660 66800 14716
rect 66736 14656 66800 14660
rect 66816 14716 66880 14720
rect 66816 14660 66820 14716
rect 66820 14660 66876 14716
rect 66876 14660 66880 14716
rect 66816 14656 66880 14660
rect 28580 14452 28644 14516
rect 28212 14316 28276 14380
rect 5796 14172 5860 14176
rect 5796 14116 5800 14172
rect 5800 14116 5856 14172
rect 5856 14116 5860 14172
rect 5796 14112 5860 14116
rect 5876 14172 5940 14176
rect 5876 14116 5880 14172
rect 5880 14116 5936 14172
rect 5936 14116 5940 14172
rect 5876 14112 5940 14116
rect 5956 14172 6020 14176
rect 5956 14116 5960 14172
rect 5960 14116 6016 14172
rect 6016 14116 6020 14172
rect 5956 14112 6020 14116
rect 6036 14172 6100 14176
rect 6036 14116 6040 14172
rect 6040 14116 6096 14172
rect 6096 14116 6100 14172
rect 6036 14112 6100 14116
rect 36516 14172 36580 14176
rect 36516 14116 36520 14172
rect 36520 14116 36576 14172
rect 36576 14116 36580 14172
rect 36516 14112 36580 14116
rect 36596 14172 36660 14176
rect 36596 14116 36600 14172
rect 36600 14116 36656 14172
rect 36656 14116 36660 14172
rect 36596 14112 36660 14116
rect 36676 14172 36740 14176
rect 36676 14116 36680 14172
rect 36680 14116 36736 14172
rect 36736 14116 36740 14172
rect 36676 14112 36740 14116
rect 36756 14172 36820 14176
rect 36756 14116 36760 14172
rect 36760 14116 36816 14172
rect 36816 14116 36820 14172
rect 36756 14112 36820 14116
rect 67236 14172 67300 14176
rect 67236 14116 67240 14172
rect 67240 14116 67296 14172
rect 67296 14116 67300 14172
rect 67236 14112 67300 14116
rect 67316 14172 67380 14176
rect 67316 14116 67320 14172
rect 67320 14116 67376 14172
rect 67376 14116 67380 14172
rect 67316 14112 67380 14116
rect 67396 14172 67460 14176
rect 67396 14116 67400 14172
rect 67400 14116 67456 14172
rect 67456 14116 67460 14172
rect 67396 14112 67460 14116
rect 67476 14172 67540 14176
rect 67476 14116 67480 14172
rect 67480 14116 67536 14172
rect 67536 14116 67540 14172
rect 67476 14112 67540 14116
rect 5136 13628 5200 13632
rect 5136 13572 5140 13628
rect 5140 13572 5196 13628
rect 5196 13572 5200 13628
rect 5136 13568 5200 13572
rect 5216 13628 5280 13632
rect 5216 13572 5220 13628
rect 5220 13572 5276 13628
rect 5276 13572 5280 13628
rect 5216 13568 5280 13572
rect 5296 13628 5360 13632
rect 5296 13572 5300 13628
rect 5300 13572 5356 13628
rect 5356 13572 5360 13628
rect 5296 13568 5360 13572
rect 5376 13628 5440 13632
rect 5376 13572 5380 13628
rect 5380 13572 5436 13628
rect 5436 13572 5440 13628
rect 5376 13568 5440 13572
rect 35856 13628 35920 13632
rect 35856 13572 35860 13628
rect 35860 13572 35916 13628
rect 35916 13572 35920 13628
rect 35856 13568 35920 13572
rect 35936 13628 36000 13632
rect 35936 13572 35940 13628
rect 35940 13572 35996 13628
rect 35996 13572 36000 13628
rect 35936 13568 36000 13572
rect 36016 13628 36080 13632
rect 36016 13572 36020 13628
rect 36020 13572 36076 13628
rect 36076 13572 36080 13628
rect 36016 13568 36080 13572
rect 36096 13628 36160 13632
rect 36096 13572 36100 13628
rect 36100 13572 36156 13628
rect 36156 13572 36160 13628
rect 36096 13568 36160 13572
rect 66576 13628 66640 13632
rect 66576 13572 66580 13628
rect 66580 13572 66636 13628
rect 66636 13572 66640 13628
rect 66576 13568 66640 13572
rect 66656 13628 66720 13632
rect 66656 13572 66660 13628
rect 66660 13572 66716 13628
rect 66716 13572 66720 13628
rect 66656 13568 66720 13572
rect 66736 13628 66800 13632
rect 66736 13572 66740 13628
rect 66740 13572 66796 13628
rect 66796 13572 66800 13628
rect 66736 13568 66800 13572
rect 66816 13628 66880 13632
rect 66816 13572 66820 13628
rect 66820 13572 66876 13628
rect 66876 13572 66880 13628
rect 66816 13568 66880 13572
rect 5796 13084 5860 13088
rect 5796 13028 5800 13084
rect 5800 13028 5856 13084
rect 5856 13028 5860 13084
rect 5796 13024 5860 13028
rect 5876 13084 5940 13088
rect 5876 13028 5880 13084
rect 5880 13028 5936 13084
rect 5936 13028 5940 13084
rect 5876 13024 5940 13028
rect 5956 13084 6020 13088
rect 5956 13028 5960 13084
rect 5960 13028 6016 13084
rect 6016 13028 6020 13084
rect 5956 13024 6020 13028
rect 6036 13084 6100 13088
rect 6036 13028 6040 13084
rect 6040 13028 6096 13084
rect 6096 13028 6100 13084
rect 6036 13024 6100 13028
rect 36516 13084 36580 13088
rect 36516 13028 36520 13084
rect 36520 13028 36576 13084
rect 36576 13028 36580 13084
rect 36516 13024 36580 13028
rect 36596 13084 36660 13088
rect 36596 13028 36600 13084
rect 36600 13028 36656 13084
rect 36656 13028 36660 13084
rect 36596 13024 36660 13028
rect 36676 13084 36740 13088
rect 36676 13028 36680 13084
rect 36680 13028 36736 13084
rect 36736 13028 36740 13084
rect 36676 13024 36740 13028
rect 36756 13084 36820 13088
rect 36756 13028 36760 13084
rect 36760 13028 36816 13084
rect 36816 13028 36820 13084
rect 36756 13024 36820 13028
rect 67236 13084 67300 13088
rect 67236 13028 67240 13084
rect 67240 13028 67296 13084
rect 67296 13028 67300 13084
rect 67236 13024 67300 13028
rect 67316 13084 67380 13088
rect 67316 13028 67320 13084
rect 67320 13028 67376 13084
rect 67376 13028 67380 13084
rect 67316 13024 67380 13028
rect 67396 13084 67460 13088
rect 67396 13028 67400 13084
rect 67400 13028 67456 13084
rect 67456 13028 67460 13084
rect 67396 13024 67460 13028
rect 67476 13084 67540 13088
rect 67476 13028 67480 13084
rect 67480 13028 67536 13084
rect 67536 13028 67540 13084
rect 67476 13024 67540 13028
rect 5136 12540 5200 12544
rect 5136 12484 5140 12540
rect 5140 12484 5196 12540
rect 5196 12484 5200 12540
rect 5136 12480 5200 12484
rect 5216 12540 5280 12544
rect 5216 12484 5220 12540
rect 5220 12484 5276 12540
rect 5276 12484 5280 12540
rect 5216 12480 5280 12484
rect 5296 12540 5360 12544
rect 5296 12484 5300 12540
rect 5300 12484 5356 12540
rect 5356 12484 5360 12540
rect 5296 12480 5360 12484
rect 5376 12540 5440 12544
rect 5376 12484 5380 12540
rect 5380 12484 5436 12540
rect 5436 12484 5440 12540
rect 5376 12480 5440 12484
rect 35856 12540 35920 12544
rect 35856 12484 35860 12540
rect 35860 12484 35916 12540
rect 35916 12484 35920 12540
rect 35856 12480 35920 12484
rect 35936 12540 36000 12544
rect 35936 12484 35940 12540
rect 35940 12484 35996 12540
rect 35996 12484 36000 12540
rect 35936 12480 36000 12484
rect 36016 12540 36080 12544
rect 36016 12484 36020 12540
rect 36020 12484 36076 12540
rect 36076 12484 36080 12540
rect 36016 12480 36080 12484
rect 36096 12540 36160 12544
rect 36096 12484 36100 12540
rect 36100 12484 36156 12540
rect 36156 12484 36160 12540
rect 36096 12480 36160 12484
rect 66576 12540 66640 12544
rect 66576 12484 66580 12540
rect 66580 12484 66636 12540
rect 66636 12484 66640 12540
rect 66576 12480 66640 12484
rect 66656 12540 66720 12544
rect 66656 12484 66660 12540
rect 66660 12484 66716 12540
rect 66716 12484 66720 12540
rect 66656 12480 66720 12484
rect 66736 12540 66800 12544
rect 66736 12484 66740 12540
rect 66740 12484 66796 12540
rect 66796 12484 66800 12540
rect 66736 12480 66800 12484
rect 66816 12540 66880 12544
rect 66816 12484 66820 12540
rect 66820 12484 66876 12540
rect 66876 12484 66880 12540
rect 66816 12480 66880 12484
rect 12756 12412 12820 12476
rect 5796 11996 5860 12000
rect 5796 11940 5800 11996
rect 5800 11940 5856 11996
rect 5856 11940 5860 11996
rect 5796 11936 5860 11940
rect 5876 11996 5940 12000
rect 5876 11940 5880 11996
rect 5880 11940 5936 11996
rect 5936 11940 5940 11996
rect 5876 11936 5940 11940
rect 5956 11996 6020 12000
rect 5956 11940 5960 11996
rect 5960 11940 6016 11996
rect 6016 11940 6020 11996
rect 5956 11936 6020 11940
rect 6036 11996 6100 12000
rect 6036 11940 6040 11996
rect 6040 11940 6096 11996
rect 6096 11940 6100 11996
rect 6036 11936 6100 11940
rect 36516 11996 36580 12000
rect 36516 11940 36520 11996
rect 36520 11940 36576 11996
rect 36576 11940 36580 11996
rect 36516 11936 36580 11940
rect 36596 11996 36660 12000
rect 36596 11940 36600 11996
rect 36600 11940 36656 11996
rect 36656 11940 36660 11996
rect 36596 11936 36660 11940
rect 36676 11996 36740 12000
rect 36676 11940 36680 11996
rect 36680 11940 36736 11996
rect 36736 11940 36740 11996
rect 36676 11936 36740 11940
rect 36756 11996 36820 12000
rect 36756 11940 36760 11996
rect 36760 11940 36816 11996
rect 36816 11940 36820 11996
rect 36756 11936 36820 11940
rect 67236 11996 67300 12000
rect 67236 11940 67240 11996
rect 67240 11940 67296 11996
rect 67296 11940 67300 11996
rect 67236 11936 67300 11940
rect 67316 11996 67380 12000
rect 67316 11940 67320 11996
rect 67320 11940 67376 11996
rect 67376 11940 67380 11996
rect 67316 11936 67380 11940
rect 67396 11996 67460 12000
rect 67396 11940 67400 11996
rect 67400 11940 67456 11996
rect 67456 11940 67460 11996
rect 67396 11936 67460 11940
rect 67476 11996 67540 12000
rect 67476 11940 67480 11996
rect 67480 11940 67536 11996
rect 67536 11940 67540 11996
rect 67476 11936 67540 11940
rect 19932 11460 19996 11524
rect 5136 11452 5200 11456
rect 5136 11396 5140 11452
rect 5140 11396 5196 11452
rect 5196 11396 5200 11452
rect 5136 11392 5200 11396
rect 5216 11452 5280 11456
rect 5216 11396 5220 11452
rect 5220 11396 5276 11452
rect 5276 11396 5280 11452
rect 5216 11392 5280 11396
rect 5296 11452 5360 11456
rect 5296 11396 5300 11452
rect 5300 11396 5356 11452
rect 5356 11396 5360 11452
rect 5296 11392 5360 11396
rect 5376 11452 5440 11456
rect 5376 11396 5380 11452
rect 5380 11396 5436 11452
rect 5436 11396 5440 11452
rect 5376 11392 5440 11396
rect 35856 11452 35920 11456
rect 35856 11396 35860 11452
rect 35860 11396 35916 11452
rect 35916 11396 35920 11452
rect 35856 11392 35920 11396
rect 35936 11452 36000 11456
rect 35936 11396 35940 11452
rect 35940 11396 35996 11452
rect 35996 11396 36000 11452
rect 35936 11392 36000 11396
rect 36016 11452 36080 11456
rect 36016 11396 36020 11452
rect 36020 11396 36076 11452
rect 36076 11396 36080 11452
rect 36016 11392 36080 11396
rect 36096 11452 36160 11456
rect 36096 11396 36100 11452
rect 36100 11396 36156 11452
rect 36156 11396 36160 11452
rect 36096 11392 36160 11396
rect 66576 11452 66640 11456
rect 66576 11396 66580 11452
rect 66580 11396 66636 11452
rect 66636 11396 66640 11452
rect 66576 11392 66640 11396
rect 66656 11452 66720 11456
rect 66656 11396 66660 11452
rect 66660 11396 66716 11452
rect 66716 11396 66720 11452
rect 66656 11392 66720 11396
rect 66736 11452 66800 11456
rect 66736 11396 66740 11452
rect 66740 11396 66796 11452
rect 66796 11396 66800 11452
rect 66736 11392 66800 11396
rect 66816 11452 66880 11456
rect 66816 11396 66820 11452
rect 66820 11396 66876 11452
rect 66876 11396 66880 11452
rect 66816 11392 66880 11396
rect 17724 11324 17788 11388
rect 15332 11188 15396 11252
rect 13308 11052 13372 11116
rect 26556 11052 26620 11116
rect 5796 10908 5860 10912
rect 5796 10852 5800 10908
rect 5800 10852 5856 10908
rect 5856 10852 5860 10908
rect 5796 10848 5860 10852
rect 5876 10908 5940 10912
rect 5876 10852 5880 10908
rect 5880 10852 5936 10908
rect 5936 10852 5940 10908
rect 5876 10848 5940 10852
rect 5956 10908 6020 10912
rect 5956 10852 5960 10908
rect 5960 10852 6016 10908
rect 6016 10852 6020 10908
rect 5956 10848 6020 10852
rect 6036 10908 6100 10912
rect 6036 10852 6040 10908
rect 6040 10852 6096 10908
rect 6096 10852 6100 10908
rect 6036 10848 6100 10852
rect 36516 10908 36580 10912
rect 36516 10852 36520 10908
rect 36520 10852 36576 10908
rect 36576 10852 36580 10908
rect 36516 10848 36580 10852
rect 36596 10908 36660 10912
rect 36596 10852 36600 10908
rect 36600 10852 36656 10908
rect 36656 10852 36660 10908
rect 36596 10848 36660 10852
rect 36676 10908 36740 10912
rect 36676 10852 36680 10908
rect 36680 10852 36736 10908
rect 36736 10852 36740 10908
rect 36676 10848 36740 10852
rect 36756 10908 36820 10912
rect 36756 10852 36760 10908
rect 36760 10852 36816 10908
rect 36816 10852 36820 10908
rect 36756 10848 36820 10852
rect 67236 10908 67300 10912
rect 67236 10852 67240 10908
rect 67240 10852 67296 10908
rect 67296 10852 67300 10908
rect 67236 10848 67300 10852
rect 67316 10908 67380 10912
rect 67316 10852 67320 10908
rect 67320 10852 67376 10908
rect 67376 10852 67380 10908
rect 67316 10848 67380 10852
rect 67396 10908 67460 10912
rect 67396 10852 67400 10908
rect 67400 10852 67456 10908
rect 67456 10852 67460 10908
rect 67396 10848 67460 10852
rect 67476 10908 67540 10912
rect 67476 10852 67480 10908
rect 67480 10852 67536 10908
rect 67536 10852 67540 10908
rect 67476 10848 67540 10852
rect 17356 10780 17420 10844
rect 10732 10644 10796 10708
rect 26188 10568 26252 10572
rect 26188 10512 26238 10568
rect 26238 10512 26252 10568
rect 26188 10508 26252 10512
rect 16436 10372 16500 10436
rect 30972 10372 31036 10436
rect 5136 10364 5200 10368
rect 5136 10308 5140 10364
rect 5140 10308 5196 10364
rect 5196 10308 5200 10364
rect 5136 10304 5200 10308
rect 5216 10364 5280 10368
rect 5216 10308 5220 10364
rect 5220 10308 5276 10364
rect 5276 10308 5280 10364
rect 5216 10304 5280 10308
rect 5296 10364 5360 10368
rect 5296 10308 5300 10364
rect 5300 10308 5356 10364
rect 5356 10308 5360 10364
rect 5296 10304 5360 10308
rect 5376 10364 5440 10368
rect 5376 10308 5380 10364
rect 5380 10308 5436 10364
rect 5436 10308 5440 10364
rect 5376 10304 5440 10308
rect 35856 10364 35920 10368
rect 35856 10308 35860 10364
rect 35860 10308 35916 10364
rect 35916 10308 35920 10364
rect 35856 10304 35920 10308
rect 35936 10364 36000 10368
rect 35936 10308 35940 10364
rect 35940 10308 35996 10364
rect 35996 10308 36000 10364
rect 35936 10304 36000 10308
rect 36016 10364 36080 10368
rect 36016 10308 36020 10364
rect 36020 10308 36076 10364
rect 36076 10308 36080 10364
rect 36016 10304 36080 10308
rect 36096 10364 36160 10368
rect 36096 10308 36100 10364
rect 36100 10308 36156 10364
rect 36156 10308 36160 10364
rect 36096 10304 36160 10308
rect 66576 10364 66640 10368
rect 66576 10308 66580 10364
rect 66580 10308 66636 10364
rect 66636 10308 66640 10364
rect 66576 10304 66640 10308
rect 66656 10364 66720 10368
rect 66656 10308 66660 10364
rect 66660 10308 66716 10364
rect 66716 10308 66720 10364
rect 66656 10304 66720 10308
rect 66736 10364 66800 10368
rect 66736 10308 66740 10364
rect 66740 10308 66796 10364
rect 66796 10308 66800 10364
rect 66736 10304 66800 10308
rect 66816 10364 66880 10368
rect 66816 10308 66820 10364
rect 66820 10308 66876 10364
rect 66876 10308 66880 10364
rect 66816 10304 66880 10308
rect 10916 10236 10980 10300
rect 23060 10236 23124 10300
rect 18092 10100 18156 10164
rect 21772 9964 21836 10028
rect 22692 9964 22756 10028
rect 23796 9964 23860 10028
rect 5796 9820 5860 9824
rect 5796 9764 5800 9820
rect 5800 9764 5856 9820
rect 5856 9764 5860 9820
rect 5796 9760 5860 9764
rect 5876 9820 5940 9824
rect 5876 9764 5880 9820
rect 5880 9764 5936 9820
rect 5936 9764 5940 9820
rect 5876 9760 5940 9764
rect 5956 9820 6020 9824
rect 5956 9764 5960 9820
rect 5960 9764 6016 9820
rect 6016 9764 6020 9820
rect 5956 9760 6020 9764
rect 6036 9820 6100 9824
rect 6036 9764 6040 9820
rect 6040 9764 6096 9820
rect 6096 9764 6100 9820
rect 6036 9760 6100 9764
rect 19748 9556 19812 9620
rect 36516 9820 36580 9824
rect 36516 9764 36520 9820
rect 36520 9764 36576 9820
rect 36576 9764 36580 9820
rect 36516 9760 36580 9764
rect 36596 9820 36660 9824
rect 36596 9764 36600 9820
rect 36600 9764 36656 9820
rect 36656 9764 36660 9820
rect 36596 9760 36660 9764
rect 36676 9820 36740 9824
rect 36676 9764 36680 9820
rect 36680 9764 36736 9820
rect 36736 9764 36740 9820
rect 36676 9760 36740 9764
rect 36756 9820 36820 9824
rect 36756 9764 36760 9820
rect 36760 9764 36816 9820
rect 36816 9764 36820 9820
rect 36756 9760 36820 9764
rect 67236 9820 67300 9824
rect 67236 9764 67240 9820
rect 67240 9764 67296 9820
rect 67296 9764 67300 9820
rect 67236 9760 67300 9764
rect 67316 9820 67380 9824
rect 67316 9764 67320 9820
rect 67320 9764 67376 9820
rect 67376 9764 67380 9820
rect 67316 9760 67380 9764
rect 67396 9820 67460 9824
rect 67396 9764 67400 9820
rect 67400 9764 67456 9820
rect 67456 9764 67460 9820
rect 67396 9760 67460 9764
rect 67476 9820 67540 9824
rect 67476 9764 67480 9820
rect 67480 9764 67536 9820
rect 67536 9764 67540 9820
rect 67476 9760 67540 9764
rect 24900 9692 24964 9756
rect 29132 9692 29196 9756
rect 30236 9752 30300 9756
rect 30236 9696 30250 9752
rect 30250 9696 30300 9752
rect 30236 9692 30300 9696
rect 24164 9284 24228 9348
rect 28948 9616 29012 9620
rect 28948 9560 28998 9616
rect 28998 9560 29012 9616
rect 28948 9556 29012 9560
rect 5136 9276 5200 9280
rect 5136 9220 5140 9276
rect 5140 9220 5196 9276
rect 5196 9220 5200 9276
rect 5136 9216 5200 9220
rect 5216 9276 5280 9280
rect 5216 9220 5220 9276
rect 5220 9220 5276 9276
rect 5276 9220 5280 9276
rect 5216 9216 5280 9220
rect 5296 9276 5360 9280
rect 5296 9220 5300 9276
rect 5300 9220 5356 9276
rect 5356 9220 5360 9276
rect 5296 9216 5360 9220
rect 5376 9276 5440 9280
rect 5376 9220 5380 9276
rect 5380 9220 5436 9276
rect 5436 9220 5440 9276
rect 5376 9216 5440 9220
rect 35856 9276 35920 9280
rect 35856 9220 35860 9276
rect 35860 9220 35916 9276
rect 35916 9220 35920 9276
rect 35856 9216 35920 9220
rect 35936 9276 36000 9280
rect 35936 9220 35940 9276
rect 35940 9220 35996 9276
rect 35996 9220 36000 9276
rect 35936 9216 36000 9220
rect 36016 9276 36080 9280
rect 36016 9220 36020 9276
rect 36020 9220 36076 9276
rect 36076 9220 36080 9276
rect 36016 9216 36080 9220
rect 36096 9276 36160 9280
rect 36096 9220 36100 9276
rect 36100 9220 36156 9276
rect 36156 9220 36160 9276
rect 36096 9216 36160 9220
rect 66576 9276 66640 9280
rect 66576 9220 66580 9276
rect 66580 9220 66636 9276
rect 66636 9220 66640 9276
rect 66576 9216 66640 9220
rect 66656 9276 66720 9280
rect 66656 9220 66660 9276
rect 66660 9220 66716 9276
rect 66716 9220 66720 9276
rect 66656 9216 66720 9220
rect 66736 9276 66800 9280
rect 66736 9220 66740 9276
rect 66740 9220 66796 9276
rect 66796 9220 66800 9276
rect 66736 9216 66800 9220
rect 66816 9276 66880 9280
rect 66816 9220 66820 9276
rect 66820 9220 66876 9276
rect 66876 9220 66880 9276
rect 66816 9216 66880 9220
rect 24716 9012 24780 9076
rect 29316 9012 29380 9076
rect 28764 8876 28828 8940
rect 17908 8740 17972 8804
rect 18644 8740 18708 8804
rect 5796 8732 5860 8736
rect 5796 8676 5800 8732
rect 5800 8676 5856 8732
rect 5856 8676 5860 8732
rect 5796 8672 5860 8676
rect 5876 8732 5940 8736
rect 5876 8676 5880 8732
rect 5880 8676 5936 8732
rect 5936 8676 5940 8732
rect 5876 8672 5940 8676
rect 5956 8732 6020 8736
rect 5956 8676 5960 8732
rect 5960 8676 6016 8732
rect 6016 8676 6020 8732
rect 5956 8672 6020 8676
rect 6036 8732 6100 8736
rect 6036 8676 6040 8732
rect 6040 8676 6096 8732
rect 6096 8676 6100 8732
rect 6036 8672 6100 8676
rect 36516 8732 36580 8736
rect 36516 8676 36520 8732
rect 36520 8676 36576 8732
rect 36576 8676 36580 8732
rect 36516 8672 36580 8676
rect 36596 8732 36660 8736
rect 36596 8676 36600 8732
rect 36600 8676 36656 8732
rect 36656 8676 36660 8732
rect 36596 8672 36660 8676
rect 36676 8732 36740 8736
rect 36676 8676 36680 8732
rect 36680 8676 36736 8732
rect 36736 8676 36740 8732
rect 36676 8672 36740 8676
rect 36756 8732 36820 8736
rect 36756 8676 36760 8732
rect 36760 8676 36816 8732
rect 36816 8676 36820 8732
rect 36756 8672 36820 8676
rect 67236 8732 67300 8736
rect 67236 8676 67240 8732
rect 67240 8676 67296 8732
rect 67296 8676 67300 8732
rect 67236 8672 67300 8676
rect 67316 8732 67380 8736
rect 67316 8676 67320 8732
rect 67320 8676 67376 8732
rect 67376 8676 67380 8732
rect 67316 8672 67380 8676
rect 67396 8732 67460 8736
rect 67396 8676 67400 8732
rect 67400 8676 67456 8732
rect 67456 8676 67460 8732
rect 67396 8672 67460 8676
rect 67476 8732 67540 8736
rect 67476 8676 67480 8732
rect 67480 8676 67536 8732
rect 67536 8676 67540 8732
rect 67476 8672 67540 8676
rect 18276 8468 18340 8532
rect 19380 8468 19444 8532
rect 18460 8332 18524 8396
rect 25268 8468 25332 8532
rect 31156 8468 31220 8532
rect 33364 8468 33428 8532
rect 37044 8468 37108 8532
rect 20668 8332 20732 8396
rect 25820 8332 25884 8396
rect 27476 8332 27540 8396
rect 31892 8332 31956 8396
rect 33180 8332 33244 8396
rect 33732 8332 33796 8396
rect 5136 8188 5200 8192
rect 5136 8132 5140 8188
rect 5140 8132 5196 8188
rect 5196 8132 5200 8188
rect 5136 8128 5200 8132
rect 5216 8188 5280 8192
rect 5216 8132 5220 8188
rect 5220 8132 5276 8188
rect 5276 8132 5280 8188
rect 5216 8128 5280 8132
rect 5296 8188 5360 8192
rect 5296 8132 5300 8188
rect 5300 8132 5356 8188
rect 5356 8132 5360 8188
rect 5296 8128 5360 8132
rect 5376 8188 5440 8192
rect 5376 8132 5380 8188
rect 5380 8132 5436 8188
rect 5436 8132 5440 8188
rect 5376 8128 5440 8132
rect 35856 8188 35920 8192
rect 35856 8132 35860 8188
rect 35860 8132 35916 8188
rect 35916 8132 35920 8188
rect 35856 8128 35920 8132
rect 35936 8188 36000 8192
rect 35936 8132 35940 8188
rect 35940 8132 35996 8188
rect 35996 8132 36000 8188
rect 35936 8128 36000 8132
rect 36016 8188 36080 8192
rect 36016 8132 36020 8188
rect 36020 8132 36076 8188
rect 36076 8132 36080 8188
rect 36016 8128 36080 8132
rect 36096 8188 36160 8192
rect 36096 8132 36100 8188
rect 36100 8132 36156 8188
rect 36156 8132 36160 8188
rect 36096 8128 36160 8132
rect 66576 8188 66640 8192
rect 66576 8132 66580 8188
rect 66580 8132 66636 8188
rect 66636 8132 66640 8188
rect 66576 8128 66640 8132
rect 66656 8188 66720 8192
rect 66656 8132 66660 8188
rect 66660 8132 66716 8188
rect 66716 8132 66720 8188
rect 66656 8128 66720 8132
rect 66736 8188 66800 8192
rect 66736 8132 66740 8188
rect 66740 8132 66796 8188
rect 66796 8132 66800 8188
rect 66736 8128 66800 8132
rect 66816 8188 66880 8192
rect 66816 8132 66820 8188
rect 66820 8132 66876 8188
rect 66876 8132 66880 8188
rect 66816 8128 66880 8132
rect 17172 8060 17236 8124
rect 24900 7924 24964 7988
rect 28212 7924 28276 7988
rect 33548 7924 33612 7988
rect 20116 7788 20180 7852
rect 30604 7848 30668 7852
rect 30604 7792 30654 7848
rect 30654 7792 30668 7848
rect 30604 7788 30668 7792
rect 32260 7848 32324 7852
rect 32260 7792 32310 7848
rect 32310 7792 32324 7848
rect 32260 7788 32324 7792
rect 13676 7652 13740 7716
rect 27108 7652 27172 7716
rect 34468 7652 34532 7716
rect 5796 7644 5860 7648
rect 5796 7588 5800 7644
rect 5800 7588 5856 7644
rect 5856 7588 5860 7644
rect 5796 7584 5860 7588
rect 5876 7644 5940 7648
rect 5876 7588 5880 7644
rect 5880 7588 5936 7644
rect 5936 7588 5940 7644
rect 5876 7584 5940 7588
rect 5956 7644 6020 7648
rect 5956 7588 5960 7644
rect 5960 7588 6016 7644
rect 6016 7588 6020 7644
rect 5956 7584 6020 7588
rect 6036 7644 6100 7648
rect 6036 7588 6040 7644
rect 6040 7588 6096 7644
rect 6096 7588 6100 7644
rect 6036 7584 6100 7588
rect 36516 7644 36580 7648
rect 36516 7588 36520 7644
rect 36520 7588 36576 7644
rect 36576 7588 36580 7644
rect 36516 7584 36580 7588
rect 36596 7644 36660 7648
rect 36596 7588 36600 7644
rect 36600 7588 36656 7644
rect 36656 7588 36660 7644
rect 36596 7584 36660 7588
rect 36676 7644 36740 7648
rect 36676 7588 36680 7644
rect 36680 7588 36736 7644
rect 36736 7588 36740 7644
rect 36676 7584 36740 7588
rect 36756 7644 36820 7648
rect 36756 7588 36760 7644
rect 36760 7588 36816 7644
rect 36816 7588 36820 7644
rect 36756 7584 36820 7588
rect 67236 7644 67300 7648
rect 67236 7588 67240 7644
rect 67240 7588 67296 7644
rect 67296 7588 67300 7644
rect 67236 7584 67300 7588
rect 67316 7644 67380 7648
rect 67316 7588 67320 7644
rect 67320 7588 67376 7644
rect 67376 7588 67380 7644
rect 67316 7584 67380 7588
rect 67396 7644 67460 7648
rect 67396 7588 67400 7644
rect 67400 7588 67456 7644
rect 67456 7588 67460 7644
rect 67396 7584 67460 7588
rect 67476 7644 67540 7648
rect 67476 7588 67480 7644
rect 67480 7588 67536 7644
rect 67536 7588 67540 7644
rect 67476 7584 67540 7588
rect 27292 7516 27356 7580
rect 23428 7380 23492 7444
rect 21220 7244 21284 7308
rect 32812 7244 32876 7308
rect 27292 7108 27356 7172
rect 5136 7100 5200 7104
rect 5136 7044 5140 7100
rect 5140 7044 5196 7100
rect 5196 7044 5200 7100
rect 5136 7040 5200 7044
rect 5216 7100 5280 7104
rect 5216 7044 5220 7100
rect 5220 7044 5276 7100
rect 5276 7044 5280 7100
rect 5216 7040 5280 7044
rect 5296 7100 5360 7104
rect 5296 7044 5300 7100
rect 5300 7044 5356 7100
rect 5356 7044 5360 7100
rect 5296 7040 5360 7044
rect 5376 7100 5440 7104
rect 5376 7044 5380 7100
rect 5380 7044 5436 7100
rect 5436 7044 5440 7100
rect 5376 7040 5440 7044
rect 5796 6556 5860 6560
rect 5796 6500 5800 6556
rect 5800 6500 5856 6556
rect 5856 6500 5860 6556
rect 5796 6496 5860 6500
rect 5876 6556 5940 6560
rect 5876 6500 5880 6556
rect 5880 6500 5936 6556
rect 5936 6500 5940 6556
rect 5876 6496 5940 6500
rect 5956 6556 6020 6560
rect 5956 6500 5960 6556
rect 5960 6500 6016 6556
rect 6016 6500 6020 6556
rect 5956 6496 6020 6500
rect 6036 6556 6100 6560
rect 6036 6500 6040 6556
rect 6040 6500 6096 6556
rect 6096 6500 6100 6556
rect 6036 6496 6100 6500
rect 35856 7100 35920 7104
rect 35856 7044 35860 7100
rect 35860 7044 35916 7100
rect 35916 7044 35920 7100
rect 35856 7040 35920 7044
rect 35936 7100 36000 7104
rect 35936 7044 35940 7100
rect 35940 7044 35996 7100
rect 35996 7044 36000 7100
rect 35936 7040 36000 7044
rect 36016 7100 36080 7104
rect 36016 7044 36020 7100
rect 36020 7044 36076 7100
rect 36076 7044 36080 7100
rect 36016 7040 36080 7044
rect 36096 7100 36160 7104
rect 36096 7044 36100 7100
rect 36100 7044 36156 7100
rect 36156 7044 36160 7100
rect 36096 7040 36160 7044
rect 66576 7100 66640 7104
rect 66576 7044 66580 7100
rect 66580 7044 66636 7100
rect 66636 7044 66640 7100
rect 66576 7040 66640 7044
rect 66656 7100 66720 7104
rect 66656 7044 66660 7100
rect 66660 7044 66716 7100
rect 66716 7044 66720 7100
rect 66656 7040 66720 7044
rect 66736 7100 66800 7104
rect 66736 7044 66740 7100
rect 66740 7044 66796 7100
rect 66796 7044 66800 7100
rect 66736 7040 66800 7044
rect 66816 7100 66880 7104
rect 66816 7044 66820 7100
rect 66820 7044 66876 7100
rect 66876 7044 66880 7100
rect 66816 7040 66880 7044
rect 30972 6836 31036 6900
rect 35020 6836 35084 6900
rect 36516 6556 36580 6560
rect 36516 6500 36520 6556
rect 36520 6500 36576 6556
rect 36576 6500 36580 6556
rect 36516 6496 36580 6500
rect 36596 6556 36660 6560
rect 36596 6500 36600 6556
rect 36600 6500 36656 6556
rect 36656 6500 36660 6556
rect 36596 6496 36660 6500
rect 36676 6556 36740 6560
rect 36676 6500 36680 6556
rect 36680 6500 36736 6556
rect 36736 6500 36740 6556
rect 36676 6496 36740 6500
rect 36756 6556 36820 6560
rect 36756 6500 36760 6556
rect 36760 6500 36816 6556
rect 36816 6500 36820 6556
rect 36756 6496 36820 6500
rect 22140 6428 22204 6492
rect 17172 6156 17236 6220
rect 67236 6556 67300 6560
rect 67236 6500 67240 6556
rect 67240 6500 67296 6556
rect 67296 6500 67300 6556
rect 67236 6496 67300 6500
rect 67316 6556 67380 6560
rect 67316 6500 67320 6556
rect 67320 6500 67376 6556
rect 67376 6500 67380 6556
rect 67316 6496 67380 6500
rect 67396 6556 67460 6560
rect 67396 6500 67400 6556
rect 67400 6500 67456 6556
rect 67456 6500 67460 6556
rect 67396 6496 67460 6500
rect 67476 6556 67540 6560
rect 67476 6500 67480 6556
rect 67480 6500 67536 6556
rect 67536 6500 67540 6556
rect 67476 6496 67540 6500
rect 16068 6020 16132 6084
rect 16436 6080 16500 6084
rect 16436 6024 16450 6080
rect 16450 6024 16500 6080
rect 16436 6020 16500 6024
rect 16988 6020 17052 6084
rect 18092 6020 18156 6084
rect 18644 6080 18708 6084
rect 18644 6024 18658 6080
rect 18658 6024 18708 6080
rect 18644 6020 18708 6024
rect 28580 6020 28644 6084
rect 5136 6012 5200 6016
rect 5136 5956 5140 6012
rect 5140 5956 5196 6012
rect 5196 5956 5200 6012
rect 5136 5952 5200 5956
rect 5216 6012 5280 6016
rect 5216 5956 5220 6012
rect 5220 5956 5276 6012
rect 5276 5956 5280 6012
rect 5216 5952 5280 5956
rect 5296 6012 5360 6016
rect 5296 5956 5300 6012
rect 5300 5956 5356 6012
rect 5356 5956 5360 6012
rect 5296 5952 5360 5956
rect 5376 6012 5440 6016
rect 5376 5956 5380 6012
rect 5380 5956 5436 6012
rect 5436 5956 5440 6012
rect 5376 5952 5440 5956
rect 20668 5884 20732 5948
rect 23796 5944 23860 5948
rect 23796 5888 23810 5944
rect 23810 5888 23860 5944
rect 23796 5884 23860 5888
rect 28396 5884 28460 5948
rect 35856 6012 35920 6016
rect 35856 5956 35860 6012
rect 35860 5956 35916 6012
rect 35916 5956 35920 6012
rect 35856 5952 35920 5956
rect 35936 6012 36000 6016
rect 35936 5956 35940 6012
rect 35940 5956 35996 6012
rect 35996 5956 36000 6012
rect 35936 5952 36000 5956
rect 36016 6012 36080 6016
rect 36016 5956 36020 6012
rect 36020 5956 36076 6012
rect 36076 5956 36080 6012
rect 36016 5952 36080 5956
rect 36096 6012 36160 6016
rect 36096 5956 36100 6012
rect 36100 5956 36156 6012
rect 36156 5956 36160 6012
rect 36096 5952 36160 5956
rect 66576 6012 66640 6016
rect 66576 5956 66580 6012
rect 66580 5956 66636 6012
rect 66636 5956 66640 6012
rect 66576 5952 66640 5956
rect 66656 6012 66720 6016
rect 66656 5956 66660 6012
rect 66660 5956 66716 6012
rect 66716 5956 66720 6012
rect 66656 5952 66720 5956
rect 66736 6012 66800 6016
rect 66736 5956 66740 6012
rect 66740 5956 66796 6012
rect 66796 5956 66800 6012
rect 66736 5952 66800 5956
rect 66816 6012 66880 6016
rect 66816 5956 66820 6012
rect 66820 5956 66876 6012
rect 66876 5956 66880 6012
rect 66816 5952 66880 5956
rect 19196 5748 19260 5812
rect 19932 5748 19996 5812
rect 21220 5748 21284 5812
rect 22692 5612 22756 5676
rect 24164 5476 24228 5540
rect 27476 5476 27540 5540
rect 5796 5468 5860 5472
rect 5796 5412 5800 5468
rect 5800 5412 5856 5468
rect 5856 5412 5860 5468
rect 5796 5408 5860 5412
rect 5876 5468 5940 5472
rect 5876 5412 5880 5468
rect 5880 5412 5936 5468
rect 5936 5412 5940 5468
rect 5876 5408 5940 5412
rect 5956 5468 6020 5472
rect 5956 5412 5960 5468
rect 5960 5412 6016 5468
rect 6016 5412 6020 5468
rect 5956 5408 6020 5412
rect 6036 5468 6100 5472
rect 6036 5412 6040 5468
rect 6040 5412 6096 5468
rect 6096 5412 6100 5468
rect 6036 5408 6100 5412
rect 36516 5468 36580 5472
rect 36516 5412 36520 5468
rect 36520 5412 36576 5468
rect 36576 5412 36580 5468
rect 36516 5408 36580 5412
rect 36596 5468 36660 5472
rect 36596 5412 36600 5468
rect 36600 5412 36656 5468
rect 36656 5412 36660 5468
rect 36596 5408 36660 5412
rect 36676 5468 36740 5472
rect 36676 5412 36680 5468
rect 36680 5412 36736 5468
rect 36736 5412 36740 5468
rect 36676 5408 36740 5412
rect 36756 5468 36820 5472
rect 36756 5412 36760 5468
rect 36760 5412 36816 5468
rect 36816 5412 36820 5468
rect 36756 5408 36820 5412
rect 67236 5468 67300 5472
rect 67236 5412 67240 5468
rect 67240 5412 67296 5468
rect 67296 5412 67300 5468
rect 67236 5408 67300 5412
rect 67316 5468 67380 5472
rect 67316 5412 67320 5468
rect 67320 5412 67376 5468
rect 67376 5412 67380 5468
rect 67316 5408 67380 5412
rect 67396 5468 67460 5472
rect 67396 5412 67400 5468
rect 67400 5412 67456 5468
rect 67456 5412 67460 5468
rect 67396 5408 67460 5412
rect 67476 5468 67540 5472
rect 67476 5412 67480 5468
rect 67480 5412 67536 5468
rect 67536 5412 67540 5468
rect 67476 5408 67540 5412
rect 15332 5340 15396 5404
rect 13308 5204 13372 5268
rect 29132 5340 29196 5404
rect 22140 5204 22204 5268
rect 32260 5264 32324 5268
rect 32260 5208 32274 5264
rect 32274 5208 32324 5264
rect 32260 5204 32324 5208
rect 28948 4992 29012 4996
rect 28948 4936 28998 4992
rect 28998 4936 29012 4992
rect 28948 4932 29012 4936
rect 5136 4924 5200 4928
rect 5136 4868 5140 4924
rect 5140 4868 5196 4924
rect 5196 4868 5200 4924
rect 5136 4864 5200 4868
rect 5216 4924 5280 4928
rect 5216 4868 5220 4924
rect 5220 4868 5276 4924
rect 5276 4868 5280 4924
rect 5216 4864 5280 4868
rect 5296 4924 5360 4928
rect 5296 4868 5300 4924
rect 5300 4868 5356 4924
rect 5356 4868 5360 4924
rect 5296 4864 5360 4868
rect 5376 4924 5440 4928
rect 5376 4868 5380 4924
rect 5380 4868 5436 4924
rect 5436 4868 5440 4924
rect 5376 4864 5440 4868
rect 35856 4924 35920 4928
rect 35856 4868 35860 4924
rect 35860 4868 35916 4924
rect 35916 4868 35920 4924
rect 35856 4864 35920 4868
rect 35936 4924 36000 4928
rect 35936 4868 35940 4924
rect 35940 4868 35996 4924
rect 35996 4868 36000 4924
rect 35936 4864 36000 4868
rect 36016 4924 36080 4928
rect 36016 4868 36020 4924
rect 36020 4868 36076 4924
rect 36076 4868 36080 4924
rect 36016 4864 36080 4868
rect 36096 4924 36160 4928
rect 36096 4868 36100 4924
rect 36100 4868 36156 4924
rect 36156 4868 36160 4924
rect 36096 4864 36160 4868
rect 66576 4924 66640 4928
rect 66576 4868 66580 4924
rect 66580 4868 66636 4924
rect 66636 4868 66640 4924
rect 66576 4864 66640 4868
rect 66656 4924 66720 4928
rect 66656 4868 66660 4924
rect 66660 4868 66716 4924
rect 66716 4868 66720 4924
rect 66656 4864 66720 4868
rect 66736 4924 66800 4928
rect 66736 4868 66740 4924
rect 66740 4868 66796 4924
rect 66796 4868 66800 4924
rect 66736 4864 66800 4868
rect 66816 4924 66880 4928
rect 66816 4868 66820 4924
rect 66820 4868 66876 4924
rect 66876 4868 66880 4924
rect 66816 4864 66880 4868
rect 12756 4796 12820 4860
rect 17356 4796 17420 4860
rect 17724 4856 17788 4860
rect 17724 4800 17738 4856
rect 17738 4800 17788 4856
rect 17724 4796 17788 4800
rect 19748 4796 19812 4860
rect 28764 4796 28828 4860
rect 15148 4388 15212 4452
rect 20116 4388 20180 4452
rect 5796 4380 5860 4384
rect 5796 4324 5800 4380
rect 5800 4324 5856 4380
rect 5856 4324 5860 4380
rect 5796 4320 5860 4324
rect 5876 4380 5940 4384
rect 5876 4324 5880 4380
rect 5880 4324 5936 4380
rect 5936 4324 5940 4380
rect 5876 4320 5940 4324
rect 5956 4380 6020 4384
rect 5956 4324 5960 4380
rect 5960 4324 6016 4380
rect 6016 4324 6020 4380
rect 5956 4320 6020 4324
rect 6036 4380 6100 4384
rect 6036 4324 6040 4380
rect 6040 4324 6096 4380
rect 6096 4324 6100 4380
rect 6036 4320 6100 4324
rect 36516 4380 36580 4384
rect 36516 4324 36520 4380
rect 36520 4324 36576 4380
rect 36576 4324 36580 4380
rect 36516 4320 36580 4324
rect 36596 4380 36660 4384
rect 36596 4324 36600 4380
rect 36600 4324 36656 4380
rect 36656 4324 36660 4380
rect 36596 4320 36660 4324
rect 36676 4380 36740 4384
rect 36676 4324 36680 4380
rect 36680 4324 36736 4380
rect 36736 4324 36740 4380
rect 36676 4320 36740 4324
rect 36756 4380 36820 4384
rect 36756 4324 36760 4380
rect 36760 4324 36816 4380
rect 36816 4324 36820 4380
rect 36756 4320 36820 4324
rect 67236 4380 67300 4384
rect 67236 4324 67240 4380
rect 67240 4324 67296 4380
rect 67296 4324 67300 4380
rect 67236 4320 67300 4324
rect 67316 4380 67380 4384
rect 67316 4324 67320 4380
rect 67320 4324 67376 4380
rect 67376 4324 67380 4380
rect 67316 4320 67380 4324
rect 67396 4380 67460 4384
rect 67396 4324 67400 4380
rect 67400 4324 67456 4380
rect 67456 4324 67460 4380
rect 67396 4320 67460 4324
rect 67476 4380 67540 4384
rect 67476 4324 67480 4380
rect 67480 4324 67536 4380
rect 67536 4324 67540 4380
rect 67476 4320 67540 4324
rect 24716 4116 24780 4180
rect 29316 4116 29380 4180
rect 10916 4040 10980 4044
rect 10916 3984 10930 4040
rect 10930 3984 10980 4040
rect 10916 3980 10980 3984
rect 21772 3980 21836 4044
rect 23060 3980 23124 4044
rect 25820 3980 25884 4044
rect 26556 3980 26620 4044
rect 11836 3844 11900 3908
rect 13676 3844 13740 3908
rect 16988 3904 17052 3908
rect 16988 3848 17002 3904
rect 17002 3848 17052 3904
rect 16988 3844 17052 3848
rect 5136 3836 5200 3840
rect 5136 3780 5140 3836
rect 5140 3780 5196 3836
rect 5196 3780 5200 3836
rect 5136 3776 5200 3780
rect 5216 3836 5280 3840
rect 5216 3780 5220 3836
rect 5220 3780 5276 3836
rect 5276 3780 5280 3836
rect 5216 3776 5280 3780
rect 5296 3836 5360 3840
rect 5296 3780 5300 3836
rect 5300 3780 5356 3836
rect 5356 3780 5360 3836
rect 5296 3776 5360 3780
rect 5376 3836 5440 3840
rect 5376 3780 5380 3836
rect 5380 3780 5436 3836
rect 5436 3780 5440 3836
rect 5376 3776 5440 3780
rect 35856 3836 35920 3840
rect 35856 3780 35860 3836
rect 35860 3780 35916 3836
rect 35916 3780 35920 3836
rect 35856 3776 35920 3780
rect 35936 3836 36000 3840
rect 35936 3780 35940 3836
rect 35940 3780 35996 3836
rect 35996 3780 36000 3836
rect 35936 3776 36000 3780
rect 36016 3836 36080 3840
rect 36016 3780 36020 3836
rect 36020 3780 36076 3836
rect 36076 3780 36080 3836
rect 36016 3776 36080 3780
rect 36096 3836 36160 3840
rect 36096 3780 36100 3836
rect 36100 3780 36156 3836
rect 36156 3780 36160 3836
rect 36096 3776 36160 3780
rect 66576 3836 66640 3840
rect 66576 3780 66580 3836
rect 66580 3780 66636 3836
rect 66636 3780 66640 3836
rect 66576 3776 66640 3780
rect 66656 3836 66720 3840
rect 66656 3780 66660 3836
rect 66660 3780 66716 3836
rect 66716 3780 66720 3836
rect 66656 3776 66720 3780
rect 66736 3836 66800 3840
rect 66736 3780 66740 3836
rect 66740 3780 66796 3836
rect 66796 3780 66800 3836
rect 66736 3776 66800 3780
rect 66816 3836 66880 3840
rect 66816 3780 66820 3836
rect 66820 3780 66876 3836
rect 66876 3780 66880 3836
rect 66816 3776 66880 3780
rect 4844 3572 4908 3636
rect 74028 3768 74092 3772
rect 74028 3712 74078 3768
rect 74078 3712 74092 3768
rect 74028 3708 74092 3712
rect 28580 3572 28644 3636
rect 16068 3300 16132 3364
rect 31892 3300 31956 3364
rect 5796 3292 5860 3296
rect 5796 3236 5800 3292
rect 5800 3236 5856 3292
rect 5856 3236 5860 3292
rect 5796 3232 5860 3236
rect 5876 3292 5940 3296
rect 5876 3236 5880 3292
rect 5880 3236 5936 3292
rect 5936 3236 5940 3292
rect 5876 3232 5940 3236
rect 5956 3292 6020 3296
rect 5956 3236 5960 3292
rect 5960 3236 6016 3292
rect 6016 3236 6020 3292
rect 5956 3232 6020 3236
rect 6036 3292 6100 3296
rect 6036 3236 6040 3292
rect 6040 3236 6096 3292
rect 6096 3236 6100 3292
rect 6036 3232 6100 3236
rect 36516 3292 36580 3296
rect 36516 3236 36520 3292
rect 36520 3236 36576 3292
rect 36576 3236 36580 3292
rect 36516 3232 36580 3236
rect 36596 3292 36660 3296
rect 36596 3236 36600 3292
rect 36600 3236 36656 3292
rect 36656 3236 36660 3292
rect 36596 3232 36660 3236
rect 36676 3292 36740 3296
rect 36676 3236 36680 3292
rect 36680 3236 36736 3292
rect 36736 3236 36740 3292
rect 36676 3232 36740 3236
rect 36756 3292 36820 3296
rect 36756 3236 36760 3292
rect 36760 3236 36816 3292
rect 36816 3236 36820 3292
rect 36756 3232 36820 3236
rect 67236 3292 67300 3296
rect 67236 3236 67240 3292
rect 67240 3236 67296 3292
rect 67296 3236 67300 3292
rect 67236 3232 67300 3236
rect 67316 3292 67380 3296
rect 67316 3236 67320 3292
rect 67320 3236 67376 3292
rect 67376 3236 67380 3292
rect 67316 3232 67380 3236
rect 67396 3292 67460 3296
rect 67396 3236 67400 3292
rect 67400 3236 67456 3292
rect 67456 3236 67460 3292
rect 67396 3232 67460 3236
rect 67476 3292 67540 3296
rect 67476 3236 67480 3292
rect 67480 3236 67536 3292
rect 67536 3236 67540 3292
rect 67476 3232 67540 3236
rect 23428 3164 23492 3228
rect 25268 3164 25332 3228
rect 27292 3088 27356 3092
rect 27292 3032 27342 3088
rect 27342 3032 27356 3088
rect 27292 3028 27356 3032
rect 37044 2892 37108 2956
rect 31156 2756 31220 2820
rect 5136 2748 5200 2752
rect 5136 2692 5140 2748
rect 5140 2692 5196 2748
rect 5196 2692 5200 2748
rect 5136 2688 5200 2692
rect 5216 2748 5280 2752
rect 5216 2692 5220 2748
rect 5220 2692 5276 2748
rect 5276 2692 5280 2748
rect 5216 2688 5280 2692
rect 5296 2748 5360 2752
rect 5296 2692 5300 2748
rect 5300 2692 5356 2748
rect 5356 2692 5360 2748
rect 5296 2688 5360 2692
rect 5376 2748 5440 2752
rect 5376 2692 5380 2748
rect 5380 2692 5436 2748
rect 5436 2692 5440 2748
rect 5376 2688 5440 2692
rect 35856 2748 35920 2752
rect 35856 2692 35860 2748
rect 35860 2692 35916 2748
rect 35916 2692 35920 2748
rect 35856 2688 35920 2692
rect 35936 2748 36000 2752
rect 35936 2692 35940 2748
rect 35940 2692 35996 2748
rect 35996 2692 36000 2748
rect 35936 2688 36000 2692
rect 36016 2748 36080 2752
rect 36016 2692 36020 2748
rect 36020 2692 36076 2748
rect 36076 2692 36080 2748
rect 36016 2688 36080 2692
rect 36096 2748 36160 2752
rect 36096 2692 36100 2748
rect 36100 2692 36156 2748
rect 36156 2692 36160 2748
rect 36096 2688 36160 2692
rect 66576 2748 66640 2752
rect 66576 2692 66580 2748
rect 66580 2692 66636 2748
rect 66636 2692 66640 2748
rect 66576 2688 66640 2692
rect 66656 2748 66720 2752
rect 66656 2692 66660 2748
rect 66660 2692 66716 2748
rect 66716 2692 66720 2748
rect 66656 2688 66720 2692
rect 66736 2748 66800 2752
rect 66736 2692 66740 2748
rect 66740 2692 66796 2748
rect 66796 2692 66800 2748
rect 66736 2688 66800 2692
rect 66816 2748 66880 2752
rect 66816 2692 66820 2748
rect 66820 2692 66876 2748
rect 66876 2692 66880 2748
rect 66816 2688 66880 2692
rect 10732 2620 10796 2684
rect 18276 2620 18340 2684
rect 33548 2620 33612 2684
rect 17908 2484 17972 2548
rect 33364 2484 33428 2548
rect 18460 2348 18524 2412
rect 24716 2348 24780 2412
rect 5796 2204 5860 2208
rect 5796 2148 5800 2204
rect 5800 2148 5856 2204
rect 5856 2148 5860 2204
rect 5796 2144 5860 2148
rect 5876 2204 5940 2208
rect 5876 2148 5880 2204
rect 5880 2148 5936 2204
rect 5936 2148 5940 2204
rect 5876 2144 5940 2148
rect 5956 2204 6020 2208
rect 5956 2148 5960 2204
rect 5960 2148 6016 2204
rect 6016 2148 6020 2204
rect 5956 2144 6020 2148
rect 6036 2204 6100 2208
rect 6036 2148 6040 2204
rect 6040 2148 6096 2204
rect 6096 2148 6100 2204
rect 6036 2144 6100 2148
rect 34468 2212 34532 2276
rect 36516 2204 36580 2208
rect 36516 2148 36520 2204
rect 36520 2148 36576 2204
rect 36576 2148 36580 2204
rect 36516 2144 36580 2148
rect 36596 2204 36660 2208
rect 36596 2148 36600 2204
rect 36600 2148 36656 2204
rect 36656 2148 36660 2204
rect 36596 2144 36660 2148
rect 36676 2204 36740 2208
rect 36676 2148 36680 2204
rect 36680 2148 36736 2204
rect 36736 2148 36740 2204
rect 36676 2144 36740 2148
rect 36756 2204 36820 2208
rect 36756 2148 36760 2204
rect 36760 2148 36816 2204
rect 36816 2148 36820 2204
rect 36756 2144 36820 2148
rect 67236 2204 67300 2208
rect 67236 2148 67240 2204
rect 67240 2148 67296 2204
rect 67296 2148 67300 2204
rect 67236 2144 67300 2148
rect 67316 2204 67380 2208
rect 67316 2148 67320 2204
rect 67320 2148 67376 2204
rect 67376 2148 67380 2204
rect 67316 2144 67380 2148
rect 67396 2204 67460 2208
rect 67396 2148 67400 2204
rect 67400 2148 67456 2204
rect 67456 2148 67460 2204
rect 67396 2144 67460 2148
rect 67476 2204 67540 2208
rect 67476 2148 67480 2204
rect 67480 2148 67536 2204
rect 67536 2148 67540 2204
rect 67476 2144 67540 2148
rect 33180 2076 33244 2140
rect 30236 1668 30300 1732
rect 19196 988 19260 1052
<< metal4 >>
rect 5128 37568 5448 37584
rect 5128 37504 5136 37568
rect 5200 37504 5216 37568
rect 5280 37504 5296 37568
rect 5360 37504 5376 37568
rect 5440 37504 5448 37568
rect 5128 36480 5448 37504
rect 5128 36416 5136 36480
rect 5200 36416 5216 36480
rect 5280 36416 5296 36480
rect 5360 36416 5376 36480
rect 5440 36416 5448 36480
rect 5128 35392 5448 36416
rect 5128 35328 5136 35392
rect 5200 35328 5216 35392
rect 5280 35328 5296 35392
rect 5360 35328 5376 35392
rect 5440 35328 5448 35392
rect 5128 34304 5448 35328
rect 5128 34240 5136 34304
rect 5200 34240 5216 34304
rect 5280 34240 5296 34304
rect 5360 34240 5376 34304
rect 5440 34240 5448 34304
rect 5128 33216 5448 34240
rect 5128 33152 5136 33216
rect 5200 33152 5216 33216
rect 5280 33152 5296 33216
rect 5360 33152 5376 33216
rect 5440 33152 5448 33216
rect 5128 32128 5448 33152
rect 5128 32064 5136 32128
rect 5200 32064 5216 32128
rect 5280 32064 5296 32128
rect 5360 32064 5376 32128
rect 5440 32064 5448 32128
rect 5128 31040 5448 32064
rect 5128 30976 5136 31040
rect 5200 30976 5216 31040
rect 5280 30976 5296 31040
rect 5360 30976 5376 31040
rect 5440 30976 5448 31040
rect 5128 29952 5448 30976
rect 5128 29888 5136 29952
rect 5200 29888 5216 29952
rect 5280 29888 5296 29952
rect 5360 29888 5376 29952
rect 5440 29888 5448 29952
rect 5128 28864 5448 29888
rect 5128 28800 5136 28864
rect 5200 28800 5216 28864
rect 5280 28800 5296 28864
rect 5360 28800 5376 28864
rect 5440 28800 5448 28864
rect 5128 27776 5448 28800
rect 5128 27712 5136 27776
rect 5200 27712 5216 27776
rect 5280 27712 5296 27776
rect 5360 27712 5376 27776
rect 5440 27712 5448 27776
rect 5128 26688 5448 27712
rect 5128 26624 5136 26688
rect 5200 26624 5216 26688
rect 5280 26624 5296 26688
rect 5360 26624 5376 26688
rect 5440 26624 5448 26688
rect 5128 25600 5448 26624
rect 5128 25536 5136 25600
rect 5200 25536 5216 25600
rect 5280 25536 5296 25600
rect 5360 25536 5376 25600
rect 5440 25536 5448 25600
rect 5128 24512 5448 25536
rect 5128 24448 5136 24512
rect 5200 24448 5216 24512
rect 5280 24448 5296 24512
rect 5360 24448 5376 24512
rect 5440 24448 5448 24512
rect 5128 23424 5448 24448
rect 5128 23360 5136 23424
rect 5200 23360 5216 23424
rect 5280 23360 5296 23424
rect 5360 23360 5376 23424
rect 5440 23360 5448 23424
rect 5128 22336 5448 23360
rect 5128 22272 5136 22336
rect 5200 22272 5216 22336
rect 5280 22272 5296 22336
rect 5360 22272 5376 22336
rect 5440 22272 5448 22336
rect 5128 21248 5448 22272
rect 5128 21184 5136 21248
rect 5200 21184 5216 21248
rect 5280 21184 5296 21248
rect 5360 21184 5376 21248
rect 5440 21184 5448 21248
rect 5128 20160 5448 21184
rect 5128 20096 5136 20160
rect 5200 20096 5216 20160
rect 5280 20096 5296 20160
rect 5360 20096 5376 20160
rect 5440 20096 5448 20160
rect 5128 19072 5448 20096
rect 5128 19008 5136 19072
rect 5200 19008 5216 19072
rect 5280 19008 5296 19072
rect 5360 19008 5376 19072
rect 5440 19008 5448 19072
rect 5128 17984 5448 19008
rect 5128 17920 5136 17984
rect 5200 17920 5216 17984
rect 5280 17920 5296 17984
rect 5360 17920 5376 17984
rect 5440 17920 5448 17984
rect 5128 16896 5448 17920
rect 5128 16832 5136 16896
rect 5200 16832 5216 16896
rect 5280 16832 5296 16896
rect 5360 16832 5376 16896
rect 5440 16832 5448 16896
rect 5128 15808 5448 16832
rect 5128 15744 5136 15808
rect 5200 15744 5216 15808
rect 5280 15744 5296 15808
rect 5360 15744 5376 15808
rect 5440 15744 5448 15808
rect 5128 14720 5448 15744
rect 5128 14656 5136 14720
rect 5200 14656 5216 14720
rect 5280 14656 5296 14720
rect 5360 14656 5376 14720
rect 5440 14656 5448 14720
rect 5128 13632 5448 14656
rect 5128 13568 5136 13632
rect 5200 13568 5216 13632
rect 5280 13568 5296 13632
rect 5360 13568 5376 13632
rect 5440 13568 5448 13632
rect 5128 12544 5448 13568
rect 5128 12480 5136 12544
rect 5200 12480 5216 12544
rect 5280 12480 5296 12544
rect 5360 12480 5376 12544
rect 5440 12480 5448 12544
rect 5128 11456 5448 12480
rect 5128 11392 5136 11456
rect 5200 11392 5216 11456
rect 5280 11392 5296 11456
rect 5360 11392 5376 11456
rect 5440 11392 5448 11456
rect 5128 10368 5448 11392
rect 5128 10304 5136 10368
rect 5200 10304 5216 10368
rect 5280 10304 5296 10368
rect 5360 10304 5376 10368
rect 5440 10304 5448 10368
rect 5128 9280 5448 10304
rect 5128 9216 5136 9280
rect 5200 9216 5216 9280
rect 5280 9216 5296 9280
rect 5360 9216 5376 9280
rect 5440 9216 5448 9280
rect 4846 3637 4906 8382
rect 5128 8192 5448 9216
rect 5128 8128 5136 8192
rect 5200 8128 5216 8192
rect 5280 8128 5296 8192
rect 5360 8128 5376 8192
rect 5440 8128 5448 8192
rect 5128 7104 5448 8128
rect 5128 7040 5136 7104
rect 5200 7040 5216 7104
rect 5280 7040 5296 7104
rect 5360 7040 5376 7104
rect 5440 7040 5448 7104
rect 5128 6016 5448 7040
rect 5128 5952 5136 6016
rect 5200 5952 5216 6016
rect 5280 5952 5296 6016
rect 5360 5952 5376 6016
rect 5440 5952 5448 6016
rect 5128 4928 5448 5952
rect 5128 4864 5136 4928
rect 5200 4864 5216 4928
rect 5280 4864 5296 4928
rect 5360 4864 5376 4928
rect 5440 4864 5448 4928
rect 5128 3840 5448 4864
rect 5128 3776 5136 3840
rect 5200 3776 5216 3840
rect 5280 3776 5296 3840
rect 5360 3776 5376 3840
rect 5440 3776 5448 3840
rect 4843 3636 4909 3637
rect 4843 3572 4844 3636
rect 4908 3572 4909 3636
rect 4843 3571 4909 3572
rect 5128 2752 5448 3776
rect 5128 2688 5136 2752
rect 5200 2688 5216 2752
rect 5280 2688 5296 2752
rect 5360 2688 5376 2752
rect 5440 2688 5448 2752
rect 5128 2128 5448 2688
rect 5788 37024 6108 37584
rect 5788 36960 5796 37024
rect 5860 36960 5876 37024
rect 5940 36960 5956 37024
rect 6020 36960 6036 37024
rect 6100 36960 6108 37024
rect 5788 35936 6108 36960
rect 35848 37568 36168 37584
rect 35848 37504 35856 37568
rect 35920 37504 35936 37568
rect 36000 37504 36016 37568
rect 36080 37504 36096 37568
rect 36160 37504 36168 37568
rect 7051 36548 7117 36549
rect 7051 36484 7052 36548
rect 7116 36484 7117 36548
rect 7051 36483 7117 36484
rect 32811 36548 32877 36549
rect 32811 36484 32812 36548
rect 32876 36484 32877 36548
rect 32811 36483 32877 36484
rect 5788 35872 5796 35936
rect 5860 35872 5876 35936
rect 5940 35872 5956 35936
rect 6020 35872 6036 35936
rect 6100 35872 6108 35936
rect 5788 34848 6108 35872
rect 5788 34784 5796 34848
rect 5860 34784 5876 34848
rect 5940 34784 5956 34848
rect 6020 34784 6036 34848
rect 6100 34784 6108 34848
rect 5788 33760 6108 34784
rect 5788 33696 5796 33760
rect 5860 33696 5876 33760
rect 5940 33696 5956 33760
rect 6020 33696 6036 33760
rect 6100 33696 6108 33760
rect 5788 32672 6108 33696
rect 5788 32608 5796 32672
rect 5860 32608 5876 32672
rect 5940 32608 5956 32672
rect 6020 32608 6036 32672
rect 6100 32608 6108 32672
rect 5788 31584 6108 32608
rect 5788 31520 5796 31584
rect 5860 31520 5876 31584
rect 5940 31520 5956 31584
rect 6020 31520 6036 31584
rect 6100 31520 6108 31584
rect 5788 30496 6108 31520
rect 5788 30432 5796 30496
rect 5860 30432 5876 30496
rect 5940 30432 5956 30496
rect 6020 30432 6036 30496
rect 6100 30432 6108 30496
rect 5788 29408 6108 30432
rect 5788 29344 5796 29408
rect 5860 29344 5876 29408
rect 5940 29344 5956 29408
rect 6020 29344 6036 29408
rect 6100 29344 6108 29408
rect 5788 28320 6108 29344
rect 5788 28256 5796 28320
rect 5860 28256 5876 28320
rect 5940 28256 5956 28320
rect 6020 28256 6036 28320
rect 6100 28256 6108 28320
rect 5788 27232 6108 28256
rect 5788 27168 5796 27232
rect 5860 27168 5876 27232
rect 5940 27168 5956 27232
rect 6020 27168 6036 27232
rect 6100 27168 6108 27232
rect 5788 26144 6108 27168
rect 5788 26080 5796 26144
rect 5860 26080 5876 26144
rect 5940 26080 5956 26144
rect 6020 26080 6036 26144
rect 6100 26080 6108 26144
rect 5788 25056 6108 26080
rect 5788 24992 5796 25056
rect 5860 24992 5876 25056
rect 5940 24992 5956 25056
rect 6020 24992 6036 25056
rect 6100 24992 6108 25056
rect 5788 23968 6108 24992
rect 5788 23904 5796 23968
rect 5860 23904 5876 23968
rect 5940 23904 5956 23968
rect 6020 23904 6036 23968
rect 6100 23904 6108 23968
rect 5788 22880 6108 23904
rect 5788 22816 5796 22880
rect 5860 22816 5876 22880
rect 5940 22816 5956 22880
rect 6020 22816 6036 22880
rect 6100 22816 6108 22880
rect 5788 21792 6108 22816
rect 5788 21728 5796 21792
rect 5860 21728 5876 21792
rect 5940 21728 5956 21792
rect 6020 21728 6036 21792
rect 6100 21728 6108 21792
rect 5788 20704 6108 21728
rect 5788 20640 5796 20704
rect 5860 20640 5876 20704
rect 5940 20640 5956 20704
rect 6020 20640 6036 20704
rect 6100 20640 6108 20704
rect 5788 19616 6108 20640
rect 5788 19552 5796 19616
rect 5860 19552 5876 19616
rect 5940 19552 5956 19616
rect 6020 19552 6036 19616
rect 6100 19552 6108 19616
rect 5788 18528 6108 19552
rect 5788 18464 5796 18528
rect 5860 18464 5876 18528
rect 5940 18464 5956 18528
rect 6020 18464 6036 18528
rect 6100 18464 6108 18528
rect 5788 17440 6108 18464
rect 5788 17376 5796 17440
rect 5860 17376 5876 17440
rect 5940 17376 5956 17440
rect 6020 17376 6036 17440
rect 6100 17376 6108 17440
rect 5788 16352 6108 17376
rect 5788 16288 5796 16352
rect 5860 16288 5876 16352
rect 5940 16288 5956 16352
rect 6020 16288 6036 16352
rect 6100 16288 6108 16352
rect 5788 15264 6108 16288
rect 5788 15200 5796 15264
rect 5860 15200 5876 15264
rect 5940 15200 5956 15264
rect 6020 15200 6036 15264
rect 6100 15200 6108 15264
rect 5788 14176 6108 15200
rect 5788 14112 5796 14176
rect 5860 14112 5876 14176
rect 5940 14112 5956 14176
rect 6020 14112 6036 14176
rect 6100 14112 6108 14176
rect 5788 13088 6108 14112
rect 5788 13024 5796 13088
rect 5860 13024 5876 13088
rect 5940 13024 5956 13088
rect 6020 13024 6036 13088
rect 6100 13024 6108 13088
rect 5788 12000 6108 13024
rect 5788 11936 5796 12000
rect 5860 11936 5876 12000
rect 5940 11936 5956 12000
rect 6020 11936 6036 12000
rect 6100 11936 6108 12000
rect 5788 10912 6108 11936
rect 5788 10848 5796 10912
rect 5860 10848 5876 10912
rect 5940 10848 5956 10912
rect 6020 10848 6036 10912
rect 6100 10848 6108 10912
rect 5788 9824 6108 10848
rect 5788 9760 5796 9824
rect 5860 9760 5876 9824
rect 5940 9760 5956 9824
rect 6020 9760 6036 9824
rect 6100 9760 6108 9824
rect 5788 8736 6108 9760
rect 5788 8672 5796 8736
rect 5860 8672 5876 8736
rect 5940 8672 5956 8736
rect 6020 8672 6036 8736
rect 6100 8672 6108 8736
rect 5788 7648 6108 8672
rect 7054 7938 7114 36483
rect 27475 29612 27541 29613
rect 27475 29548 27476 29612
rect 27540 29548 27541 29612
rect 27475 29547 27541 29548
rect 27291 18052 27357 18053
rect 27291 17988 27292 18052
rect 27356 17988 27357 18052
rect 27291 17987 27357 17988
rect 27294 16590 27354 17987
rect 27110 16530 27354 16590
rect 12755 12476 12821 12477
rect 12755 12412 12756 12476
rect 12820 12412 12821 12476
rect 12755 12411 12821 12412
rect 10731 10708 10797 10709
rect 10731 10644 10732 10708
rect 10796 10644 10797 10708
rect 10731 10643 10797 10644
rect 5788 7584 5796 7648
rect 5860 7584 5876 7648
rect 5940 7584 5956 7648
rect 6020 7584 6036 7648
rect 6100 7584 6108 7648
rect 5788 6560 6108 7584
rect 5788 6496 5796 6560
rect 5860 6496 5876 6560
rect 5940 6496 5956 6560
rect 6020 6496 6036 6560
rect 6100 6496 6108 6560
rect 5788 5472 6108 6496
rect 5788 5408 5796 5472
rect 5860 5408 5876 5472
rect 5940 5408 5956 5472
rect 6020 5408 6036 5472
rect 6100 5408 6108 5472
rect 5788 4384 6108 5408
rect 5788 4320 5796 4384
rect 5860 4320 5876 4384
rect 5940 4320 5956 4384
rect 6020 4320 6036 4384
rect 6100 4320 6108 4384
rect 5788 3296 6108 4320
rect 5788 3232 5796 3296
rect 5860 3232 5876 3296
rect 5940 3232 5956 3296
rect 6020 3232 6036 3296
rect 6100 3232 6108 3296
rect 5788 2208 6108 3232
rect 10734 2685 10794 10643
rect 10915 10300 10981 10301
rect 10915 10236 10916 10300
rect 10980 10236 10981 10300
rect 10915 10235 10981 10236
rect 10918 4045 10978 10235
rect 10915 4044 10981 4045
rect 10915 3980 10916 4044
rect 10980 3980 10981 4044
rect 10915 3979 10981 3980
rect 11838 3909 11898 10422
rect 12758 4861 12818 12411
rect 19931 11524 19997 11525
rect 19931 11460 19932 11524
rect 19996 11460 19997 11524
rect 19931 11459 19997 11460
rect 17723 11388 17789 11389
rect 17723 11324 17724 11388
rect 17788 11324 17789 11388
rect 17723 11323 17789 11324
rect 15331 11252 15397 11253
rect 15331 11188 15332 11252
rect 15396 11188 15397 11252
rect 15331 11187 15397 11188
rect 13307 11116 13373 11117
rect 13307 11052 13308 11116
rect 13372 11052 13373 11116
rect 13307 11051 13373 11052
rect 13310 5269 13370 11051
rect 13675 7716 13741 7717
rect 13675 7652 13676 7716
rect 13740 7652 13741 7716
rect 13675 7651 13741 7652
rect 13307 5268 13373 5269
rect 13307 5204 13308 5268
rect 13372 5204 13373 5268
rect 13307 5203 13373 5204
rect 12755 4860 12821 4861
rect 12755 4796 12756 4860
rect 12820 4796 12821 4860
rect 12755 4795 12821 4796
rect 13678 3909 13738 7651
rect 15334 5405 15394 11187
rect 17355 10844 17421 10845
rect 17355 10780 17356 10844
rect 17420 10780 17421 10844
rect 17355 10779 17421 10780
rect 16435 10436 16501 10437
rect 16435 10372 16436 10436
rect 16500 10372 16501 10436
rect 16435 10371 16501 10372
rect 16438 6085 16498 10371
rect 17171 8124 17237 8125
rect 17171 8060 17172 8124
rect 17236 8060 17237 8124
rect 17171 8059 17237 8060
rect 17174 6221 17234 8059
rect 17171 6220 17237 6221
rect 17171 6156 17172 6220
rect 17236 6156 17237 6220
rect 17171 6155 17237 6156
rect 16067 6084 16133 6085
rect 16067 6020 16068 6084
rect 16132 6020 16133 6084
rect 16067 6019 16133 6020
rect 16435 6084 16501 6085
rect 16435 6020 16436 6084
rect 16500 6020 16501 6084
rect 16435 6019 16501 6020
rect 16987 6084 17053 6085
rect 16987 6020 16988 6084
rect 17052 6020 17053 6084
rect 16987 6019 17053 6020
rect 15331 5404 15397 5405
rect 15331 5340 15332 5404
rect 15396 5340 15397 5404
rect 15331 5339 15397 5340
rect 11835 3908 11901 3909
rect 11835 3844 11836 3908
rect 11900 3844 11901 3908
rect 11835 3843 11901 3844
rect 13675 3908 13741 3909
rect 13675 3844 13676 3908
rect 13740 3844 13741 3908
rect 16070 3858 16130 6019
rect 16990 3909 17050 6019
rect 17358 4861 17418 10779
rect 17726 4861 17786 11323
rect 18091 10164 18157 10165
rect 18091 10100 18092 10164
rect 18156 10100 18157 10164
rect 18091 10099 18157 10100
rect 17907 8804 17973 8805
rect 17907 8740 17908 8804
rect 17972 8740 17973 8804
rect 17907 8739 17973 8740
rect 17355 4860 17421 4861
rect 17355 4796 17356 4860
rect 17420 4796 17421 4860
rect 17355 4795 17421 4796
rect 17723 4860 17789 4861
rect 17723 4796 17724 4860
rect 17788 4796 17789 4860
rect 17723 4795 17789 4796
rect 16987 3908 17053 3909
rect 13675 3843 13741 3844
rect 16987 3844 16988 3908
rect 17052 3844 17053 3908
rect 16987 3843 17053 3844
rect 16070 3365 16130 3622
rect 16067 3364 16133 3365
rect 16067 3300 16068 3364
rect 16132 3300 16133 3364
rect 16067 3299 16133 3300
rect 10731 2684 10797 2685
rect 10731 2620 10732 2684
rect 10796 2620 10797 2684
rect 10731 2619 10797 2620
rect 17910 2549 17970 8739
rect 18094 6085 18154 10099
rect 19747 9620 19813 9621
rect 19747 9556 19748 9620
rect 19812 9556 19813 9620
rect 19747 9555 19813 9556
rect 18643 8804 18709 8805
rect 18643 8740 18644 8804
rect 18708 8740 18709 8804
rect 18643 8739 18709 8740
rect 18275 8532 18341 8533
rect 18275 8468 18276 8532
rect 18340 8468 18341 8532
rect 18275 8467 18341 8468
rect 18091 6084 18157 6085
rect 18091 6020 18092 6084
rect 18156 6020 18157 6084
rect 18091 6019 18157 6020
rect 18278 2685 18338 8467
rect 18459 8396 18525 8397
rect 18459 8332 18460 8396
rect 18524 8332 18525 8396
rect 18459 8331 18525 8332
rect 18275 2684 18341 2685
rect 18275 2620 18276 2684
rect 18340 2620 18341 2684
rect 18275 2619 18341 2620
rect 17907 2548 17973 2549
rect 17907 2484 17908 2548
rect 17972 2484 17973 2548
rect 17907 2483 17973 2484
rect 18462 2413 18522 8331
rect 18646 6085 18706 8739
rect 18643 6084 18709 6085
rect 18643 6020 18644 6084
rect 18708 6020 18709 6084
rect 18643 6019 18709 6020
rect 19195 5812 19261 5813
rect 19195 5748 19196 5812
rect 19260 5748 19261 5812
rect 19195 5747 19261 5748
rect 18459 2412 18525 2413
rect 18459 2348 18460 2412
rect 18524 2348 18525 2412
rect 18459 2347 18525 2348
rect 5788 2144 5796 2208
rect 5860 2144 5876 2208
rect 5940 2144 5956 2208
rect 6020 2144 6036 2208
rect 6100 2144 6108 2208
rect 5788 2128 6108 2144
rect 19198 1053 19258 5747
rect 19750 4861 19810 9555
rect 19934 5813 19994 11459
rect 26555 11116 26621 11117
rect 26555 11052 26556 11116
rect 26620 11052 26621 11116
rect 26555 11051 26621 11052
rect 23059 10300 23125 10301
rect 23059 10236 23060 10300
rect 23124 10236 23125 10300
rect 23059 10235 23125 10236
rect 21771 10028 21837 10029
rect 21771 9964 21772 10028
rect 21836 9964 21837 10028
rect 21771 9963 21837 9964
rect 22691 10028 22757 10029
rect 22691 9964 22692 10028
rect 22756 9964 22757 10028
rect 22691 9963 22757 9964
rect 20667 8396 20733 8397
rect 20667 8332 20668 8396
rect 20732 8332 20733 8396
rect 20667 8331 20733 8332
rect 20115 7852 20181 7853
rect 20115 7788 20116 7852
rect 20180 7788 20181 7852
rect 20115 7787 20181 7788
rect 19931 5812 19997 5813
rect 19931 5748 19932 5812
rect 19996 5748 19997 5812
rect 19931 5747 19997 5748
rect 19747 4860 19813 4861
rect 19747 4796 19748 4860
rect 19812 4796 19813 4860
rect 19747 4795 19813 4796
rect 20118 4453 20178 7787
rect 20670 5949 20730 8331
rect 21219 7308 21285 7309
rect 21219 7244 21220 7308
rect 21284 7244 21285 7308
rect 21219 7243 21285 7244
rect 20667 5948 20733 5949
rect 20667 5884 20668 5948
rect 20732 5884 20733 5948
rect 20667 5883 20733 5884
rect 21222 5813 21282 7243
rect 21219 5812 21285 5813
rect 21219 5748 21220 5812
rect 21284 5748 21285 5812
rect 21219 5747 21285 5748
rect 20115 4452 20181 4453
rect 20115 4388 20116 4452
rect 20180 4388 20181 4452
rect 20115 4387 20181 4388
rect 21774 4045 21834 9963
rect 22139 6492 22205 6493
rect 22139 6428 22140 6492
rect 22204 6428 22205 6492
rect 22139 6427 22205 6428
rect 22142 5269 22202 6427
rect 22694 5677 22754 9963
rect 22691 5676 22757 5677
rect 22691 5612 22692 5676
rect 22756 5612 22757 5676
rect 22691 5611 22757 5612
rect 22139 5268 22205 5269
rect 22139 5204 22140 5268
rect 22204 5204 22205 5268
rect 22139 5203 22205 5204
rect 23062 4045 23122 10235
rect 23795 10028 23861 10029
rect 23795 9964 23796 10028
rect 23860 9964 23861 10028
rect 23795 9963 23861 9964
rect 23427 7444 23493 7445
rect 23427 7380 23428 7444
rect 23492 7380 23493 7444
rect 23427 7379 23493 7380
rect 21771 4044 21837 4045
rect 21771 3980 21772 4044
rect 21836 3980 21837 4044
rect 21771 3979 21837 3980
rect 23059 4044 23125 4045
rect 23059 3980 23060 4044
rect 23124 3980 23125 4044
rect 23059 3979 23125 3980
rect 23430 3229 23490 7379
rect 23798 5949 23858 9963
rect 24899 9756 24965 9757
rect 24899 9692 24900 9756
rect 24964 9692 24965 9756
rect 24899 9691 24965 9692
rect 24163 9348 24229 9349
rect 24163 9284 24164 9348
rect 24228 9284 24229 9348
rect 24163 9283 24229 9284
rect 23795 5948 23861 5949
rect 23795 5884 23796 5948
rect 23860 5884 23861 5948
rect 23795 5883 23861 5884
rect 24166 5541 24226 9283
rect 24715 9076 24781 9077
rect 24715 9012 24716 9076
rect 24780 9012 24781 9076
rect 24715 9011 24781 9012
rect 24163 5540 24229 5541
rect 24163 5476 24164 5540
rect 24228 5476 24229 5540
rect 24163 5475 24229 5476
rect 24718 4181 24778 9011
rect 24902 7989 24962 9691
rect 25267 8532 25333 8533
rect 25267 8468 25268 8532
rect 25332 8468 25333 8532
rect 25267 8467 25333 8468
rect 24899 7988 24965 7989
rect 24899 7924 24900 7988
rect 24964 7924 24965 7988
rect 24899 7923 24965 7924
rect 25270 4538 25330 8467
rect 25819 8396 25885 8397
rect 25819 8332 25820 8396
rect 25884 8332 25885 8396
rect 25819 8331 25885 8332
rect 24715 4180 24781 4181
rect 24715 4116 24716 4180
rect 24780 4116 24781 4180
rect 24715 4115 24781 4116
rect 25270 3229 25330 4302
rect 25822 4045 25882 8331
rect 26558 4045 26618 11051
rect 27110 7717 27170 16530
rect 27478 12450 27538 29547
rect 28395 26892 28461 26893
rect 28395 26828 28396 26892
rect 28460 26828 28461 26892
rect 28395 26827 28461 26828
rect 28211 14380 28277 14381
rect 28211 14316 28212 14380
rect 28276 14316 28277 14380
rect 28211 14315 28277 14316
rect 27294 12390 27538 12450
rect 27107 7716 27173 7717
rect 27107 7652 27108 7716
rect 27172 7652 27173 7716
rect 27107 7651 27173 7652
rect 27294 7581 27354 12390
rect 27475 8396 27541 8397
rect 27475 8332 27476 8396
rect 27540 8332 27541 8396
rect 27475 8331 27541 8332
rect 27291 7580 27357 7581
rect 27291 7516 27292 7580
rect 27356 7516 27357 7580
rect 27291 7515 27357 7516
rect 27291 7172 27357 7173
rect 27291 7108 27292 7172
rect 27356 7108 27357 7172
rect 27291 7107 27357 7108
rect 25819 4044 25885 4045
rect 25819 3980 25820 4044
rect 25884 3980 25885 4044
rect 25819 3979 25885 3980
rect 26555 4044 26621 4045
rect 26555 3980 26556 4044
rect 26620 3980 26621 4044
rect 26555 3979 26621 3980
rect 23427 3228 23493 3229
rect 23427 3164 23428 3228
rect 23492 3164 23493 3228
rect 23427 3163 23493 3164
rect 25267 3228 25333 3229
rect 25267 3164 25268 3228
rect 25332 3164 25333 3228
rect 25267 3163 25333 3164
rect 27294 3093 27354 7107
rect 27478 5541 27538 8331
rect 28214 7989 28274 14315
rect 28211 7988 28277 7989
rect 28211 7924 28212 7988
rect 28276 7924 28277 7988
rect 28211 7923 28277 7924
rect 28398 5949 28458 26827
rect 28579 14516 28645 14517
rect 28579 14452 28580 14516
rect 28644 14452 28645 14516
rect 28579 14451 28645 14452
rect 28582 6085 28642 14451
rect 30971 10436 31037 10437
rect 30971 10372 30972 10436
rect 31036 10372 31037 10436
rect 30971 10371 31037 10372
rect 29131 9756 29197 9757
rect 29131 9692 29132 9756
rect 29196 9692 29197 9756
rect 29131 9691 29197 9692
rect 30235 9756 30301 9757
rect 30235 9692 30236 9756
rect 30300 9692 30301 9756
rect 30235 9691 30301 9692
rect 28947 9620 29013 9621
rect 28947 9556 28948 9620
rect 29012 9556 29013 9620
rect 28947 9555 29013 9556
rect 28763 8940 28829 8941
rect 28763 8876 28764 8940
rect 28828 8876 28829 8940
rect 28763 8875 28829 8876
rect 28579 6084 28645 6085
rect 28579 6020 28580 6084
rect 28644 6020 28645 6084
rect 28579 6019 28645 6020
rect 28395 5948 28461 5949
rect 28395 5884 28396 5948
rect 28460 5884 28461 5948
rect 28395 5883 28461 5884
rect 27475 5540 27541 5541
rect 27475 5476 27476 5540
rect 27540 5476 27541 5540
rect 27475 5475 27541 5476
rect 28582 3637 28642 6019
rect 28766 4861 28826 8875
rect 28950 4997 29010 9555
rect 29134 5405 29194 9691
rect 29315 9076 29381 9077
rect 29315 9012 29316 9076
rect 29380 9012 29381 9076
rect 29315 9011 29381 9012
rect 29131 5404 29197 5405
rect 29131 5340 29132 5404
rect 29196 5340 29197 5404
rect 29131 5339 29197 5340
rect 28947 4996 29013 4997
rect 28947 4932 28948 4996
rect 29012 4932 29013 4996
rect 28947 4931 29013 4932
rect 28763 4860 28829 4861
rect 28763 4796 28764 4860
rect 28828 4796 28829 4860
rect 28763 4795 28829 4796
rect 29318 4181 29378 9011
rect 29315 4180 29381 4181
rect 29315 4116 29316 4180
rect 29380 4116 29381 4180
rect 29315 4115 29381 4116
rect 28579 3636 28645 3637
rect 28579 3572 28580 3636
rect 28644 3572 28645 3636
rect 28579 3571 28645 3572
rect 27291 3092 27357 3093
rect 27291 3028 27292 3092
rect 27356 3028 27357 3092
rect 27291 3027 27357 3028
rect 30238 1733 30298 9691
rect 30974 6901 31034 10371
rect 31155 8532 31221 8533
rect 31155 8468 31156 8532
rect 31220 8468 31221 8532
rect 31155 8467 31221 8468
rect 30971 6900 31037 6901
rect 30971 6836 30972 6900
rect 31036 6836 31037 6900
rect 30971 6835 31037 6836
rect 31158 2821 31218 8467
rect 31891 8396 31957 8397
rect 31891 8332 31892 8396
rect 31956 8332 31957 8396
rect 31891 8331 31957 8332
rect 31894 3365 31954 8331
rect 32259 7852 32325 7853
rect 32259 7788 32260 7852
rect 32324 7788 32325 7852
rect 32259 7787 32325 7788
rect 32262 5269 32322 7787
rect 32814 7309 32874 36483
rect 35848 36480 36168 37504
rect 35848 36416 35856 36480
rect 35920 36416 35936 36480
rect 36000 36416 36016 36480
rect 36080 36416 36096 36480
rect 36160 36416 36168 36480
rect 35848 35392 36168 36416
rect 35848 35328 35856 35392
rect 35920 35328 35936 35392
rect 36000 35328 36016 35392
rect 36080 35328 36096 35392
rect 36160 35328 36168 35392
rect 35848 34304 36168 35328
rect 35848 34240 35856 34304
rect 35920 34240 35936 34304
rect 36000 34240 36016 34304
rect 36080 34240 36096 34304
rect 36160 34240 36168 34304
rect 35848 33216 36168 34240
rect 35848 33152 35856 33216
rect 35920 33152 35936 33216
rect 36000 33152 36016 33216
rect 36080 33152 36096 33216
rect 36160 33152 36168 33216
rect 35848 32128 36168 33152
rect 35848 32064 35856 32128
rect 35920 32064 35936 32128
rect 36000 32064 36016 32128
rect 36080 32064 36096 32128
rect 36160 32064 36168 32128
rect 35848 31040 36168 32064
rect 35848 30976 35856 31040
rect 35920 30976 35936 31040
rect 36000 30976 36016 31040
rect 36080 30976 36096 31040
rect 36160 30976 36168 31040
rect 35848 29952 36168 30976
rect 35848 29888 35856 29952
rect 35920 29888 35936 29952
rect 36000 29888 36016 29952
rect 36080 29888 36096 29952
rect 36160 29888 36168 29952
rect 35848 28864 36168 29888
rect 35848 28800 35856 28864
rect 35920 28800 35936 28864
rect 36000 28800 36016 28864
rect 36080 28800 36096 28864
rect 36160 28800 36168 28864
rect 35848 27776 36168 28800
rect 35848 27712 35856 27776
rect 35920 27712 35936 27776
rect 36000 27712 36016 27776
rect 36080 27712 36096 27776
rect 36160 27712 36168 27776
rect 35848 26688 36168 27712
rect 35848 26624 35856 26688
rect 35920 26624 35936 26688
rect 36000 26624 36016 26688
rect 36080 26624 36096 26688
rect 36160 26624 36168 26688
rect 35848 25600 36168 26624
rect 35848 25536 35856 25600
rect 35920 25536 35936 25600
rect 36000 25536 36016 25600
rect 36080 25536 36096 25600
rect 36160 25536 36168 25600
rect 35848 24512 36168 25536
rect 35848 24448 35856 24512
rect 35920 24448 35936 24512
rect 36000 24448 36016 24512
rect 36080 24448 36096 24512
rect 36160 24448 36168 24512
rect 35019 24172 35085 24173
rect 35019 24108 35020 24172
rect 35084 24108 35085 24172
rect 35019 24107 35085 24108
rect 33363 8532 33429 8533
rect 33363 8468 33364 8532
rect 33428 8468 33429 8532
rect 33363 8467 33429 8468
rect 33179 8396 33245 8397
rect 33179 8332 33180 8396
rect 33244 8332 33245 8396
rect 33179 8331 33245 8332
rect 32811 7308 32877 7309
rect 32811 7244 32812 7308
rect 32876 7244 32877 7308
rect 32811 7243 32877 7244
rect 32259 5268 32325 5269
rect 32259 5204 32260 5268
rect 32324 5204 32325 5268
rect 32259 5203 32325 5204
rect 31891 3364 31957 3365
rect 31891 3300 31892 3364
rect 31956 3300 31957 3364
rect 31891 3299 31957 3300
rect 31155 2820 31221 2821
rect 31155 2756 31156 2820
rect 31220 2756 31221 2820
rect 31155 2755 31221 2756
rect 33182 2141 33242 8331
rect 33366 2549 33426 8467
rect 33731 8396 33797 8397
rect 33731 8332 33732 8396
rect 33796 8332 33797 8396
rect 33731 8331 33797 8332
rect 33547 7988 33613 7989
rect 33547 7924 33548 7988
rect 33612 7924 33613 7988
rect 33547 7923 33613 7924
rect 33550 2685 33610 7923
rect 33547 2684 33613 2685
rect 33547 2620 33548 2684
rect 33612 2620 33613 2684
rect 33547 2619 33613 2620
rect 33363 2548 33429 2549
rect 33363 2484 33364 2548
rect 33428 2484 33429 2548
rect 33734 2498 33794 8331
rect 34467 7716 34533 7717
rect 34467 7652 34468 7716
rect 34532 7652 34533 7716
rect 34467 7651 34533 7652
rect 33363 2483 33429 2484
rect 34470 2277 34530 7651
rect 35022 6901 35082 24107
rect 35848 23424 36168 24448
rect 35848 23360 35856 23424
rect 35920 23360 35936 23424
rect 36000 23360 36016 23424
rect 36080 23360 36096 23424
rect 36160 23360 36168 23424
rect 35848 22336 36168 23360
rect 35848 22272 35856 22336
rect 35920 22272 35936 22336
rect 36000 22272 36016 22336
rect 36080 22272 36096 22336
rect 36160 22272 36168 22336
rect 35848 21248 36168 22272
rect 35848 21184 35856 21248
rect 35920 21184 35936 21248
rect 36000 21184 36016 21248
rect 36080 21184 36096 21248
rect 36160 21184 36168 21248
rect 35848 20160 36168 21184
rect 35848 20096 35856 20160
rect 35920 20096 35936 20160
rect 36000 20096 36016 20160
rect 36080 20096 36096 20160
rect 36160 20096 36168 20160
rect 35848 19072 36168 20096
rect 35848 19008 35856 19072
rect 35920 19008 35936 19072
rect 36000 19008 36016 19072
rect 36080 19008 36096 19072
rect 36160 19008 36168 19072
rect 35848 17984 36168 19008
rect 35848 17920 35856 17984
rect 35920 17920 35936 17984
rect 36000 17920 36016 17984
rect 36080 17920 36096 17984
rect 36160 17920 36168 17984
rect 35848 16896 36168 17920
rect 35848 16832 35856 16896
rect 35920 16832 35936 16896
rect 36000 16832 36016 16896
rect 36080 16832 36096 16896
rect 36160 16832 36168 16896
rect 35848 15808 36168 16832
rect 35848 15744 35856 15808
rect 35920 15744 35936 15808
rect 36000 15744 36016 15808
rect 36080 15744 36096 15808
rect 36160 15744 36168 15808
rect 35848 14720 36168 15744
rect 35848 14656 35856 14720
rect 35920 14656 35936 14720
rect 36000 14656 36016 14720
rect 36080 14656 36096 14720
rect 36160 14656 36168 14720
rect 35848 13632 36168 14656
rect 35848 13568 35856 13632
rect 35920 13568 35936 13632
rect 36000 13568 36016 13632
rect 36080 13568 36096 13632
rect 36160 13568 36168 13632
rect 35848 12544 36168 13568
rect 35848 12480 35856 12544
rect 35920 12480 35936 12544
rect 36000 12480 36016 12544
rect 36080 12480 36096 12544
rect 36160 12480 36168 12544
rect 35848 11456 36168 12480
rect 35848 11392 35856 11456
rect 35920 11392 35936 11456
rect 36000 11392 36016 11456
rect 36080 11392 36096 11456
rect 36160 11392 36168 11456
rect 35848 10368 36168 11392
rect 35848 10304 35856 10368
rect 35920 10304 35936 10368
rect 36000 10304 36016 10368
rect 36080 10304 36096 10368
rect 36160 10304 36168 10368
rect 35848 9280 36168 10304
rect 35848 9216 35856 9280
rect 35920 9216 35936 9280
rect 36000 9216 36016 9280
rect 36080 9216 36096 9280
rect 36160 9216 36168 9280
rect 35848 8192 36168 9216
rect 35848 8128 35856 8192
rect 35920 8128 35936 8192
rect 36000 8128 36016 8192
rect 36080 8128 36096 8192
rect 36160 8128 36168 8192
rect 35848 7104 36168 8128
rect 35848 7040 35856 7104
rect 35920 7040 35936 7104
rect 36000 7040 36016 7104
rect 36080 7040 36096 7104
rect 36160 7040 36168 7104
rect 35019 6900 35085 6901
rect 35019 6836 35020 6900
rect 35084 6836 35085 6900
rect 35019 6835 35085 6836
rect 35848 6016 36168 7040
rect 35848 5952 35856 6016
rect 35920 5952 35936 6016
rect 36000 5952 36016 6016
rect 36080 5952 36096 6016
rect 36160 5952 36168 6016
rect 35848 4928 36168 5952
rect 35848 4864 35856 4928
rect 35920 4864 35936 4928
rect 36000 4864 36016 4928
rect 36080 4864 36096 4928
rect 36160 4864 36168 4928
rect 35848 3840 36168 4864
rect 35848 3776 35856 3840
rect 35920 3776 35936 3840
rect 36000 3776 36016 3840
rect 36080 3776 36096 3840
rect 36160 3776 36168 3840
rect 35848 2752 36168 3776
rect 35848 2688 35856 2752
rect 35920 2688 35936 2752
rect 36000 2688 36016 2752
rect 36080 2688 36096 2752
rect 36160 2688 36168 2752
rect 34467 2276 34533 2277
rect 34467 2212 34468 2276
rect 34532 2212 34533 2276
rect 34467 2211 34533 2212
rect 33179 2140 33245 2141
rect 33179 2076 33180 2140
rect 33244 2076 33245 2140
rect 35848 2128 36168 2688
rect 36508 37024 36828 37584
rect 36508 36960 36516 37024
rect 36580 36960 36596 37024
rect 36660 36960 36676 37024
rect 36740 36960 36756 37024
rect 36820 36960 36828 37024
rect 36508 35936 36828 36960
rect 36508 35872 36516 35936
rect 36580 35872 36596 35936
rect 36660 35872 36676 35936
rect 36740 35872 36756 35936
rect 36820 35872 36828 35936
rect 36508 34848 36828 35872
rect 36508 34784 36516 34848
rect 36580 34784 36596 34848
rect 36660 34784 36676 34848
rect 36740 34784 36756 34848
rect 36820 34784 36828 34848
rect 36508 33760 36828 34784
rect 36508 33696 36516 33760
rect 36580 33696 36596 33760
rect 36660 33696 36676 33760
rect 36740 33696 36756 33760
rect 36820 33696 36828 33760
rect 36508 32672 36828 33696
rect 36508 32608 36516 32672
rect 36580 32608 36596 32672
rect 36660 32608 36676 32672
rect 36740 32608 36756 32672
rect 36820 32608 36828 32672
rect 36508 31584 36828 32608
rect 36508 31520 36516 31584
rect 36580 31520 36596 31584
rect 36660 31520 36676 31584
rect 36740 31520 36756 31584
rect 36820 31520 36828 31584
rect 36508 30496 36828 31520
rect 36508 30432 36516 30496
rect 36580 30432 36596 30496
rect 36660 30432 36676 30496
rect 36740 30432 36756 30496
rect 36820 30432 36828 30496
rect 36508 29408 36828 30432
rect 36508 29344 36516 29408
rect 36580 29344 36596 29408
rect 36660 29344 36676 29408
rect 36740 29344 36756 29408
rect 36820 29344 36828 29408
rect 36508 28320 36828 29344
rect 36508 28256 36516 28320
rect 36580 28256 36596 28320
rect 36660 28256 36676 28320
rect 36740 28256 36756 28320
rect 36820 28256 36828 28320
rect 36508 27232 36828 28256
rect 36508 27168 36516 27232
rect 36580 27168 36596 27232
rect 36660 27168 36676 27232
rect 36740 27168 36756 27232
rect 36820 27168 36828 27232
rect 36508 26144 36828 27168
rect 36508 26080 36516 26144
rect 36580 26080 36596 26144
rect 36660 26080 36676 26144
rect 36740 26080 36756 26144
rect 36820 26080 36828 26144
rect 36508 25056 36828 26080
rect 36508 24992 36516 25056
rect 36580 24992 36596 25056
rect 36660 24992 36676 25056
rect 36740 24992 36756 25056
rect 36820 24992 36828 25056
rect 36508 23968 36828 24992
rect 36508 23904 36516 23968
rect 36580 23904 36596 23968
rect 36660 23904 36676 23968
rect 36740 23904 36756 23968
rect 36820 23904 36828 23968
rect 36508 22880 36828 23904
rect 36508 22816 36516 22880
rect 36580 22816 36596 22880
rect 36660 22816 36676 22880
rect 36740 22816 36756 22880
rect 36820 22816 36828 22880
rect 36508 21792 36828 22816
rect 36508 21728 36516 21792
rect 36580 21728 36596 21792
rect 36660 21728 36676 21792
rect 36740 21728 36756 21792
rect 36820 21728 36828 21792
rect 36508 20704 36828 21728
rect 36508 20640 36516 20704
rect 36580 20640 36596 20704
rect 36660 20640 36676 20704
rect 36740 20640 36756 20704
rect 36820 20640 36828 20704
rect 36508 19616 36828 20640
rect 36508 19552 36516 19616
rect 36580 19552 36596 19616
rect 36660 19552 36676 19616
rect 36740 19552 36756 19616
rect 36820 19552 36828 19616
rect 36508 18528 36828 19552
rect 36508 18464 36516 18528
rect 36580 18464 36596 18528
rect 36660 18464 36676 18528
rect 36740 18464 36756 18528
rect 36820 18464 36828 18528
rect 36508 17440 36828 18464
rect 36508 17376 36516 17440
rect 36580 17376 36596 17440
rect 36660 17376 36676 17440
rect 36740 17376 36756 17440
rect 36820 17376 36828 17440
rect 36508 16352 36828 17376
rect 36508 16288 36516 16352
rect 36580 16288 36596 16352
rect 36660 16288 36676 16352
rect 36740 16288 36756 16352
rect 36820 16288 36828 16352
rect 36508 15264 36828 16288
rect 36508 15200 36516 15264
rect 36580 15200 36596 15264
rect 36660 15200 36676 15264
rect 36740 15200 36756 15264
rect 36820 15200 36828 15264
rect 36508 14176 36828 15200
rect 36508 14112 36516 14176
rect 36580 14112 36596 14176
rect 36660 14112 36676 14176
rect 36740 14112 36756 14176
rect 36820 14112 36828 14176
rect 36508 13088 36828 14112
rect 36508 13024 36516 13088
rect 36580 13024 36596 13088
rect 36660 13024 36676 13088
rect 36740 13024 36756 13088
rect 36820 13024 36828 13088
rect 36508 12000 36828 13024
rect 36508 11936 36516 12000
rect 36580 11936 36596 12000
rect 36660 11936 36676 12000
rect 36740 11936 36756 12000
rect 36820 11936 36828 12000
rect 36508 10912 36828 11936
rect 36508 10848 36516 10912
rect 36580 10848 36596 10912
rect 36660 10848 36676 10912
rect 36740 10848 36756 10912
rect 36820 10848 36828 10912
rect 36508 9824 36828 10848
rect 36508 9760 36516 9824
rect 36580 9760 36596 9824
rect 36660 9760 36676 9824
rect 36740 9760 36756 9824
rect 36820 9760 36828 9824
rect 36508 8736 36828 9760
rect 36508 8672 36516 8736
rect 36580 8672 36596 8736
rect 36660 8672 36676 8736
rect 36740 8672 36756 8736
rect 36820 8672 36828 8736
rect 36508 7648 36828 8672
rect 66568 37568 66888 37584
rect 66568 37504 66576 37568
rect 66640 37504 66656 37568
rect 66720 37504 66736 37568
rect 66800 37504 66816 37568
rect 66880 37504 66888 37568
rect 66568 36480 66888 37504
rect 66568 36416 66576 36480
rect 66640 36416 66656 36480
rect 66720 36416 66736 36480
rect 66800 36416 66816 36480
rect 66880 36416 66888 36480
rect 66568 35392 66888 36416
rect 66568 35328 66576 35392
rect 66640 35328 66656 35392
rect 66720 35328 66736 35392
rect 66800 35328 66816 35392
rect 66880 35328 66888 35392
rect 66568 34304 66888 35328
rect 66568 34240 66576 34304
rect 66640 34240 66656 34304
rect 66720 34240 66736 34304
rect 66800 34240 66816 34304
rect 66880 34240 66888 34304
rect 66568 33216 66888 34240
rect 66568 33152 66576 33216
rect 66640 33152 66656 33216
rect 66720 33152 66736 33216
rect 66800 33152 66816 33216
rect 66880 33152 66888 33216
rect 66568 32128 66888 33152
rect 66568 32064 66576 32128
rect 66640 32064 66656 32128
rect 66720 32064 66736 32128
rect 66800 32064 66816 32128
rect 66880 32064 66888 32128
rect 66568 31040 66888 32064
rect 66568 30976 66576 31040
rect 66640 30976 66656 31040
rect 66720 30976 66736 31040
rect 66800 30976 66816 31040
rect 66880 30976 66888 31040
rect 66568 29952 66888 30976
rect 66568 29888 66576 29952
rect 66640 29888 66656 29952
rect 66720 29888 66736 29952
rect 66800 29888 66816 29952
rect 66880 29888 66888 29952
rect 66568 28864 66888 29888
rect 66568 28800 66576 28864
rect 66640 28800 66656 28864
rect 66720 28800 66736 28864
rect 66800 28800 66816 28864
rect 66880 28800 66888 28864
rect 66568 27776 66888 28800
rect 66568 27712 66576 27776
rect 66640 27712 66656 27776
rect 66720 27712 66736 27776
rect 66800 27712 66816 27776
rect 66880 27712 66888 27776
rect 66568 26688 66888 27712
rect 66568 26624 66576 26688
rect 66640 26624 66656 26688
rect 66720 26624 66736 26688
rect 66800 26624 66816 26688
rect 66880 26624 66888 26688
rect 66568 25600 66888 26624
rect 66568 25536 66576 25600
rect 66640 25536 66656 25600
rect 66720 25536 66736 25600
rect 66800 25536 66816 25600
rect 66880 25536 66888 25600
rect 66568 24512 66888 25536
rect 66568 24448 66576 24512
rect 66640 24448 66656 24512
rect 66720 24448 66736 24512
rect 66800 24448 66816 24512
rect 66880 24448 66888 24512
rect 66568 23424 66888 24448
rect 66568 23360 66576 23424
rect 66640 23360 66656 23424
rect 66720 23360 66736 23424
rect 66800 23360 66816 23424
rect 66880 23360 66888 23424
rect 66568 22336 66888 23360
rect 66568 22272 66576 22336
rect 66640 22272 66656 22336
rect 66720 22272 66736 22336
rect 66800 22272 66816 22336
rect 66880 22272 66888 22336
rect 66568 21248 66888 22272
rect 66568 21184 66576 21248
rect 66640 21184 66656 21248
rect 66720 21184 66736 21248
rect 66800 21184 66816 21248
rect 66880 21184 66888 21248
rect 66568 20160 66888 21184
rect 66568 20096 66576 20160
rect 66640 20096 66656 20160
rect 66720 20096 66736 20160
rect 66800 20096 66816 20160
rect 66880 20096 66888 20160
rect 66568 19072 66888 20096
rect 66568 19008 66576 19072
rect 66640 19008 66656 19072
rect 66720 19008 66736 19072
rect 66800 19008 66816 19072
rect 66880 19008 66888 19072
rect 66568 17984 66888 19008
rect 66568 17920 66576 17984
rect 66640 17920 66656 17984
rect 66720 17920 66736 17984
rect 66800 17920 66816 17984
rect 66880 17920 66888 17984
rect 66568 16896 66888 17920
rect 66568 16832 66576 16896
rect 66640 16832 66656 16896
rect 66720 16832 66736 16896
rect 66800 16832 66816 16896
rect 66880 16832 66888 16896
rect 66568 15808 66888 16832
rect 66568 15744 66576 15808
rect 66640 15744 66656 15808
rect 66720 15744 66736 15808
rect 66800 15744 66816 15808
rect 66880 15744 66888 15808
rect 66568 14720 66888 15744
rect 66568 14656 66576 14720
rect 66640 14656 66656 14720
rect 66720 14656 66736 14720
rect 66800 14656 66816 14720
rect 66880 14656 66888 14720
rect 66568 13632 66888 14656
rect 66568 13568 66576 13632
rect 66640 13568 66656 13632
rect 66720 13568 66736 13632
rect 66800 13568 66816 13632
rect 66880 13568 66888 13632
rect 66568 12544 66888 13568
rect 66568 12480 66576 12544
rect 66640 12480 66656 12544
rect 66720 12480 66736 12544
rect 66800 12480 66816 12544
rect 66880 12480 66888 12544
rect 66568 11456 66888 12480
rect 66568 11392 66576 11456
rect 66640 11392 66656 11456
rect 66720 11392 66736 11456
rect 66800 11392 66816 11456
rect 66880 11392 66888 11456
rect 66568 10368 66888 11392
rect 66568 10304 66576 10368
rect 66640 10304 66656 10368
rect 66720 10304 66736 10368
rect 66800 10304 66816 10368
rect 66880 10304 66888 10368
rect 66568 9280 66888 10304
rect 66568 9216 66576 9280
rect 66640 9216 66656 9280
rect 66720 9216 66736 9280
rect 66800 9216 66816 9280
rect 66880 9216 66888 9280
rect 37043 8532 37109 8533
rect 37043 8468 37044 8532
rect 37108 8468 37109 8532
rect 37043 8467 37109 8468
rect 36508 7584 36516 7648
rect 36580 7584 36596 7648
rect 36660 7584 36676 7648
rect 36740 7584 36756 7648
rect 36820 7584 36828 7648
rect 36508 6560 36828 7584
rect 36508 6496 36516 6560
rect 36580 6496 36596 6560
rect 36660 6496 36676 6560
rect 36740 6496 36756 6560
rect 36820 6496 36828 6560
rect 36508 5472 36828 6496
rect 36508 5408 36516 5472
rect 36580 5408 36596 5472
rect 36660 5408 36676 5472
rect 36740 5408 36756 5472
rect 36820 5408 36828 5472
rect 36508 4384 36828 5408
rect 36508 4320 36516 4384
rect 36580 4320 36596 4384
rect 36660 4320 36676 4384
rect 36740 4320 36756 4384
rect 36820 4320 36828 4384
rect 36508 3296 36828 4320
rect 36508 3232 36516 3296
rect 36580 3232 36596 3296
rect 36660 3232 36676 3296
rect 36740 3232 36756 3296
rect 36820 3232 36828 3296
rect 36508 2208 36828 3232
rect 37046 2957 37106 8467
rect 66568 8192 66888 9216
rect 66568 8128 66576 8192
rect 66640 8128 66656 8192
rect 66720 8128 66736 8192
rect 66800 8128 66816 8192
rect 66880 8128 66888 8192
rect 66568 7104 66888 8128
rect 66568 7040 66576 7104
rect 66640 7040 66656 7104
rect 66720 7040 66736 7104
rect 66800 7040 66816 7104
rect 66880 7040 66888 7104
rect 66568 6016 66888 7040
rect 66568 5952 66576 6016
rect 66640 5952 66656 6016
rect 66720 5952 66736 6016
rect 66800 5952 66816 6016
rect 66880 5952 66888 6016
rect 66568 4928 66888 5952
rect 66568 4864 66576 4928
rect 66640 4864 66656 4928
rect 66720 4864 66736 4928
rect 66800 4864 66816 4928
rect 66880 4864 66888 4928
rect 66568 3840 66888 4864
rect 66568 3776 66576 3840
rect 66640 3776 66656 3840
rect 66720 3776 66736 3840
rect 66800 3776 66816 3840
rect 66880 3776 66888 3840
rect 37043 2956 37109 2957
rect 37043 2892 37044 2956
rect 37108 2892 37109 2956
rect 37043 2891 37109 2892
rect 36508 2144 36516 2208
rect 36580 2144 36596 2208
rect 36660 2144 36676 2208
rect 36740 2144 36756 2208
rect 36820 2144 36828 2208
rect 36508 2128 36828 2144
rect 66568 2752 66888 3776
rect 66568 2688 66576 2752
rect 66640 2688 66656 2752
rect 66720 2688 66736 2752
rect 66800 2688 66816 2752
rect 66880 2688 66888 2752
rect 66568 2128 66888 2688
rect 67228 37024 67548 37584
rect 67228 36960 67236 37024
rect 67300 36960 67316 37024
rect 67380 36960 67396 37024
rect 67460 36960 67476 37024
rect 67540 36960 67548 37024
rect 67228 35936 67548 36960
rect 67228 35872 67236 35936
rect 67300 35872 67316 35936
rect 67380 35872 67396 35936
rect 67460 35872 67476 35936
rect 67540 35872 67548 35936
rect 67228 34848 67548 35872
rect 67228 34784 67236 34848
rect 67300 34784 67316 34848
rect 67380 34784 67396 34848
rect 67460 34784 67476 34848
rect 67540 34784 67548 34848
rect 67228 33760 67548 34784
rect 67228 33696 67236 33760
rect 67300 33696 67316 33760
rect 67380 33696 67396 33760
rect 67460 33696 67476 33760
rect 67540 33696 67548 33760
rect 67228 32672 67548 33696
rect 67228 32608 67236 32672
rect 67300 32608 67316 32672
rect 67380 32608 67396 32672
rect 67460 32608 67476 32672
rect 67540 32608 67548 32672
rect 67228 31584 67548 32608
rect 67228 31520 67236 31584
rect 67300 31520 67316 31584
rect 67380 31520 67396 31584
rect 67460 31520 67476 31584
rect 67540 31520 67548 31584
rect 67228 30496 67548 31520
rect 67228 30432 67236 30496
rect 67300 30432 67316 30496
rect 67380 30432 67396 30496
rect 67460 30432 67476 30496
rect 67540 30432 67548 30496
rect 67228 29408 67548 30432
rect 67228 29344 67236 29408
rect 67300 29344 67316 29408
rect 67380 29344 67396 29408
rect 67460 29344 67476 29408
rect 67540 29344 67548 29408
rect 67228 28320 67548 29344
rect 67228 28256 67236 28320
rect 67300 28256 67316 28320
rect 67380 28256 67396 28320
rect 67460 28256 67476 28320
rect 67540 28256 67548 28320
rect 67228 27232 67548 28256
rect 67228 27168 67236 27232
rect 67300 27168 67316 27232
rect 67380 27168 67396 27232
rect 67460 27168 67476 27232
rect 67540 27168 67548 27232
rect 67228 26144 67548 27168
rect 67228 26080 67236 26144
rect 67300 26080 67316 26144
rect 67380 26080 67396 26144
rect 67460 26080 67476 26144
rect 67540 26080 67548 26144
rect 67228 25056 67548 26080
rect 67228 24992 67236 25056
rect 67300 24992 67316 25056
rect 67380 24992 67396 25056
rect 67460 24992 67476 25056
rect 67540 24992 67548 25056
rect 67228 23968 67548 24992
rect 67228 23904 67236 23968
rect 67300 23904 67316 23968
rect 67380 23904 67396 23968
rect 67460 23904 67476 23968
rect 67540 23904 67548 23968
rect 67228 22880 67548 23904
rect 67228 22816 67236 22880
rect 67300 22816 67316 22880
rect 67380 22816 67396 22880
rect 67460 22816 67476 22880
rect 67540 22816 67548 22880
rect 67228 21792 67548 22816
rect 67228 21728 67236 21792
rect 67300 21728 67316 21792
rect 67380 21728 67396 21792
rect 67460 21728 67476 21792
rect 67540 21728 67548 21792
rect 67228 20704 67548 21728
rect 67228 20640 67236 20704
rect 67300 20640 67316 20704
rect 67380 20640 67396 20704
rect 67460 20640 67476 20704
rect 67540 20640 67548 20704
rect 67228 19616 67548 20640
rect 67228 19552 67236 19616
rect 67300 19552 67316 19616
rect 67380 19552 67396 19616
rect 67460 19552 67476 19616
rect 67540 19552 67548 19616
rect 67228 18528 67548 19552
rect 67228 18464 67236 18528
rect 67300 18464 67316 18528
rect 67380 18464 67396 18528
rect 67460 18464 67476 18528
rect 67540 18464 67548 18528
rect 67228 17440 67548 18464
rect 67228 17376 67236 17440
rect 67300 17376 67316 17440
rect 67380 17376 67396 17440
rect 67460 17376 67476 17440
rect 67540 17376 67548 17440
rect 67228 16352 67548 17376
rect 67228 16288 67236 16352
rect 67300 16288 67316 16352
rect 67380 16288 67396 16352
rect 67460 16288 67476 16352
rect 67540 16288 67548 16352
rect 67228 15264 67548 16288
rect 67228 15200 67236 15264
rect 67300 15200 67316 15264
rect 67380 15200 67396 15264
rect 67460 15200 67476 15264
rect 67540 15200 67548 15264
rect 67228 14176 67548 15200
rect 67228 14112 67236 14176
rect 67300 14112 67316 14176
rect 67380 14112 67396 14176
rect 67460 14112 67476 14176
rect 67540 14112 67548 14176
rect 67228 13088 67548 14112
rect 67228 13024 67236 13088
rect 67300 13024 67316 13088
rect 67380 13024 67396 13088
rect 67460 13024 67476 13088
rect 67540 13024 67548 13088
rect 67228 12000 67548 13024
rect 67228 11936 67236 12000
rect 67300 11936 67316 12000
rect 67380 11936 67396 12000
rect 67460 11936 67476 12000
rect 67540 11936 67548 12000
rect 67228 10912 67548 11936
rect 67228 10848 67236 10912
rect 67300 10848 67316 10912
rect 67380 10848 67396 10912
rect 67460 10848 67476 10912
rect 67540 10848 67548 10912
rect 67228 9824 67548 10848
rect 67228 9760 67236 9824
rect 67300 9760 67316 9824
rect 67380 9760 67396 9824
rect 67460 9760 67476 9824
rect 67540 9760 67548 9824
rect 67228 8736 67548 9760
rect 67228 8672 67236 8736
rect 67300 8672 67316 8736
rect 67380 8672 67396 8736
rect 67460 8672 67476 8736
rect 67540 8672 67548 8736
rect 67228 7648 67548 8672
rect 67228 7584 67236 7648
rect 67300 7584 67316 7648
rect 67380 7584 67396 7648
rect 67460 7584 67476 7648
rect 67540 7584 67548 7648
rect 67228 6560 67548 7584
rect 67228 6496 67236 6560
rect 67300 6496 67316 6560
rect 67380 6496 67396 6560
rect 67460 6496 67476 6560
rect 67540 6496 67548 6560
rect 67228 5472 67548 6496
rect 67228 5408 67236 5472
rect 67300 5408 67316 5472
rect 67380 5408 67396 5472
rect 67460 5408 67476 5472
rect 67540 5408 67548 5472
rect 67228 4384 67548 5408
rect 67228 4320 67236 4384
rect 67300 4320 67316 4384
rect 67380 4320 67396 4384
rect 67460 4320 67476 4384
rect 67540 4320 67548 4384
rect 67228 3296 67548 4320
rect 67228 3232 67236 3296
rect 67300 3232 67316 3296
rect 67380 3232 67396 3296
rect 67460 3232 67476 3296
rect 67540 3232 67548 3296
rect 67228 2208 67548 3232
rect 67228 2144 67236 2208
rect 67300 2144 67316 2208
rect 67380 2144 67396 2208
rect 67460 2144 67476 2208
rect 67540 2144 67548 2208
rect 67228 2128 67548 2144
rect 33179 2075 33245 2076
rect 30235 1732 30301 1733
rect 30235 1668 30236 1732
rect 30300 1668 30301 1732
rect 30235 1667 30301 1668
rect 19195 1052 19261 1053
rect 19195 988 19196 1052
rect 19260 988 19261 1052
rect 19195 987 19261 988
<< via4 >>
rect 4758 8382 4994 8618
rect 6966 7702 7202 7938
rect 11750 10422 11986 10658
rect 15062 4452 15298 4538
rect 15062 4388 15148 4452
rect 15148 4388 15212 4452
rect 15212 4388 15298 4452
rect 15062 4302 15298 4388
rect 15982 3622 16218 3858
rect 19294 8532 19530 8618
rect 19294 8468 19380 8532
rect 19380 8468 19444 8532
rect 19444 8468 19530 8532
rect 19294 8382 19530 8468
rect 26102 10572 26338 10658
rect 26102 10508 26188 10572
rect 26188 10508 26252 10572
rect 26252 10508 26338 10572
rect 26102 10422 26338 10508
rect 25182 4302 25418 4538
rect 24630 2412 24866 2498
rect 24630 2348 24716 2412
rect 24716 2348 24780 2412
rect 24780 2348 24866 2412
rect 24630 2262 24866 2348
rect 30518 7852 30754 7938
rect 30518 7788 30604 7852
rect 30604 7788 30668 7852
rect 30668 7788 30754 7852
rect 30518 7702 30754 7788
rect 33646 2262 33882 2498
rect 73942 3772 74178 3858
rect 73942 3708 74028 3772
rect 74028 3708 74092 3772
rect 74092 3708 74178 3772
rect 73942 3622 74178 3708
<< metal5 >>
rect 11708 10658 26380 10700
rect 11708 10422 11750 10658
rect 11986 10422 26102 10658
rect 26338 10422 26380 10658
rect 11708 10380 26380 10422
rect 4716 8618 19572 8660
rect 4716 8382 4758 8618
rect 4994 8382 19294 8618
rect 19530 8382 19572 8618
rect 4716 8340 19572 8382
rect 6924 7938 30796 7980
rect 6924 7702 6966 7938
rect 7202 7702 30518 7938
rect 30754 7702 30796 7938
rect 6924 7660 30796 7702
rect 15020 4538 25460 4580
rect 15020 4302 15062 4538
rect 15298 4302 25182 4538
rect 25418 4302 25460 4538
rect 15020 4260 25460 4302
rect 15940 3858 74220 3900
rect 15940 3622 15982 3858
rect 16218 3622 73942 3858
rect 74178 3622 74220 3858
rect 15940 3580 74220 3622
rect 24588 2498 33924 2540
rect 24588 2262 24630 2498
rect 24866 2262 33646 2498
rect 33882 2262 33924 2498
rect 24588 2220 33924 2262
use sky130_fd_sc_hd__inv_2  _099_
timestamp 25201
transform 1 0 21252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 25201
transform 1 0 32568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 25201
transform -1 0 32936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 25201
transform -1 0 39008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 25201
transform -1 0 11960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _104_
timestamp 25201
transform -1 0 43884 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _105_
timestamp 25201
transform -1 0 27784 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _106_
timestamp 25201
transform 1 0 28152 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _107_
timestamp 25201
transform 1 0 17204 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_4  _108_
timestamp 25201
transform -1 0 39744 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_4  _109_
timestamp 25201
transform 1 0 12420 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _110_
timestamp 25201
transform 1 0 20424 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 25201
transform 1 0 12420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _112_
timestamp 25201
transform -1 0 19780 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _113_
timestamp 25201
transform 1 0 17572 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _114_
timestamp 25201
transform 1 0 21528 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _115_
timestamp 25201
transform -1 0 22632 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _116_
timestamp 25201
transform 1 0 12512 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _117_
timestamp 25201
transform 1 0 22724 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _118_
timestamp 25201
transform -1 0 23276 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _119_
timestamp 25201
transform 1 0 29256 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _120_
timestamp 25201
transform 1 0 30544 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _121_
timestamp 25201
transform -1 0 32384 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _122_
timestamp 25201
transform -1 0 34776 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _123_
timestamp 25201
transform -1 0 30912 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _124_
timestamp 25201
transform 1 0 35604 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _125_
timestamp 25201
transform 1 0 40112 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _126_
timestamp 25201
transform -1 0 43148 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _127_
timestamp 25201
transform 1 0 33028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _128_
timestamp 25201
transform -1 0 43240 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _129_
timestamp 25201
transform 1 0 15180 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_2  _130_
timestamp 25201
transform -1 0 11960 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _131_
timestamp 25201
transform -1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _132_
timestamp 25201
transform -1 0 19504 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _133_
timestamp 25201
transform 1 0 20792 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _134_
timestamp 25201
transform -1 0 24656 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _135_
timestamp 25201
transform 1 0 19596 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _136_
timestamp 25201
transform -1 0 27508 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 25201
transform -1 0 35880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _138_
timestamp 25201
transform -1 0 20424 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _139_
timestamp 25201
transform 1 0 21620 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _140_
timestamp 25201
transform -1 0 15640 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _141_
timestamp 25201
transform 1 0 21344 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _142_
timestamp 25201
transform 1 0 20516 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _143_
timestamp 25201
transform 1 0 17572 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _144_
timestamp 25201
transform -1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _145_
timestamp 25201
transform -1 0 21160 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _146_
timestamp 25201
transform 1 0 24196 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _147_
timestamp 25201
transform 1 0 20424 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _148_
timestamp 25201
transform 1 0 20148 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _149_
timestamp 25201
transform 1 0 21160 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _150_
timestamp 25201
transform -1 0 25944 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _151_
timestamp 25201
transform 1 0 22264 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _152_
timestamp 25201
transform -1 0 26772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _153_
timestamp 25201
transform -1 0 25024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _154_
timestamp 25201
transform 1 0 24564 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _155_
timestamp 25201
transform -1 0 24472 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _156_
timestamp 25201
transform 1 0 26036 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _157_
timestamp 25201
transform -1 0 24196 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _158_
timestamp 25201
transform -1 0 25668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _159_
timestamp 25201
transform 1 0 22172 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _160_
timestamp 25201
transform 1 0 27876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _161_
timestamp 25201
transform 1 0 26864 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _162_
timestamp 25201
transform -1 0 28152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _163_
timestamp 25201
transform -1 0 22632 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _164_
timestamp 25201
transform 1 0 25300 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _165_
timestamp 25201
transform 1 0 21988 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _166_
timestamp 25201
transform 1 0 29532 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _167_
timestamp 25201
transform 1 0 28060 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _168_
timestamp 25201
transform 1 0 33028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _169_
timestamp 25201
transform 1 0 30452 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _170_
timestamp 25201
transform -1 0 29900 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _171_
timestamp 25201
transform 1 0 31004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _172_
timestamp 25201
transform -1 0 27784 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _173_
timestamp 25201
transform -1 0 32200 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _174_
timestamp 25201
transform 1 0 33028 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _175_
timestamp 25201
transform 1 0 32200 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _176_
timestamp 25201
transform -1 0 31096 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _177_
timestamp 25201
transform 1 0 33028 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _178_
timestamp 25201
transform 1 0 35604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _179_
timestamp 25201
transform 1 0 34868 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _180_
timestamp 25201
transform 1 0 27140 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _181_
timestamp 25201
transform 1 0 33856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _182_
timestamp 25201
transform 1 0 34132 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _183_
timestamp 25201
transform -1 0 34040 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _184_
timestamp 25201
transform -1 0 42228 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 25201
transform 1 0 36984 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _186_
timestamp 25201
transform -1 0 32200 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _187_
timestamp 25201
transform 1 0 27876 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _188_
timestamp 25201
transform -1 0 38456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _189_
timestamp 25201
transform -1 0 34776 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _190_
timestamp 25201
transform 1 0 30452 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _191_
timestamp 25201
transform -1 0 32108 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _192_
timestamp 25201
transform -1 0 34684 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _193_
timestamp 25201
transform -1 0 25944 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _194_
timestamp 25201
transform -1 0 35512 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _195_
timestamp 25201
transform 1 0 40204 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _196_
timestamp 25201
transform 1 0 34040 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _197_
timestamp 25201
transform -1 0 36616 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _198_
timestamp 25201
transform 1 0 11224 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _199_
timestamp 25201
transform 1 0 12420 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _200_
timestamp 25201
transform 1 0 14996 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _201_
timestamp 25201
transform 1 0 17572 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _202_
timestamp 25201
transform 1 0 19504 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _203_
timestamp 25201
transform 1 0 20884 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _204_
timestamp 25201
transform 1 0 22908 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp 25201
transform 1 0 25668 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 25201
transform 1 0 27876 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _207_
timestamp 25201
transform 1 0 29900 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 25201
transform 1 0 31372 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 25201
transform 1 0 33028 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 25201
transform 1 0 34684 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _211_
timestamp 25201
transform -1 0 36616 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 25201
transform 1 0 40756 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 25201
transform -1 0 41400 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 25201
transform 1 0 44804 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _215_
timestamp 25201
transform -1 0 44896 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _216_
timestamp 25201
transform 1 0 14904 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _217_
timestamp 25201
transform 1 0 18952 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _218_
timestamp 25201
transform 1 0 20148 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _219_
timestamp 25201
transform 1 0 22080 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _220_
timestamp 25201
transform 1 0 24012 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _221_
timestamp 25201
transform 1 0 24288 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _222_
timestamp 25201
transform 1 0 25024 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _223_
timestamp 25201
transform 1 0 26680 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _224_
timestamp 25201
transform 1 0 29624 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _225_
timestamp 25201
transform 1 0 29716 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _226_
timestamp 25201
transform 1 0 30544 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _227_
timestamp 25201
transform -1 0 34224 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _228_
timestamp 25201
transform 1 0 34776 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _229_
timestamp 25201
transform -1 0 38088 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _230_
timestamp 25201
transform 1 0 37812 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _231_
timestamp 25201
transform 1 0 38180 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _232_
timestamp 25201
transform 1 0 33028 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _233_
timestamp 25201
transform 1 0 37352 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _234_
timestamp 25201
transform 1 0 10488 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _235_
timestamp 25201
transform 1 0 11960 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _236_
timestamp 25201
transform 1 0 13064 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _237_
timestamp 25201
transform -1 0 18216 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _238_
timestamp 25201
transform 1 0 18308 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _239_
timestamp 25201
transform 1 0 20148 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _240_
timestamp 25201
transform 1 0 23184 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _241_
timestamp 25201
transform 1 0 25300 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _242_
timestamp 25201
transform 1 0 26680 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _243_
timestamp 25201
transform -1 0 30360 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _244_
timestamp 25201
transform 1 0 30912 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _245_
timestamp 25201
transform 1 0 32384 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _246_
timestamp 25201
transform -1 0 35972 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _247_
timestamp 25201
transform -1 0 37996 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _248_
timestamp 25201
transform 1 0 38640 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _249_
timestamp 25201
transform -1 0 42044 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _250_
timestamp 25201
transform 1 0 41400 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _251_
timestamp 25201
transform 1 0 42228 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _258_
timestamp 25201
transform 1 0 47840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _259_
timestamp 25201
transform 1 0 51060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _260_
timestamp 25201
transform -1 0 53912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _261_
timestamp 25201
transform 1 0 57132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _262_
timestamp 25201
transform 1 0 60720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _263_
timestamp 25201
transform 1 0 64492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _264_
timestamp 25201
transform 1 0 66976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _265_
timestamp 25201
transform -1 0 69368 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _266_
timestamp 25201
transform 1 0 70656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _267_
timestamp 25201
transform 1 0 74244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _268_
timestamp 25201
transform 1 0 58420 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _269_
timestamp 25201
transform 1 0 55384 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _270_
timestamp 25201
transform 1 0 51704 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _271_
timestamp 25201
transform 1 0 48024 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _272_
timestamp 25201
transform 1 0 44344 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _273_
timestamp 25201
transform 1 0 40664 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _274_
timestamp 25201
transform -1 0 37260 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _275_
timestamp 25201
transform -1 0 34040 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _276_
timestamp 25201
transform 1 0 29624 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _277_
timestamp 25201
transform 1 0 25944 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _278_
timestamp 25201
transform 1 0 22264 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _279_
timestamp 25201
transform -1 0 19320 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _280_
timestamp 25201
transform 1 0 14904 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _281_
timestamp 25201
transform -1 0 12144 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _282_
timestamp 25201
transform 1 0 7544 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_116
timestamp 25201
transform -1 0 50968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_117
timestamp 25201
transform -1 0 55752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_118
timestamp 25201
transform -1 0 59616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_119
timestamp 25201
transform -1 0 63480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_120
timestamp 25201
transform -1 0 73416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_121
timestamp 25201
transform -1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 25201
transform 1 0 21252 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 25201
transform -1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 25201
transform -1 0 33304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 25201
transform -1 0 7544 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 25201
transform 1 0 9936 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 25201
transform -1 0 25484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 25201
transform -1 0 19872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 25201
transform -1 0 35144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 25201
transform -1 0 28060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 25201
transform 1 0 23276 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 25201
transform 1 0 24012 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 25201
transform -1 0 36156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 25201
transform -1 0 13432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 25201
transform -1 0 28796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 25201
transform 1 0 27968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 25201
transform -1 0 26128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 25201
transform 1 0 26496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 25201
transform 1 0 27324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 25201
transform -1 0 18584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 25201
transform 1 0 16192 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 25201
transform -1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 25201
transform -1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 25201
transform 1 0 28888 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 25201
transform 1 0 26036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 25201
transform 1 0 30544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 25201
transform 1 0 27876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 25201
transform -1 0 19504 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 25201
transform -1 0 15180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 25201
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 25201
transform -1 0 12328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 25201
transform 1 0 15916 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 25201
transform 1 0 28520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_HCLK
timestamp 25201
transform 1 0 26864 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_HCLK
timestamp 25201
transform -1 0 19504 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_HCLK
timestamp 25201
transform 1 0 22724 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_HCLK
timestamp 25201
transform 1 0 36892 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_HCLK
timestamp 25201
transform 1 0 32292 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_2  clkload0
timestamp 25201
transform -1 0 15456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp 25201
transform -1 0 18216 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload2
timestamp 25201
transform -1 0 31004 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout97
timestamp 25201
transform -1 0 23552 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout98
timestamp 25201
transform 1 0 31740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout99
timestamp 25201
transform -1 0 23092 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout100
timestamp 25201
transform -1 0 20700 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout101
timestamp 25201
transform -1 0 37812 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout102
timestamp 25201
transform 1 0 15824 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout105
timestamp 25201
transform -1 0 20056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout106
timestamp 25201
transform 1 0 28520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout107
timestamp 25201
transform -1 0 11868 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout108
timestamp 25201
transform 1 0 33396 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout109
timestamp 25201
transform -1 0 10120 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp 25201
transform 1 0 14904 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout111
timestamp 25201
transform -1 0 29256 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout112
timestamp 25201
transform 1 0 12512 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout113
timestamp 25201
transform 1 0 9936 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout114
timestamp 25201
transform -1 0 10488 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout115
timestamp 25201
transform 1 0 31096 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636993656
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 25201
transform 1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 25201
transform 1 0 7268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 25201
transform 1 0 9844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109
timestamp 25201
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_309
timestamp 25201
transform 1 0 30452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_337
timestamp 25201
transform 1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_410
timestamp 25201
transform 1 0 39744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 25201
transform 1 0 45632 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_533
timestamp 25201
transform 1 0 51060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_555
timestamp 25201
transform 1 0 53084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 25201
transform 1 0 53452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_577
timestamp 25201
transform 1 0 55108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_584
timestamp 25201
transform 1 0 55752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_589
timestamp 25201
transform 1 0 56212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_597
timestamp 25201
transform 1 0 56948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_633
timestamp 25201
transform 1 0 60260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 25201
transform 1 0 60996 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_661
timestamp 25201
transform 1 0 62836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_668
timestamp 25201
transform 1 0 63480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_673
timestamp 25201
transform 1 0 63940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_681
timestamp 25201
transform 1 0 64676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_701
timestamp 25201
transform 1 0 66516 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_723
timestamp 25201
transform 1 0 68540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_727
timestamp 25201
transform 1 0 68908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_745
timestamp 25201
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_749
timestamp 25201
transform 1 0 70932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_755
timestamp 25201
transform 1 0 71484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_785
timestamp 25201
transform 1 0 74244 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_807
timestamp 25201
transform 1 0 76268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_811
timestamp 25201
transform 1 0 76636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_821
timestamp 25201
transform 1 0 77556 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636993656
transform 1 0 2300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 25201
transform 1 0 3404 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_23
timestamp 25201
transform 1 0 4140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 25201
transform 1 0 7268 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 25201
transform 1 0 12420 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 25201
transform 1 0 32752 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 25201
transform 1 0 37996 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_396
timestamp 25201
transform 1 0 38456 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_418
timestamp 25201
transform 1 0 40480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 25201
transform 1 0 48484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_530
timestamp 25201
transform 1 0 50784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_564
timestamp 25201
transform 1 0 53912 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_589
timestamp 25201
transform 1 0 56212 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_597
timestamp 25201
transform 1 0 56948 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_610
timestamp 25201
transform 1 0 58144 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_617
timestamp 25201
transform 1 0 58788 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_626
timestamp 1636993656
transform 1 0 59616 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 25201
transform 1 0 63204 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 25201
transform 1 0 63756 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_673
timestamp 25201
transform 1 0 63940 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_709
timestamp 25201
transform 1 0 67252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_732
timestamp 25201
transform 1 0 69368 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_757
timestamp 25201
transform 1 0 71668 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_774
timestamp 25201
transform 1 0 73232 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_782
timestamp 25201
transform 1 0 73968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_820
timestamp 25201
transform 1 0 77464 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636993656
transform 1 0 2300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636993656
transform 1 0 3404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 25201
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 25201
transform 1 0 4968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 25201
transform 1 0 9844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_104
timestamp 25201
transform 1 0 11592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_128
timestamp 25201
transform 1 0 13800 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_215
timestamp 25201
transform 1 0 21804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_387
timestamp 25201
transform 1 0 37628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 25201
transform 1 0 45632 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_480
timestamp 25201
transform 1 0 46184 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_497
timestamp 25201
transform 1 0 47748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_529
timestamp 25201
transform 1 0 50692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_533
timestamp 25201
transform 1 0 51060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_539
timestamp 25201
transform 1 0 51612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_556
timestamp 25201
transform 1 0 53176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_560
timestamp 25201
transform 1 0 53544 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_577
timestamp 25201
transform 1 0 55108 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_585
timestamp 25201
transform 1 0 55844 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636993656
transform 1 0 56212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_601
timestamp 25201
transform 1 0 57316 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_618
timestamp 1636993656
transform 1 0 58880 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_630
timestamp 1636993656
transform 1 0 59984 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_642
timestamp 25201
transform 1 0 61088 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_661
timestamp 1636993656
transform 1 0 62836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_673
timestamp 1636993656
transform 1 0 63940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_685
timestamp 25201
transform 1 0 65044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_694
timestamp 25201
transform 1 0 65872 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_701
timestamp 25201
transform 1 0 66516 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_707
timestamp 25201
transform 1 0 67068 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_724
timestamp 25201
transform 1 0 68632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_728
timestamp 25201
transform 1 0 69000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_745
timestamp 25201
transform 1 0 70564 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_753
timestamp 25201
transform 1 0 71300 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_773
timestamp 1636993656
transform 1 0 73140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_785
timestamp 25201
transform 1 0 74244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_813
timestamp 25201
transform 1 0 76820 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636993656
transform 1 0 2300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636993656
transform 1 0 3404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636993656
transform 1 0 4508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_39
timestamp 25201
transform 1 0 5612 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 25201
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 25201
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_60
timestamp 25201
transform 1 0 7544 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp 25201
transform 1 0 17572 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_199
timestamp 25201
transform 1 0 20332 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_225
timestamp 25201
transform 1 0 22724 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_269
timestamp 25201
transform 1 0 26772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_281
timestamp 25201
transform 1 0 27876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_364
timestamp 25201
transform 1 0 35512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_396
timestamp 25201
transform 1 0 38456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_413
timestamp 25201
transform 1 0 40020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_443
timestamp 25201
transform 1 0 42780 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 25201
transform 1 0 43148 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_449
timestamp 25201
transform 1 0 43332 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_501
timestamp 25201
transform 1 0 48116 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636993656
transform 1 0 50692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_541
timestamp 25201
transform 1 0 51796 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_555
timestamp 25201
transform 1 0 53084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 25201
transform 1 0 53452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636993656
transform 1 0 53636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636993656
transform 1 0 54740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636993656
transform 1 0 55844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636993656
transform 1 0 56948 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 25201
transform 1 0 58052 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 25201
transform 1 0 58604 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636993656
transform 1 0 58788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636993656
transform 1 0 59892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636993656
transform 1 0 60996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636993656
transform 1 0 62100 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 25201
transform 1 0 63204 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 25201
transform 1 0 63756 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636993656
transform 1 0 63940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_685
timestamp 25201
transform 1 0 65044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_689
timestamp 25201
transform 1 0 65412 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_698
timestamp 1636993656
transform 1 0 66240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_710
timestamp 25201
transform 1 0 67344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_720
timestamp 25201
transform 1 0 68264 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636993656
transform 1 0 69092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636993656
transform 1 0 70196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_753
timestamp 25201
transform 1 0 71300 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_762
timestamp 1636993656
transform 1 0 72128 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_774
timestamp 25201
transform 1 0 73232 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_782
timestamp 25201
transform 1 0 73968 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_785
timestamp 25201
transform 1 0 74244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_789
timestamp 25201
transform 1 0 74612 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636993656
transform 1 0 2300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636993656
transform 1 0 3404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 25201
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636993656
transform 1 0 4692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_41
timestamp 25201
transform 1 0 5796 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_49
timestamp 25201
transform 1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 25201
transform 1 0 9844 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_262
timestamp 25201
transform 1 0 26128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_290
timestamp 25201
transform 1 0 28704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 25201
transform 1 0 30452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_328
timestamp 25201
transform 1 0 32200 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_365
timestamp 25201
transform 1 0 35604 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_421
timestamp 25201
transform 1 0 40756 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_433
timestamp 25201
transform 1 0 41860 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_517
timestamp 1636993656
transform 1 0 49588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_529
timestamp 25201
transform 1 0 50692 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636993656
transform 1 0 51060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636993656
transform 1 0 52164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1636993656
transform 1 0 53268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1636993656
transform 1 0 54372 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 25201
transform 1 0 55476 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 25201
transform 1 0 56028 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636993656
transform 1 0 56212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636993656
transform 1 0 57316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1636993656
transform 1 0 58420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1636993656
transform 1 0 59524 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 25201
transform 1 0 60628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 25201
transform 1 0 61180 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636993656
transform 1 0 61364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636993656
transform 1 0 62468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1636993656
transform 1 0 63572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1636993656
transform 1 0 64676 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 25201
transform 1 0 65780 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 25201
transform 1 0 66332 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636993656
transform 1 0 66516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636993656
transform 1 0 67620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1636993656
transform 1 0 68724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1636993656
transform 1 0 69828 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 25201
transform 1 0 70932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 25201
transform 1 0 71484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636993656
transform 1 0 71668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636993656
transform 1 0 72772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1636993656
transform 1 0 73876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1636993656
transform 1 0 74980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 25201
transform 1 0 76084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 25201
transform 1 0 76636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_813
timestamp 25201
transform 1 0 76820 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636993656
transform 1 0 2300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636993656
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636993656
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636993656
transform 1 0 5612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 25201
transform 1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 25201
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 25201
transform 1 0 7268 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp 25201
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 25201
transform 1 0 12420 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_283
timestamp 25201
transform 1 0 28060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_308
timestamp 25201
transform 1 0 30360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_337
timestamp 25201
transform 1 0 33028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_389
timestamp 25201
transform 1 0 37812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 25201
transform 1 0 43148 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_489
timestamp 1636993656
transform 1 0 47012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_501
timestamp 25201
transform 1 0 48116 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1636993656
transform 1 0 48484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1636993656
transform 1 0 49588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1636993656
transform 1 0 50692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1636993656
transform 1 0 51796 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 25201
transform 1 0 52900 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 25201
transform 1 0 53452 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1636993656
transform 1 0 53636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1636993656
transform 1 0 54740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1636993656
transform 1 0 55844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1636993656
transform 1 0 56948 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 25201
transform 1 0 58052 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 25201
transform 1 0 58604 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1636993656
transform 1 0 58788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1636993656
transform 1 0 59892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1636993656
transform 1 0 60996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1636993656
transform 1 0 62100 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 25201
transform 1 0 63204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 25201
transform 1 0 63756 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1636993656
transform 1 0 63940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1636993656
transform 1 0 65044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1636993656
transform 1 0 66148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1636993656
transform 1 0 67252 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 25201
transform 1 0 68356 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 25201
transform 1 0 68908 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1636993656
transform 1 0 69092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1636993656
transform 1 0 70196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1636993656
transform 1 0 71300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1636993656
transform 1 0 72404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 25201
transform 1 0 73508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 25201
transform 1 0 74060 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1636993656
transform 1 0 74244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1636993656
transform 1 0 75348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_809
timestamp 25201
transform 1 0 76452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_813
timestamp 25201
transform 1 0 76820 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636993656
transform 1 0 2300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636993656
transform 1 0 3404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 25201
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636993656
transform 1 0 4692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636993656
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636993656
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 25201
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_73
timestamp 25201
transform 1 0 8740 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 25201
transform 1 0 9844 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 25201
transform 1 0 10304 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_153
timestamp 25201
transform 1 0 16100 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_253
timestamp 25201
transform 1 0 25300 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_290
timestamp 25201
transform 1 0 28704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_318
timestamp 25201
transform 1 0 31280 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_328
timestamp 25201
transform 1 0 32200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp 25201
transform 1 0 40480 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_471
timestamp 25201
transform 1 0 45356 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 25201
transform 1 0 45724 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_485
timestamp 1636993656
transform 1 0 46644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_497
timestamp 1636993656
transform 1 0 47748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_509
timestamp 1636993656
transform 1 0 48852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_521
timestamp 25201
transform 1 0 49956 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_529
timestamp 25201
transform 1 0 50692 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1636993656
transform 1 0 51060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1636993656
transform 1 0 52164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1636993656
transform 1 0 53268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1636993656
transform 1 0 54372 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 25201
transform 1 0 55476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 25201
transform 1 0 56028 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1636993656
transform 1 0 56212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1636993656
transform 1 0 57316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1636993656
transform 1 0 58420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1636993656
transform 1 0 59524 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 25201
transform 1 0 60628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 25201
transform 1 0 61180 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1636993656
transform 1 0 61364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1636993656
transform 1 0 62468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1636993656
transform 1 0 63572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1636993656
transform 1 0 64676 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 25201
transform 1 0 65780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 25201
transform 1 0 66332 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1636993656
transform 1 0 66516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1636993656
transform 1 0 67620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1636993656
transform 1 0 68724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1636993656
transform 1 0 69828 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 25201
transform 1 0 70932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 25201
transform 1 0 71484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1636993656
transform 1 0 71668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1636993656
transform 1 0 72772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1636993656
transform 1 0 73876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1636993656
transform 1 0 74980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 25201
transform 1 0 76084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 25201
transform 1 0 76636 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_813
timestamp 25201
transform 1 0 76820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_821
timestamp 25201
transform 1 0 77556 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636993656
transform 1 0 2300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636993656
transform 1 0 3404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636993656
transform 1 0 4508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636993656
transform 1 0 5612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 25201
transform 1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 25201
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636993656
transform 1 0 7268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636993656
transform 1 0 8372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_102
timestamp 25201
transform 1 0 11408 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 25201
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 25201
transform 1 0 17572 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_268
timestamp 25201
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 25201
transform 1 0 27692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp 25201
transform 1 0 27876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 25201
transform 1 0 32844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_416
timestamp 25201
transform 1 0 40296 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1636993656
transform 1 0 43332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1636993656
transform 1 0 44436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1636993656
transform 1 0 45540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1636993656
transform 1 0 46644 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 25201
transform 1 0 47748 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 25201
transform 1 0 48300 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1636993656
transform 1 0 48484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1636993656
transform 1 0 49588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1636993656
transform 1 0 50692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1636993656
transform 1 0 51796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 25201
transform 1 0 52900 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 25201
transform 1 0 53452 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1636993656
transform 1 0 53636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1636993656
transform 1 0 54740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1636993656
transform 1 0 55844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1636993656
transform 1 0 56948 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 25201
transform 1 0 58052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 25201
transform 1 0 58604 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1636993656
transform 1 0 58788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1636993656
transform 1 0 59892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1636993656
transform 1 0 60996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1636993656
transform 1 0 62100 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 25201
transform 1 0 63204 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 25201
transform 1 0 63756 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1636993656
transform 1 0 63940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1636993656
transform 1 0 65044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1636993656
transform 1 0 66148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1636993656
transform 1 0 67252 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 25201
transform 1 0 68356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 25201
transform 1 0 68908 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1636993656
transform 1 0 69092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1636993656
transform 1 0 70196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1636993656
transform 1 0 71300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1636993656
transform 1 0 72404 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 25201
transform 1 0 73508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 25201
transform 1 0 74060 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1636993656
transform 1 0 74244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1636993656
transform 1 0 75348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1636993656
transform 1 0 76452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_821
timestamp 25201
transform 1 0 77556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636993656
transform 1 0 2300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636993656
transform 1 0 3404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 25201
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636993656
transform 1 0 4692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636993656
transform 1 0 5796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636993656
transform 1 0 6900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636993656
transform 1 0 8004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 25201
transform 1 0 9108 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 25201
transform 1 0 9660 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 25201
transform 1 0 9844 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 25201
transform 1 0 10396 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_108
timestamp 25201
transform 1 0 11960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 25201
transform 1 0 24932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_291
timestamp 25201
transform 1 0 28796 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1636993656
transform 1 0 42964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1636993656
transform 1 0 44068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 25201
transform 1 0 45172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 25201
transform 1 0 45724 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1636993656
transform 1 0 45908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1636993656
transform 1 0 47012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1636993656
transform 1 0 48116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1636993656
transform 1 0 49220 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 25201
transform 1 0 50324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 25201
transform 1 0 50876 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1636993656
transform 1 0 51060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1636993656
transform 1 0 52164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1636993656
transform 1 0 53268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1636993656
transform 1 0 54372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 25201
transform 1 0 55476 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 25201
transform 1 0 56028 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1636993656
transform 1 0 56212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1636993656
transform 1 0 57316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1636993656
transform 1 0 58420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1636993656
transform 1 0 59524 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 25201
transform 1 0 60628 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 25201
transform 1 0 61180 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1636993656
transform 1 0 61364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1636993656
transform 1 0 62468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1636993656
transform 1 0 63572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1636993656
transform 1 0 64676 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 25201
transform 1 0 65780 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 25201
transform 1 0 66332 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1636993656
transform 1 0 66516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1636993656
transform 1 0 67620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1636993656
transform 1 0 68724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1636993656
transform 1 0 69828 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 25201
transform 1 0 70932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 25201
transform 1 0 71484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1636993656
transform 1 0 71668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1636993656
transform 1 0 72772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1636993656
transform 1 0 73876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1636993656
transform 1 0 74980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 25201
transform 1 0 76084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 25201
transform 1 0 76636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_813
timestamp 25201
transform 1 0 76820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_821
timestamp 25201
transform 1 0 77556 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636993656
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636993656
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636993656
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636993656
transform 1 0 5612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 25201
transform 1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 25201
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636993656
transform 1 0 7268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636993656
transform 1 0 8372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636993656
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636993656
transform 1 0 10580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 25201
transform 1 0 11684 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 25201
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 25201
transform 1 0 12420 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_117
timestamp 1636993656
transform 1 0 12788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 25201
transform 1 0 13892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_241
timestamp 25201
transform 1 0 24196 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_281
timestamp 25201
transform 1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_300
timestamp 25201
transform 1 0 29624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp 25201
transform 1 0 33028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_364
timestamp 25201
transform 1 0 35512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_383
timestamp 25201
transform 1 0 37260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_401
timestamp 25201
transform 1 0 38916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_411
timestamp 25201
transform 1 0 39836 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1636993656
transform 1 0 41492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 25201
transform 1 0 42596 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 25201
transform 1 0 43148 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1636993656
transform 1 0 43332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1636993656
transform 1 0 44436 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1636993656
transform 1 0 45540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1636993656
transform 1 0 46644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 25201
transform 1 0 47748 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 25201
transform 1 0 48300 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1636993656
transform 1 0 48484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1636993656
transform 1 0 49588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1636993656
transform 1 0 50692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1636993656
transform 1 0 51796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 25201
transform 1 0 52900 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 25201
transform 1 0 53452 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1636993656
transform 1 0 53636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1636993656
transform 1 0 54740 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1636993656
transform 1 0 55844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1636993656
transform 1 0 56948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 25201
transform 1 0 58052 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 25201
transform 1 0 58604 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1636993656
transform 1 0 58788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1636993656
transform 1 0 59892 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1636993656
transform 1 0 60996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1636993656
transform 1 0 62100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 25201
transform 1 0 63204 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 25201
transform 1 0 63756 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1636993656
transform 1 0 63940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1636993656
transform 1 0 65044 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1636993656
transform 1 0 66148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1636993656
transform 1 0 67252 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 25201
transform 1 0 68356 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 25201
transform 1 0 68908 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1636993656
transform 1 0 69092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1636993656
transform 1 0 70196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_753
timestamp 1636993656
transform 1 0 71300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_765
timestamp 1636993656
transform 1 0 72404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 25201
transform 1 0 73508 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 25201
transform 1 0 74060 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1636993656
transform 1 0 74244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1636993656
transform 1 0 75348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_809
timestamp 1636993656
transform 1 0 76452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_821
timestamp 25201
transform 1 0 77556 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636993656
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636993656
transform 1 0 3404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 25201
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636993656
transform 1 0 4692 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636993656
transform 1 0 5796 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636993656
transform 1 0 6900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1636993656
transform 1 0 8004 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 25201
transform 1 0 9108 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 25201
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636993656
transform 1 0 9844 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636993656
transform 1 0 10948 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636993656
transform 1 0 12052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636993656
transform 1 0 13156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_133
timestamp 25201
transform 1 0 14260 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 25201
transform 1 0 14996 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_166
timestamp 25201
transform 1 0 17296 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 25201
transform 1 0 19872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 25201
transform 1 0 20148 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_216
timestamp 25201
transform 1 0 21896 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 25201
transform 1 0 25300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_368
timestamp 25201
transform 1 0 35880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_400
timestamp 25201
transform 1 0 38824 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1636993656
transform 1 0 40756 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1636993656
transform 1 0 41860 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1636993656
transform 1 0 42964 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1636993656
transform 1 0 44068 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 25201
transform 1 0 45172 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 25201
transform 1 0 45724 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1636993656
transform 1 0 45908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1636993656
transform 1 0 47012 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1636993656
transform 1 0 48116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1636993656
transform 1 0 49220 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 25201
transform 1 0 50324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 25201
transform 1 0 50876 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1636993656
transform 1 0 51060 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1636993656
transform 1 0 52164 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1636993656
transform 1 0 53268 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1636993656
transform 1 0 54372 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 25201
transform 1 0 55476 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 25201
transform 1 0 56028 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1636993656
transform 1 0 56212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1636993656
transform 1 0 57316 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1636993656
transform 1 0 58420 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1636993656
transform 1 0 59524 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 25201
transform 1 0 60628 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 25201
transform 1 0 61180 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1636993656
transform 1 0 61364 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1636993656
transform 1 0 62468 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1636993656
transform 1 0 63572 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1636993656
transform 1 0 64676 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 25201
transform 1 0 65780 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 25201
transform 1 0 66332 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1636993656
transform 1 0 66516 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1636993656
transform 1 0 67620 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_725
timestamp 1636993656
transform 1 0 68724 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_737
timestamp 1636993656
transform 1 0 69828 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 25201
transform 1 0 70932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 25201
transform 1 0 71484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1636993656
transform 1 0 71668 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_769
timestamp 1636993656
transform 1 0 72772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_781
timestamp 1636993656
transform 1 0 73876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_793
timestamp 1636993656
transform 1 0 74980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 25201
transform 1 0 76084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 25201
transform 1 0 76636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_813
timestamp 25201
transform 1 0 76820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_821
timestamp 25201
transform 1 0 77556 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636993656
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636993656
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636993656
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636993656
transform 1 0 5612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 25201
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 25201
transform 1 0 7084 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636993656
transform 1 0 7268 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1636993656
transform 1 0 8372 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1636993656
transform 1 0 9476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1636993656
transform 1 0 10580 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 25201
transform 1 0 11684 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 25201
transform 1 0 12236 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1636993656
transform 1 0 12420 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1636993656
transform 1 0 13524 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_137
timestamp 25201
transform 1 0 14628 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_145
timestamp 25201
transform 1 0 15364 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_154
timestamp 25201
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_158
timestamp 25201
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 25201
transform 1 0 17388 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 25201
transform 1 0 17572 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_190
timestamp 25201
transform 1 0 19504 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 25201
transform 1 0 22724 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_236
timestamp 25201
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_262
timestamp 25201
transform 1 0 26128 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_327
timestamp 25201
transform 1 0 32108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_340
timestamp 25201
transform 1 0 33304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_387
timestamp 25201
transform 1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 25201
transform 1 0 37996 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_401
timestamp 25201
transform 1 0 38916 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_423
timestamp 1636993656
transform 1 0 40940 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_435
timestamp 1636993656
transform 1 0 42044 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 25201
transform 1 0 43148 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1636993656
transform 1 0 43332 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1636993656
transform 1 0 44436 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1636993656
transform 1 0 45540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1636993656
transform 1 0 46644 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 25201
transform 1 0 47748 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 25201
transform 1 0 48300 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1636993656
transform 1 0 48484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1636993656
transform 1 0 49588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1636993656
transform 1 0 50692 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1636993656
transform 1 0 51796 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 25201
transform 1 0 52900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 25201
transform 1 0 53452 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1636993656
transform 1 0 53636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1636993656
transform 1 0 54740 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1636993656
transform 1 0 55844 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1636993656
transform 1 0 56948 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 25201
transform 1 0 58052 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 25201
transform 1 0 58604 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1636993656
transform 1 0 58788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1636993656
transform 1 0 59892 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1636993656
transform 1 0 60996 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1636993656
transform 1 0 62100 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 25201
transform 1 0 63204 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 25201
transform 1 0 63756 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1636993656
transform 1 0 63940 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1636993656
transform 1 0 65044 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1636993656
transform 1 0 66148 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1636993656
transform 1 0 67252 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 25201
transform 1 0 68356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 25201
transform 1 0 68908 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_729
timestamp 1636993656
transform 1 0 69092 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_741
timestamp 1636993656
transform 1 0 70196 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1636993656
transform 1 0 71300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1636993656
transform 1 0 72404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 25201
transform 1 0 73508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 25201
transform 1 0 74060 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_785
timestamp 1636993656
transform 1 0 74244 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_797
timestamp 1636993656
transform 1 0 75348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_809
timestamp 1636993656
transform 1 0 76452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_821
timestamp 25201
transform 1 0 77556 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636993656
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636993656
transform 1 0 3404 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 25201
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636993656
transform 1 0 4692 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636993656
transform 1 0 5796 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636993656
transform 1 0 6900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1636993656
transform 1 0 8004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 25201
transform 1 0 9108 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 25201
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1636993656
transform 1 0 9844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_97
timestamp 25201
transform 1 0 10948 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_108
timestamp 1636993656
transform 1 0 11960 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_120
timestamp 1636993656
transform 1 0 13064 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp 25201
transform 1 0 14168 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636993656
transform 1 0 14996 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636993656
transform 1 0 16100 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_176
timestamp 25201
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_224
timestamp 25201
transform 1 0 22632 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_255
timestamp 25201
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_299
timestamp 25201
transform 1 0 29532 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_339
timestamp 25201
transform 1 0 33212 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 25201
transform 1 0 35144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_381
timestamp 25201
transform 1 0 37076 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_402
timestamp 1636993656
transform 1 0 39008 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_414
timestamp 25201
transform 1 0 40112 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1636993656
transform 1 0 40756 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1636993656
transform 1 0 41860 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1636993656
transform 1 0 42964 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1636993656
transform 1 0 44068 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 25201
transform 1 0 45172 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 25201
transform 1 0 45724 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1636993656
transform 1 0 45908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1636993656
transform 1 0 47012 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1636993656
transform 1 0 48116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1636993656
transform 1 0 49220 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 25201
transform 1 0 50324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 25201
transform 1 0 50876 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1636993656
transform 1 0 51060 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1636993656
transform 1 0 52164 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1636993656
transform 1 0 53268 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1636993656
transform 1 0 54372 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 25201
transform 1 0 55476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 25201
transform 1 0 56028 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1636993656
transform 1 0 56212 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1636993656
transform 1 0 57316 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1636993656
transform 1 0 58420 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1636993656
transform 1 0 59524 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 25201
transform 1 0 60628 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 25201
transform 1 0 61180 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1636993656
transform 1 0 61364 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1636993656
transform 1 0 62468 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1636993656
transform 1 0 63572 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1636993656
transform 1 0 64676 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 25201
transform 1 0 65780 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 25201
transform 1 0 66332 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1636993656
transform 1 0 66516 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1636993656
transform 1 0 67620 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_725
timestamp 1636993656
transform 1 0 68724 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_737
timestamp 1636993656
transform 1 0 69828 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 25201
transform 1 0 70932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 25201
transform 1 0 71484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1636993656
transform 1 0 71668 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1636993656
transform 1 0 72772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1636993656
transform 1 0 73876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_793
timestamp 1636993656
transform 1 0 74980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 25201
transform 1 0 76084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 25201
transform 1 0 76636 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_813
timestamp 25201
transform 1 0 76820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_821
timestamp 25201
transform 1 0 77556 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636993656
transform 1 0 2300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636993656
transform 1 0 3404 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636993656
transform 1 0 4508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636993656
transform 1 0 5612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 25201
transform 1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 25201
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636993656
transform 1 0 7268 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1636993656
transform 1 0 8372 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1636993656
transform 1 0 9476 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1636993656
transform 1 0 10580 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 25201
transform 1 0 11684 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 25201
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1636993656
transform 1 0 12420 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1636993656
transform 1 0 13524 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1636993656
transform 1 0 14628 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1636993656
transform 1 0 15732 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 25201
transform 1 0 16836 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 25201
transform 1 0 17388 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636993656
transform 1 0 17572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_211
timestamp 25201
transform 1 0 21436 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_262
timestamp 25201
transform 1 0 26128 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_274
timestamp 25201
transform 1 0 27232 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_360
timestamp 25201
transform 1 0 35144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 25201
transform 1 0 37444 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 25201
transform 1 0 37996 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_401
timestamp 1636993656
transform 1 0 38916 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_413
timestamp 1636993656
transform 1 0 40020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_425
timestamp 1636993656
transform 1 0 41124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_437
timestamp 25201
transform 1 0 42228 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_445
timestamp 25201
transform 1 0 42964 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1636993656
transform 1 0 43332 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1636993656
transform 1 0 44436 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1636993656
transform 1 0 45540 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1636993656
transform 1 0 46644 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 25201
transform 1 0 47748 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 25201
transform 1 0 48300 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1636993656
transform 1 0 48484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1636993656
transform 1 0 49588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1636993656
transform 1 0 50692 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1636993656
transform 1 0 51796 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 25201
transform 1 0 52900 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 25201
transform 1 0 53452 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1636993656
transform 1 0 53636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1636993656
transform 1 0 54740 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1636993656
transform 1 0 55844 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1636993656
transform 1 0 56948 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 25201
transform 1 0 58052 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 25201
transform 1 0 58604 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1636993656
transform 1 0 58788 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1636993656
transform 1 0 59892 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1636993656
transform 1 0 60996 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1636993656
transform 1 0 62100 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 25201
transform 1 0 63204 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 25201
transform 1 0 63756 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1636993656
transform 1 0 63940 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1636993656
transform 1 0 65044 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1636993656
transform 1 0 66148 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1636993656
transform 1 0 67252 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 25201
transform 1 0 68356 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 25201
transform 1 0 68908 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_729
timestamp 1636993656
transform 1 0 69092 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_741
timestamp 1636993656
transform 1 0 70196 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_753
timestamp 1636993656
transform 1 0 71300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_765
timestamp 1636993656
transform 1 0 72404 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 25201
transform 1 0 73508 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 25201
transform 1 0 74060 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_785
timestamp 1636993656
transform 1 0 74244 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_797
timestamp 1636993656
transform 1 0 75348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_809
timestamp 1636993656
transform 1 0 76452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_821
timestamp 25201
transform 1 0 77556 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636993656
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636993656
transform 1 0 3404 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 25201
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636993656
transform 1 0 4692 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636993656
transform 1 0 5796 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636993656
transform 1 0 6900 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1636993656
transform 1 0 8004 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 25201
transform 1 0 9108 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 25201
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636993656
transform 1 0 9844 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1636993656
transform 1 0 10948 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1636993656
transform 1 0 12052 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1636993656
transform 1 0 13156 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 25201
transform 1 0 14260 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 25201
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1636993656
transform 1 0 14996 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1636993656
transform 1 0 16100 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1636993656
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1636993656
transform 1 0 18308 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 25201
transform 1 0 19412 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 25201
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_217
timestamp 25201
transform 1 0 21988 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_242
timestamp 25201
transform 1 0 24288 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_291
timestamp 25201
transform 1 0 28796 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_294
timestamp 25201
transform 1 0 29072 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_341
timestamp 25201
transform 1 0 33396 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_358
timestamp 25201
transform 1 0 34960 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_373
timestamp 25201
transform 1 0 36340 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_384
timestamp 1636993656
transform 1 0 37352 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_396
timestamp 1636993656
transform 1 0 38456 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_408
timestamp 1636993656
transform 1 0 39560 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1636993656
transform 1 0 40756 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1636993656
transform 1 0 41860 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1636993656
transform 1 0 42964 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1636993656
transform 1 0 44068 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 25201
transform 1 0 45172 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 25201
transform 1 0 45724 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1636993656
transform 1 0 45908 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1636993656
transform 1 0 47012 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1636993656
transform 1 0 48116 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1636993656
transform 1 0 49220 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 25201
transform 1 0 50324 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 25201
transform 1 0 50876 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1636993656
transform 1 0 51060 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1636993656
transform 1 0 52164 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1636993656
transform 1 0 53268 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1636993656
transform 1 0 54372 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 25201
transform 1 0 55476 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 25201
transform 1 0 56028 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1636993656
transform 1 0 56212 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1636993656
transform 1 0 57316 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1636993656
transform 1 0 58420 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1636993656
transform 1 0 59524 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 25201
transform 1 0 60628 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 25201
transform 1 0 61180 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1636993656
transform 1 0 61364 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1636993656
transform 1 0 62468 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1636993656
transform 1 0 63572 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1636993656
transform 1 0 64676 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 25201
transform 1 0 65780 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 25201
transform 1 0 66332 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1636993656
transform 1 0 66516 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1636993656
transform 1 0 67620 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_725
timestamp 1636993656
transform 1 0 68724 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_737
timestamp 1636993656
transform 1 0 69828 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 25201
transform 1 0 70932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 25201
transform 1 0 71484 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_757
timestamp 1636993656
transform 1 0 71668 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_769
timestamp 1636993656
transform 1 0 72772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_781
timestamp 1636993656
transform 1 0 73876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_793
timestamp 1636993656
transform 1 0 74980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 25201
transform 1 0 76084 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 25201
transform 1 0 76636 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_813
timestamp 25201
transform 1 0 76820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_821
timestamp 25201
transform 1 0 77556 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636993656
transform 1 0 2300 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636993656
transform 1 0 3404 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636993656
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636993656
transform 1 0 5612 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 25201
transform 1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 25201
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636993656
transform 1 0 7268 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1636993656
transform 1 0 8372 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1636993656
transform 1 0 9476 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1636993656
transform 1 0 10580 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 25201
transform 1 0 11684 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 25201
transform 1 0 12236 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1636993656
transform 1 0 12420 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1636993656
transform 1 0 13524 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1636993656
transform 1 0 14628 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1636993656
transform 1 0 15732 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 25201
transform 1 0 16836 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 25201
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1636993656
transform 1 0 17572 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1636993656
transform 1 0 18676 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_193
timestamp 25201
transform 1 0 19780 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_199
timestamp 25201
transform 1 0 20332 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_205
timestamp 25201
transform 1 0 20884 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_242
timestamp 25201
transform 1 0 24288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_252
timestamp 25201
transform 1 0 25208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_271
timestamp 25201
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_322
timestamp 1636993656
transform 1 0 31648 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 25201
transform 1 0 32752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_354
timestamp 25201
transform 1 0 34592 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_364
timestamp 1636993656
transform 1 0 35512 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_376
timestamp 1636993656
transform 1 0 36616 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_388
timestamp 25201
transform 1 0 37720 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1636993656
transform 1 0 38180 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1636993656
transform 1 0 39284 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1636993656
transform 1 0 40388 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1636993656
transform 1 0 41492 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 25201
transform 1 0 42596 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 25201
transform 1 0 43148 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1636993656
transform 1 0 43332 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1636993656
transform 1 0 44436 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1636993656
transform 1 0 45540 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1636993656
transform 1 0 46644 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 25201
transform 1 0 47748 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 25201
transform 1 0 48300 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1636993656
transform 1 0 48484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1636993656
transform 1 0 49588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1636993656
transform 1 0 50692 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1636993656
transform 1 0 51796 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 25201
transform 1 0 52900 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 25201
transform 1 0 53452 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1636993656
transform 1 0 53636 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1636993656
transform 1 0 54740 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1636993656
transform 1 0 55844 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1636993656
transform 1 0 56948 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 25201
transform 1 0 58052 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 25201
transform 1 0 58604 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1636993656
transform 1 0 58788 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1636993656
transform 1 0 59892 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1636993656
transform 1 0 60996 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1636993656
transform 1 0 62100 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 25201
transform 1 0 63204 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 25201
transform 1 0 63756 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1636993656
transform 1 0 63940 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1636993656
transform 1 0 65044 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1636993656
transform 1 0 66148 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1636993656
transform 1 0 67252 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 25201
transform 1 0 68356 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 25201
transform 1 0 68908 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_729
timestamp 1636993656
transform 1 0 69092 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_741
timestamp 1636993656
transform 1 0 70196 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_753
timestamp 1636993656
transform 1 0 71300 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_765
timestamp 1636993656
transform 1 0 72404 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 25201
transform 1 0 73508 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 25201
transform 1 0 74060 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_785
timestamp 1636993656
transform 1 0 74244 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_797
timestamp 1636993656
transform 1 0 75348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_809
timestamp 1636993656
transform 1 0 76452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_821
timestamp 25201
transform 1 0 77556 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636993656
transform 1 0 2300 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636993656
transform 1 0 3404 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 25201
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636993656
transform 1 0 4692 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636993656
transform 1 0 5796 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636993656
transform 1 0 6900 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1636993656
transform 1 0 8004 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 25201
transform 1 0 9108 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 25201
transform 1 0 9660 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636993656
transform 1 0 9844 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1636993656
transform 1 0 10948 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1636993656
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1636993656
transform 1 0 13156 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 25201
transform 1 0 14260 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 25201
transform 1 0 14812 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636993656
transform 1 0 14996 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1636993656
transform 1 0 16100 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1636993656
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1636993656
transform 1 0 18308 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 25201
transform 1 0 19412 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 25201
transform 1 0 19964 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1636993656
transform 1 0 20148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_209
timestamp 25201
transform 1 0 21252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_215
timestamp 25201
transform 1 0 21804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_223
timestamp 25201
transform 1 0 22540 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 25201
transform 1 0 23092 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 25201
transform 1 0 25024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_260
timestamp 25201
transform 1 0 25944 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_268
timestamp 25201
transform 1 0 26680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_277
timestamp 25201
transform 1 0 27508 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_281
timestamp 25201
transform 1 0 27876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_293
timestamp 25201
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 25201
transform 1 0 29900 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 25201
transform 1 0 30268 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1636993656
transform 1 0 30452 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1636993656
transform 1 0 31556 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1636993656
transform 1 0 32660 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1636993656
transform 1 0 33764 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 25201
transform 1 0 34868 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 25201
transform 1 0 35420 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1636993656
transform 1 0 35604 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1636993656
transform 1 0 36708 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1636993656
transform 1 0 37812 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1636993656
transform 1 0 38916 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 25201
transform 1 0 40020 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 25201
transform 1 0 40572 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1636993656
transform 1 0 40756 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1636993656
transform 1 0 41860 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1636993656
transform 1 0 42964 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1636993656
transform 1 0 44068 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 25201
transform 1 0 45172 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 25201
transform 1 0 45724 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1636993656
transform 1 0 45908 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1636993656
transform 1 0 47012 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1636993656
transform 1 0 48116 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1636993656
transform 1 0 49220 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 25201
transform 1 0 50324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 25201
transform 1 0 50876 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1636993656
transform 1 0 51060 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1636993656
transform 1 0 52164 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1636993656
transform 1 0 53268 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1636993656
transform 1 0 54372 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 25201
transform 1 0 55476 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 25201
transform 1 0 56028 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1636993656
transform 1 0 56212 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1636993656
transform 1 0 57316 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1636993656
transform 1 0 58420 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1636993656
transform 1 0 59524 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 25201
transform 1 0 60628 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 25201
transform 1 0 61180 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1636993656
transform 1 0 61364 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1636993656
transform 1 0 62468 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1636993656
transform 1 0 63572 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1636993656
transform 1 0 64676 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 25201
transform 1 0 65780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 25201
transform 1 0 66332 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1636993656
transform 1 0 66516 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1636993656
transform 1 0 67620 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_725
timestamp 1636993656
transform 1 0 68724 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_737
timestamp 1636993656
transform 1 0 69828 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 25201
transform 1 0 70932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 25201
transform 1 0 71484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_757
timestamp 1636993656
transform 1 0 71668 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_769
timestamp 1636993656
transform 1 0 72772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_781
timestamp 1636993656
transform 1 0 73876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_793
timestamp 1636993656
transform 1 0 74980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 25201
transform 1 0 76084 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 25201
transform 1 0 76636 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_813
timestamp 25201
transform 1 0 76820 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_821
timestamp 25201
transform 1 0 77556 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636993656
transform 1 0 2300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636993656
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1636993656
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1636993656
transform 1 0 5612 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 25201
transform 1 0 6716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 25201
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636993656
transform 1 0 7268 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636993656
transform 1 0 8372 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1636993656
transform 1 0 9476 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1636993656
transform 1 0 10580 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 25201
transform 1 0 11684 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 25201
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636993656
transform 1 0 12420 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1636993656
transform 1 0 13524 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1636993656
transform 1 0 14628 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1636993656
transform 1 0 15732 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 25201
transform 1 0 16836 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 25201
transform 1 0 17388 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636993656
transform 1 0 17572 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1636993656
transform 1 0 18676 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1636993656
transform 1 0 19780 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1636993656
transform 1 0 20884 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 25201
transform 1 0 21988 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 25201
transform 1 0 22540 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1636993656
transform 1 0 22724 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1636993656
transform 1 0 23828 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1636993656
transform 1 0 24932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1636993656
transform 1 0 26036 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 25201
transform 1 0 27140 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 25201
transform 1 0 27692 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_281
timestamp 25201
transform 1 0 27876 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_287
timestamp 25201
transform 1 0 28428 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_302
timestamp 1636993656
transform 1 0 29808 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_314
timestamp 1636993656
transform 1 0 30912 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_326
timestamp 25201
transform 1 0 32016 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 25201
transform 1 0 32752 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1636993656
transform 1 0 33028 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1636993656
transform 1 0 34132 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1636993656
transform 1 0 35236 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1636993656
transform 1 0 36340 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 25201
transform 1 0 37444 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 25201
transform 1 0 37996 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1636993656
transform 1 0 38180 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1636993656
transform 1 0 39284 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1636993656
transform 1 0 40388 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1636993656
transform 1 0 41492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 25201
transform 1 0 42596 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 25201
transform 1 0 43148 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1636993656
transform 1 0 43332 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1636993656
transform 1 0 44436 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1636993656
transform 1 0 45540 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1636993656
transform 1 0 46644 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 25201
transform 1 0 47748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 25201
transform 1 0 48300 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1636993656
transform 1 0 48484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1636993656
transform 1 0 49588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1636993656
transform 1 0 50692 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1636993656
transform 1 0 51796 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 25201
transform 1 0 52900 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 25201
transform 1 0 53452 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1636993656
transform 1 0 53636 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1636993656
transform 1 0 54740 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1636993656
transform 1 0 55844 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1636993656
transform 1 0 56948 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 25201
transform 1 0 58052 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 25201
transform 1 0 58604 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1636993656
transform 1 0 58788 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1636993656
transform 1 0 59892 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1636993656
transform 1 0 60996 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1636993656
transform 1 0 62100 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 25201
transform 1 0 63204 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 25201
transform 1 0 63756 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1636993656
transform 1 0 63940 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1636993656
transform 1 0 65044 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1636993656
transform 1 0 66148 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1636993656
transform 1 0 67252 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 25201
transform 1 0 68356 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 25201
transform 1 0 68908 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_729
timestamp 1636993656
transform 1 0 69092 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_741
timestamp 1636993656
transform 1 0 70196 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_753
timestamp 1636993656
transform 1 0 71300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_765
timestamp 1636993656
transform 1 0 72404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 25201
transform 1 0 73508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 25201
transform 1 0 74060 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_785
timestamp 1636993656
transform 1 0 74244 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_797
timestamp 1636993656
transform 1 0 75348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_809
timestamp 1636993656
transform 1 0 76452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_821
timestamp 25201
transform 1 0 77556 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636993656
transform 1 0 2300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636993656
transform 1 0 3404 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 25201
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636993656
transform 1 0 4692 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636993656
transform 1 0 5796 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636993656
transform 1 0 6900 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1636993656
transform 1 0 8004 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 25201
transform 1 0 9108 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 25201
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636993656
transform 1 0 9844 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636993656
transform 1 0 10948 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1636993656
transform 1 0 12052 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1636993656
transform 1 0 13156 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 25201
transform 1 0 14260 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 25201
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636993656
transform 1 0 14996 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636993656
transform 1 0 16100 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1636993656
transform 1 0 17204 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1636993656
transform 1 0 18308 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 25201
transform 1 0 19412 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 25201
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1636993656
transform 1 0 20148 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1636993656
transform 1 0 21252 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1636993656
transform 1 0 22356 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1636993656
transform 1 0 23460 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 25201
transform 1 0 24564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 25201
transform 1 0 25116 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1636993656
transform 1 0 25300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1636993656
transform 1 0 26404 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1636993656
transform 1 0 27508 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1636993656
transform 1 0 28612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 25201
transform 1 0 29716 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 25201
transform 1 0 30268 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1636993656
transform 1 0 30452 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1636993656
transform 1 0 31556 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1636993656
transform 1 0 32660 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1636993656
transform 1 0 33764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 25201
transform 1 0 34868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 25201
transform 1 0 35420 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1636993656
transform 1 0 35604 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1636993656
transform 1 0 36708 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1636993656
transform 1 0 37812 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1636993656
transform 1 0 38916 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 25201
transform 1 0 40020 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 25201
transform 1 0 40572 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1636993656
transform 1 0 40756 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1636993656
transform 1 0 41860 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1636993656
transform 1 0 42964 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1636993656
transform 1 0 44068 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 25201
transform 1 0 45172 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 25201
transform 1 0 45724 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1636993656
transform 1 0 45908 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1636993656
transform 1 0 47012 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1636993656
transform 1 0 48116 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1636993656
transform 1 0 49220 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 25201
transform 1 0 50324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 25201
transform 1 0 50876 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1636993656
transform 1 0 51060 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1636993656
transform 1 0 52164 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1636993656
transform 1 0 53268 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1636993656
transform 1 0 54372 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 25201
transform 1 0 55476 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 25201
transform 1 0 56028 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1636993656
transform 1 0 56212 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1636993656
transform 1 0 57316 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1636993656
transform 1 0 58420 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1636993656
transform 1 0 59524 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 25201
transform 1 0 60628 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 25201
transform 1 0 61180 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1636993656
transform 1 0 61364 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1636993656
transform 1 0 62468 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1636993656
transform 1 0 63572 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1636993656
transform 1 0 64676 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 25201
transform 1 0 65780 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 25201
transform 1 0 66332 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1636993656
transform 1 0 66516 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1636993656
transform 1 0 67620 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_725
timestamp 1636993656
transform 1 0 68724 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_737
timestamp 1636993656
transform 1 0 69828 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 25201
transform 1 0 70932 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 25201
transform 1 0 71484 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_757
timestamp 1636993656
transform 1 0 71668 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_769
timestamp 1636993656
transform 1 0 72772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_781
timestamp 1636993656
transform 1 0 73876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_793
timestamp 1636993656
transform 1 0 74980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_805
timestamp 25201
transform 1 0 76084 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_811
timestamp 25201
transform 1 0 76636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_813
timestamp 25201
transform 1 0 76820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_821
timestamp 25201
transform 1 0 77556 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636993656
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636993656
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636993656
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1636993656
transform 1 0 5612 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 25201
transform 1 0 6716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 25201
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636993656
transform 1 0 7268 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1636993656
transform 1 0 8372 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1636993656
transform 1 0 9476 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1636993656
transform 1 0 10580 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 25201
transform 1 0 11684 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 25201
transform 1 0 12236 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636993656
transform 1 0 12420 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1636993656
transform 1 0 13524 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1636993656
transform 1 0 14628 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1636993656
transform 1 0 15732 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 25201
transform 1 0 16836 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 25201
transform 1 0 17388 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636993656
transform 1 0 17572 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1636993656
transform 1 0 18676 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1636993656
transform 1 0 19780 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1636993656
transform 1 0 20884 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 25201
transform 1 0 21988 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 25201
transform 1 0 22540 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636993656
transform 1 0 22724 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1636993656
transform 1 0 23828 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1636993656
transform 1 0 24932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1636993656
transform 1 0 26036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 25201
transform 1 0 27140 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 25201
transform 1 0 27692 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1636993656
transform 1 0 27876 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1636993656
transform 1 0 28980 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1636993656
transform 1 0 30084 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1636993656
transform 1 0 31188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 25201
transform 1 0 32292 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 25201
transform 1 0 32844 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1636993656
transform 1 0 33028 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1636993656
transform 1 0 34132 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1636993656
transform 1 0 35236 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1636993656
transform 1 0 36340 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 25201
transform 1 0 37444 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 25201
transform 1 0 37996 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1636993656
transform 1 0 38180 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1636993656
transform 1 0 39284 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1636993656
transform 1 0 40388 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1636993656
transform 1 0 41492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 25201
transform 1 0 42596 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 25201
transform 1 0 43148 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1636993656
transform 1 0 43332 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1636993656
transform 1 0 44436 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1636993656
transform 1 0 45540 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1636993656
transform 1 0 46644 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 25201
transform 1 0 47748 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 25201
transform 1 0 48300 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1636993656
transform 1 0 48484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1636993656
transform 1 0 49588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1636993656
transform 1 0 50692 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1636993656
transform 1 0 51796 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 25201
transform 1 0 52900 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 25201
transform 1 0 53452 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1636993656
transform 1 0 53636 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1636993656
transform 1 0 54740 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1636993656
transform 1 0 55844 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1636993656
transform 1 0 56948 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 25201
transform 1 0 58052 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 25201
transform 1 0 58604 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1636993656
transform 1 0 58788 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1636993656
transform 1 0 59892 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1636993656
transform 1 0 60996 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1636993656
transform 1 0 62100 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 25201
transform 1 0 63204 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 25201
transform 1 0 63756 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1636993656
transform 1 0 63940 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1636993656
transform 1 0 65044 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1636993656
transform 1 0 66148 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1636993656
transform 1 0 67252 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 25201
transform 1 0 68356 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 25201
transform 1 0 68908 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_729
timestamp 1636993656
transform 1 0 69092 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_741
timestamp 1636993656
transform 1 0 70196 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_753
timestamp 1636993656
transform 1 0 71300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_765
timestamp 1636993656
transform 1 0 72404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_777
timestamp 25201
transform 1 0 73508 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 25201
transform 1 0 74060 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_785
timestamp 1636993656
transform 1 0 74244 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_797
timestamp 1636993656
transform 1 0 75348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_809
timestamp 1636993656
transform 1 0 76452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_821
timestamp 25201
transform 1 0 77556 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636993656
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636993656
transform 1 0 3404 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 25201
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636993656
transform 1 0 4692 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636993656
transform 1 0 5796 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636993656
transform 1 0 6900 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1636993656
transform 1 0 8004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 25201
transform 1 0 9108 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 25201
transform 1 0 9660 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636993656
transform 1 0 9844 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1636993656
transform 1 0 10948 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1636993656
transform 1 0 12052 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1636993656
transform 1 0 13156 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 25201
transform 1 0 14260 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 25201
transform 1 0 14812 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1636993656
transform 1 0 14996 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1636993656
transform 1 0 16100 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1636993656
transform 1 0 17204 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1636993656
transform 1 0 18308 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 25201
transform 1 0 19412 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 25201
transform 1 0 19964 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1636993656
transform 1 0 20148 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1636993656
transform 1 0 21252 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1636993656
transform 1 0 22356 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1636993656
transform 1 0 23460 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 25201
transform 1 0 24564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 25201
transform 1 0 25116 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1636993656
transform 1 0 25300 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1636993656
transform 1 0 26404 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1636993656
transform 1 0 27508 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1636993656
transform 1 0 28612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 25201
transform 1 0 29716 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 25201
transform 1 0 30268 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1636993656
transform 1 0 30452 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1636993656
transform 1 0 31556 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1636993656
transform 1 0 32660 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1636993656
transform 1 0 33764 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 25201
transform 1 0 34868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 25201
transform 1 0 35420 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1636993656
transform 1 0 35604 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1636993656
transform 1 0 36708 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1636993656
transform 1 0 37812 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1636993656
transform 1 0 38916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 25201
transform 1 0 40020 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 25201
transform 1 0 40572 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1636993656
transform 1 0 40756 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1636993656
transform 1 0 41860 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1636993656
transform 1 0 42964 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1636993656
transform 1 0 44068 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 25201
transform 1 0 45172 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 25201
transform 1 0 45724 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1636993656
transform 1 0 45908 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1636993656
transform 1 0 47012 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1636993656
transform 1 0 48116 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1636993656
transform 1 0 49220 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 25201
transform 1 0 50324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 25201
transform 1 0 50876 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1636993656
transform 1 0 51060 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1636993656
transform 1 0 52164 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1636993656
transform 1 0 53268 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1636993656
transform 1 0 54372 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 25201
transform 1 0 55476 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 25201
transform 1 0 56028 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1636993656
transform 1 0 56212 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1636993656
transform 1 0 57316 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1636993656
transform 1 0 58420 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1636993656
transform 1 0 59524 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 25201
transform 1 0 60628 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 25201
transform 1 0 61180 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1636993656
transform 1 0 61364 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1636993656
transform 1 0 62468 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1636993656
transform 1 0 63572 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1636993656
transform 1 0 64676 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 25201
transform 1 0 65780 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 25201
transform 1 0 66332 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1636993656
transform 1 0 66516 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_713
timestamp 1636993656
transform 1 0 67620 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_725
timestamp 1636993656
transform 1 0 68724 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_737
timestamp 1636993656
transform 1 0 69828 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_749
timestamp 25201
transform 1 0 70932 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_755
timestamp 25201
transform 1 0 71484 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_757
timestamp 1636993656
transform 1 0 71668 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_769
timestamp 1636993656
transform 1 0 72772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_781
timestamp 1636993656
transform 1 0 73876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_793
timestamp 1636993656
transform 1 0 74980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_805
timestamp 25201
transform 1 0 76084 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_811
timestamp 25201
transform 1 0 76636 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_813
timestamp 25201
transform 1 0 76820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_821
timestamp 25201
transform 1 0 77556 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636993656
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636993656
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636993656
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1636993656
transform 1 0 5612 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 25201
transform 1 0 6716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 25201
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636993656
transform 1 0 7268 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1636993656
transform 1 0 8372 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1636993656
transform 1 0 9476 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1636993656
transform 1 0 10580 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 25201
transform 1 0 11684 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 25201
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1636993656
transform 1 0 12420 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1636993656
transform 1 0 13524 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1636993656
transform 1 0 14628 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1636993656
transform 1 0 15732 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 25201
transform 1 0 16836 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 25201
transform 1 0 17388 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1636993656
transform 1 0 17572 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1636993656
transform 1 0 18676 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1636993656
transform 1 0 19780 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1636993656
transform 1 0 20884 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 25201
transform 1 0 21988 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 25201
transform 1 0 22540 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1636993656
transform 1 0 22724 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1636993656
transform 1 0 23828 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1636993656
transform 1 0 24932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1636993656
transform 1 0 26036 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 25201
transform 1 0 27140 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 25201
transform 1 0 27692 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1636993656
transform 1 0 27876 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1636993656
transform 1 0 28980 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1636993656
transform 1 0 30084 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1636993656
transform 1 0 31188 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 25201
transform 1 0 32292 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 25201
transform 1 0 32844 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1636993656
transform 1 0 33028 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1636993656
transform 1 0 34132 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1636993656
transform 1 0 35236 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1636993656
transform 1 0 36340 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 25201
transform 1 0 37444 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 25201
transform 1 0 37996 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1636993656
transform 1 0 38180 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1636993656
transform 1 0 39284 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1636993656
transform 1 0 40388 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1636993656
transform 1 0 41492 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 25201
transform 1 0 42596 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 25201
transform 1 0 43148 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1636993656
transform 1 0 43332 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1636993656
transform 1 0 44436 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1636993656
transform 1 0 45540 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1636993656
transform 1 0 46644 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 25201
transform 1 0 47748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 25201
transform 1 0 48300 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1636993656
transform 1 0 48484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1636993656
transform 1 0 49588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1636993656
transform 1 0 50692 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1636993656
transform 1 0 51796 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 25201
transform 1 0 52900 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 25201
transform 1 0 53452 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1636993656
transform 1 0 53636 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1636993656
transform 1 0 54740 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1636993656
transform 1 0 55844 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1636993656
transform 1 0 56948 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 25201
transform 1 0 58052 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 25201
transform 1 0 58604 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1636993656
transform 1 0 58788 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1636993656
transform 1 0 59892 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1636993656
transform 1 0 60996 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1636993656
transform 1 0 62100 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 25201
transform 1 0 63204 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 25201
transform 1 0 63756 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1636993656
transform 1 0 63940 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1636993656
transform 1 0 65044 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_697
timestamp 1636993656
transform 1 0 66148 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_709
timestamp 1636993656
transform 1 0 67252 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 25201
transform 1 0 68356 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 25201
transform 1 0 68908 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_729
timestamp 1636993656
transform 1 0 69092 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_741
timestamp 1636993656
transform 1 0 70196 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_753
timestamp 1636993656
transform 1 0 71300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_765
timestamp 1636993656
transform 1 0 72404 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_777
timestamp 25201
transform 1 0 73508 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_783
timestamp 25201
transform 1 0 74060 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_785
timestamp 1636993656
transform 1 0 74244 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_797
timestamp 1636993656
transform 1 0 75348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_809
timestamp 1636993656
transform 1 0 76452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_821
timestamp 25201
transform 1 0 77556 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636993656
transform 1 0 2300 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636993656
transform 1 0 3404 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 25201
transform 1 0 4508 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636993656
transform 1 0 4692 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636993656
transform 1 0 5796 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636993656
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1636993656
transform 1 0 8004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 25201
transform 1 0 9108 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 25201
transform 1 0 9660 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636993656
transform 1 0 9844 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1636993656
transform 1 0 10948 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1636993656
transform 1 0 12052 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1636993656
transform 1 0 13156 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 25201
transform 1 0 14260 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 25201
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636993656
transform 1 0 14996 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1636993656
transform 1 0 16100 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1636993656
transform 1 0 17204 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1636993656
transform 1 0 18308 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 25201
transform 1 0 19412 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 25201
transform 1 0 19964 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1636993656
transform 1 0 20148 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1636993656
transform 1 0 21252 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1636993656
transform 1 0 22356 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1636993656
transform 1 0 23460 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 25201
transform 1 0 24564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 25201
transform 1 0 25116 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1636993656
transform 1 0 25300 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1636993656
transform 1 0 26404 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1636993656
transform 1 0 27508 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1636993656
transform 1 0 28612 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 25201
transform 1 0 29716 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 25201
transform 1 0 30268 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1636993656
transform 1 0 30452 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1636993656
transform 1 0 31556 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1636993656
transform 1 0 32660 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1636993656
transform 1 0 33764 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 25201
transform 1 0 34868 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 25201
transform 1 0 35420 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1636993656
transform 1 0 35604 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1636993656
transform 1 0 36708 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1636993656
transform 1 0 37812 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1636993656
transform 1 0 38916 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 25201
transform 1 0 40020 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 25201
transform 1 0 40572 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1636993656
transform 1 0 40756 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1636993656
transform 1 0 41860 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1636993656
transform 1 0 42964 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1636993656
transform 1 0 44068 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 25201
transform 1 0 45172 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 25201
transform 1 0 45724 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1636993656
transform 1 0 45908 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1636993656
transform 1 0 47012 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1636993656
transform 1 0 48116 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1636993656
transform 1 0 49220 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 25201
transform 1 0 50324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 25201
transform 1 0 50876 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1636993656
transform 1 0 51060 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1636993656
transform 1 0 52164 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1636993656
transform 1 0 53268 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1636993656
transform 1 0 54372 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 25201
transform 1 0 55476 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 25201
transform 1 0 56028 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1636993656
transform 1 0 56212 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1636993656
transform 1 0 57316 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1636993656
transform 1 0 58420 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_625
timestamp 1636993656
transform 1 0 59524 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 25201
transform 1 0 60628 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 25201
transform 1 0 61180 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1636993656
transform 1 0 61364 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1636993656
transform 1 0 62468 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1636993656
transform 1 0 63572 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_681
timestamp 1636993656
transform 1 0 64676 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 25201
transform 1 0 65780 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 25201
transform 1 0 66332 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_701
timestamp 1636993656
transform 1 0 66516 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_713
timestamp 1636993656
transform 1 0 67620 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_725
timestamp 1636993656
transform 1 0 68724 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_737
timestamp 1636993656
transform 1 0 69828 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_749
timestamp 25201
transform 1 0 70932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_755
timestamp 25201
transform 1 0 71484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_757
timestamp 1636993656
transform 1 0 71668 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_769
timestamp 1636993656
transform 1 0 72772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_781
timestamp 1636993656
transform 1 0 73876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_793
timestamp 1636993656
transform 1 0 74980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_805
timestamp 25201
transform 1 0 76084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_811
timestamp 25201
transform 1 0 76636 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_813
timestamp 25201
transform 1 0 76820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_821
timestamp 25201
transform 1 0 77556 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636993656
transform 1 0 2300 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636993656
transform 1 0 3404 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636993656
transform 1 0 4508 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636993656
transform 1 0 5612 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 25201
transform 1 0 6716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 25201
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636993656
transform 1 0 7268 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1636993656
transform 1 0 8372 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1636993656
transform 1 0 9476 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1636993656
transform 1 0 10580 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 25201
transform 1 0 11684 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 25201
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1636993656
transform 1 0 12420 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1636993656
transform 1 0 13524 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1636993656
transform 1 0 14628 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1636993656
transform 1 0 15732 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 25201
transform 1 0 16836 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 25201
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636993656
transform 1 0 17572 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1636993656
transform 1 0 18676 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1636993656
transform 1 0 19780 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1636993656
transform 1 0 20884 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 25201
transform 1 0 21988 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 25201
transform 1 0 22540 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1636993656
transform 1 0 22724 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1636993656
transform 1 0 23828 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1636993656
transform 1 0 24932 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1636993656
transform 1 0 26036 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 25201
transform 1 0 27140 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 25201
transform 1 0 27692 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1636993656
transform 1 0 27876 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1636993656
transform 1 0 28980 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1636993656
transform 1 0 30084 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1636993656
transform 1 0 31188 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 25201
transform 1 0 32292 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 25201
transform 1 0 32844 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1636993656
transform 1 0 33028 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1636993656
transform 1 0 34132 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1636993656
transform 1 0 35236 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1636993656
transform 1 0 36340 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 25201
transform 1 0 37444 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 25201
transform 1 0 37996 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1636993656
transform 1 0 38180 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1636993656
transform 1 0 39284 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1636993656
transform 1 0 40388 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1636993656
transform 1 0 41492 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 25201
transform 1 0 42596 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 25201
transform 1 0 43148 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1636993656
transform 1 0 43332 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1636993656
transform 1 0 44436 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1636993656
transform 1 0 45540 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1636993656
transform 1 0 46644 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 25201
transform 1 0 47748 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 25201
transform 1 0 48300 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1636993656
transform 1 0 48484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1636993656
transform 1 0 49588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1636993656
transform 1 0 50692 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1636993656
transform 1 0 51796 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 25201
transform 1 0 52900 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 25201
transform 1 0 53452 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1636993656
transform 1 0 53636 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1636993656
transform 1 0 54740 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1636993656
transform 1 0 55844 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1636993656
transform 1 0 56948 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 25201
transform 1 0 58052 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 25201
transform 1 0 58604 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1636993656
transform 1 0 58788 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1636993656
transform 1 0 59892 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1636993656
transform 1 0 60996 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1636993656
transform 1 0 62100 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 25201
transform 1 0 63204 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 25201
transform 1 0 63756 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_673
timestamp 1636993656
transform 1 0 63940 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_685
timestamp 1636993656
transform 1 0 65044 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_697
timestamp 1636993656
transform 1 0 66148 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_709
timestamp 1636993656
transform 1 0 67252 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 25201
transform 1 0 68356 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 25201
transform 1 0 68908 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_729
timestamp 1636993656
transform 1 0 69092 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_741
timestamp 1636993656
transform 1 0 70196 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_753
timestamp 1636993656
transform 1 0 71300 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_765
timestamp 1636993656
transform 1 0 72404 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_777
timestamp 25201
transform 1 0 73508 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_783
timestamp 25201
transform 1 0 74060 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_785
timestamp 1636993656
transform 1 0 74244 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_797
timestamp 1636993656
transform 1 0 75348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_809
timestamp 1636993656
transform 1 0 76452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_821
timestamp 25201
transform 1 0 77556 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636993656
transform 1 0 2300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636993656
transform 1 0 3404 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 25201
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636993656
transform 1 0 4692 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636993656
transform 1 0 5796 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636993656
transform 1 0 6900 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1636993656
transform 1 0 8004 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 25201
transform 1 0 9108 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 25201
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1636993656
transform 1 0 9844 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1636993656
transform 1 0 10948 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1636993656
transform 1 0 12052 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1636993656
transform 1 0 13156 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 25201
transform 1 0 14260 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 25201
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1636993656
transform 1 0 14996 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1636993656
transform 1 0 16100 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1636993656
transform 1 0 17204 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1636993656
transform 1 0 18308 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 25201
transform 1 0 19412 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 25201
transform 1 0 19964 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1636993656
transform 1 0 20148 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1636993656
transform 1 0 21252 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1636993656
transform 1 0 22356 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1636993656
transform 1 0 23460 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 25201
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 25201
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1636993656
transform 1 0 25300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1636993656
transform 1 0 26404 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1636993656
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1636993656
transform 1 0 28612 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 25201
transform 1 0 29716 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 25201
transform 1 0 30268 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1636993656
transform 1 0 30452 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1636993656
transform 1 0 31556 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1636993656
transform 1 0 32660 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1636993656
transform 1 0 33764 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 25201
transform 1 0 34868 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 25201
transform 1 0 35420 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1636993656
transform 1 0 35604 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1636993656
transform 1 0 36708 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1636993656
transform 1 0 37812 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1636993656
transform 1 0 38916 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 25201
transform 1 0 40020 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 25201
transform 1 0 40572 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1636993656
transform 1 0 40756 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1636993656
transform 1 0 41860 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1636993656
transform 1 0 42964 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1636993656
transform 1 0 44068 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 25201
transform 1 0 45172 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 25201
transform 1 0 45724 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1636993656
transform 1 0 45908 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1636993656
transform 1 0 47012 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1636993656
transform 1 0 48116 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1636993656
transform 1 0 49220 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 25201
transform 1 0 50324 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 25201
transform 1 0 50876 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1636993656
transform 1 0 51060 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1636993656
transform 1 0 52164 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1636993656
transform 1 0 53268 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1636993656
transform 1 0 54372 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 25201
transform 1 0 55476 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 25201
transform 1 0 56028 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1636993656
transform 1 0 56212 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1636993656
transform 1 0 57316 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1636993656
transform 1 0 58420 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1636993656
transform 1 0 59524 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 25201
transform 1 0 60628 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 25201
transform 1 0 61180 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1636993656
transform 1 0 61364 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1636993656
transform 1 0 62468 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1636993656
transform 1 0 63572 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_681
timestamp 1636993656
transform 1 0 64676 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 25201
transform 1 0 65780 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 25201
transform 1 0 66332 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_701
timestamp 1636993656
transform 1 0 66516 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_713
timestamp 1636993656
transform 1 0 67620 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_725
timestamp 1636993656
transform 1 0 68724 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_737
timestamp 1636993656
transform 1 0 69828 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_749
timestamp 25201
transform 1 0 70932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_755
timestamp 25201
transform 1 0 71484 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_757
timestamp 1636993656
transform 1 0 71668 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_769
timestamp 1636993656
transform 1 0 72772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_781
timestamp 1636993656
transform 1 0 73876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_793
timestamp 1636993656
transform 1 0 74980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_805
timestamp 25201
transform 1 0 76084 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_811
timestamp 25201
transform 1 0 76636 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_813
timestamp 25201
transform 1 0 76820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_821
timestamp 25201
transform 1 0 77556 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636993656
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636993656
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1636993656
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1636993656
transform 1 0 5612 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 25201
transform 1 0 6716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 25201
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636993656
transform 1 0 7268 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1636993656
transform 1 0 8372 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1636993656
transform 1 0 9476 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1636993656
transform 1 0 10580 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 25201
transform 1 0 11684 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 25201
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1636993656
transform 1 0 12420 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1636993656
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1636993656
transform 1 0 14628 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1636993656
transform 1 0 15732 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 25201
transform 1 0 16836 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 25201
transform 1 0 17388 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1636993656
transform 1 0 17572 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1636993656
transform 1 0 18676 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1636993656
transform 1 0 19780 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1636993656
transform 1 0 20884 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 25201
transform 1 0 21988 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 25201
transform 1 0 22540 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636993656
transform 1 0 22724 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1636993656
transform 1 0 23828 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1636993656
transform 1 0 24932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1636993656
transform 1 0 26036 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 25201
transform 1 0 27140 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 25201
transform 1 0 27692 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1636993656
transform 1 0 27876 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1636993656
transform 1 0 28980 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1636993656
transform 1 0 30084 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1636993656
transform 1 0 31188 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 25201
transform 1 0 32292 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 25201
transform 1 0 32844 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1636993656
transform 1 0 33028 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1636993656
transform 1 0 34132 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1636993656
transform 1 0 35236 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1636993656
transform 1 0 36340 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 25201
transform 1 0 37444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 25201
transform 1 0 37996 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1636993656
transform 1 0 38180 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1636993656
transform 1 0 39284 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1636993656
transform 1 0 40388 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1636993656
transform 1 0 41492 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 25201
transform 1 0 42596 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 25201
transform 1 0 43148 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1636993656
transform 1 0 43332 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1636993656
transform 1 0 44436 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1636993656
transform 1 0 45540 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1636993656
transform 1 0 46644 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 25201
transform 1 0 47748 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 25201
transform 1 0 48300 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1636993656
transform 1 0 48484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1636993656
transform 1 0 49588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1636993656
transform 1 0 50692 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1636993656
transform 1 0 51796 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 25201
transform 1 0 52900 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 25201
transform 1 0 53452 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1636993656
transform 1 0 53636 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1636993656
transform 1 0 54740 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1636993656
transform 1 0 55844 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1636993656
transform 1 0 56948 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 25201
transform 1 0 58052 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 25201
transform 1 0 58604 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1636993656
transform 1 0 58788 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1636993656
transform 1 0 59892 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1636993656
transform 1 0 60996 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1636993656
transform 1 0 62100 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 25201
transform 1 0 63204 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 25201
transform 1 0 63756 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1636993656
transform 1 0 63940 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1636993656
transform 1 0 65044 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1636993656
transform 1 0 66148 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_709
timestamp 1636993656
transform 1 0 67252 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 25201
transform 1 0 68356 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 25201
transform 1 0 68908 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_729
timestamp 1636993656
transform 1 0 69092 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_741
timestamp 1636993656
transform 1 0 70196 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_753
timestamp 1636993656
transform 1 0 71300 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_765
timestamp 1636993656
transform 1 0 72404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_777
timestamp 25201
transform 1 0 73508 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_783
timestamp 25201
transform 1 0 74060 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_785
timestamp 1636993656
transform 1 0 74244 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_797
timestamp 1636993656
transform 1 0 75348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_809
timestamp 1636993656
transform 1 0 76452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_821
timestamp 25201
transform 1 0 77556 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636993656
transform 1 0 2300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636993656
transform 1 0 3404 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 25201
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636993656
transform 1 0 4692 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636993656
transform 1 0 5796 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636993656
transform 1 0 6900 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1636993656
transform 1 0 8004 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 25201
transform 1 0 9108 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 25201
transform 1 0 9660 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636993656
transform 1 0 9844 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1636993656
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1636993656
transform 1 0 12052 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1636993656
transform 1 0 13156 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 25201
transform 1 0 14260 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 25201
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636993656
transform 1 0 14996 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1636993656
transform 1 0 16100 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1636993656
transform 1 0 17204 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1636993656
transform 1 0 18308 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 25201
transform 1 0 19412 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 25201
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636993656
transform 1 0 20148 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1636993656
transform 1 0 21252 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1636993656
transform 1 0 22356 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1636993656
transform 1 0 23460 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 25201
transform 1 0 24564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 25201
transform 1 0 25116 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1636993656
transform 1 0 25300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1636993656
transform 1 0 26404 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1636993656
transform 1 0 27508 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1636993656
transform 1 0 28612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 25201
transform 1 0 29716 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 25201
transform 1 0 30268 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1636993656
transform 1 0 30452 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1636993656
transform 1 0 31556 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1636993656
transform 1 0 32660 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1636993656
transform 1 0 33764 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 25201
transform 1 0 34868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 25201
transform 1 0 35420 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1636993656
transform 1 0 35604 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1636993656
transform 1 0 36708 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1636993656
transform 1 0 37812 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1636993656
transform 1 0 38916 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 25201
transform 1 0 40020 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 25201
transform 1 0 40572 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1636993656
transform 1 0 40756 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1636993656
transform 1 0 41860 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1636993656
transform 1 0 42964 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1636993656
transform 1 0 44068 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 25201
transform 1 0 45172 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 25201
transform 1 0 45724 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1636993656
transform 1 0 45908 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1636993656
transform 1 0 47012 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1636993656
transform 1 0 48116 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1636993656
transform 1 0 49220 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 25201
transform 1 0 50324 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 25201
transform 1 0 50876 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1636993656
transform 1 0 51060 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1636993656
transform 1 0 52164 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1636993656
transform 1 0 53268 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1636993656
transform 1 0 54372 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 25201
transform 1 0 55476 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 25201
transform 1 0 56028 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1636993656
transform 1 0 56212 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1636993656
transform 1 0 57316 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1636993656
transform 1 0 58420 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1636993656
transform 1 0 59524 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 25201
transform 1 0 60628 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 25201
transform 1 0 61180 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1636993656
transform 1 0 61364 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1636993656
transform 1 0 62468 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1636993656
transform 1 0 63572 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1636993656
transform 1 0 64676 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 25201
transform 1 0 65780 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 25201
transform 1 0 66332 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1636993656
transform 1 0 66516 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_713
timestamp 1636993656
transform 1 0 67620 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_725
timestamp 1636993656
transform 1 0 68724 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_737
timestamp 1636993656
transform 1 0 69828 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_749
timestamp 25201
transform 1 0 70932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_755
timestamp 25201
transform 1 0 71484 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_757
timestamp 1636993656
transform 1 0 71668 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_769
timestamp 1636993656
transform 1 0 72772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_781
timestamp 1636993656
transform 1 0 73876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_793
timestamp 1636993656
transform 1 0 74980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_805
timestamp 25201
transform 1 0 76084 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_811
timestamp 25201
transform 1 0 76636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_813
timestamp 25201
transform 1 0 76820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_821
timestamp 25201
transform 1 0 77556 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636993656
transform 1 0 2300 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636993656
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636993656
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636993656
transform 1 0 5612 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 25201
transform 1 0 6716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 25201
transform 1 0 7084 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636993656
transform 1 0 7268 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1636993656
transform 1 0 8372 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1636993656
transform 1 0 9476 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1636993656
transform 1 0 10580 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 25201
transform 1 0 11684 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 25201
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1636993656
transform 1 0 12420 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1636993656
transform 1 0 13524 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1636993656
transform 1 0 14628 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1636993656
transform 1 0 15732 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 25201
transform 1 0 16836 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 25201
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1636993656
transform 1 0 17572 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1636993656
transform 1 0 18676 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1636993656
transform 1 0 19780 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1636993656
transform 1 0 20884 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 25201
transform 1 0 21988 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 25201
transform 1 0 22540 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1636993656
transform 1 0 22724 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1636993656
transform 1 0 23828 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1636993656
transform 1 0 24932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1636993656
transform 1 0 26036 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 25201
transform 1 0 27140 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 25201
transform 1 0 27692 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1636993656
transform 1 0 27876 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1636993656
transform 1 0 28980 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1636993656
transform 1 0 30084 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1636993656
transform 1 0 31188 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 25201
transform 1 0 32292 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 25201
transform 1 0 32844 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1636993656
transform 1 0 33028 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1636993656
transform 1 0 34132 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1636993656
transform 1 0 35236 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1636993656
transform 1 0 36340 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 25201
transform 1 0 37444 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 25201
transform 1 0 37996 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1636993656
transform 1 0 38180 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1636993656
transform 1 0 39284 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1636993656
transform 1 0 40388 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1636993656
transform 1 0 41492 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 25201
transform 1 0 42596 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 25201
transform 1 0 43148 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1636993656
transform 1 0 43332 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1636993656
transform 1 0 44436 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1636993656
transform 1 0 45540 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1636993656
transform 1 0 46644 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 25201
transform 1 0 47748 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 25201
transform 1 0 48300 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1636993656
transform 1 0 48484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1636993656
transform 1 0 49588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1636993656
transform 1 0 50692 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1636993656
transform 1 0 51796 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 25201
transform 1 0 52900 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 25201
transform 1 0 53452 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1636993656
transform 1 0 53636 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1636993656
transform 1 0 54740 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1636993656
transform 1 0 55844 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1636993656
transform 1 0 56948 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 25201
transform 1 0 58052 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 25201
transform 1 0 58604 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1636993656
transform 1 0 58788 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1636993656
transform 1 0 59892 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1636993656
transform 1 0 60996 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1636993656
transform 1 0 62100 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 25201
transform 1 0 63204 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 25201
transform 1 0 63756 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_673
timestamp 1636993656
transform 1 0 63940 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_685
timestamp 1636993656
transform 1 0 65044 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1636993656
transform 1 0 66148 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_709
timestamp 1636993656
transform 1 0 67252 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 25201
transform 1 0 68356 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 25201
transform 1 0 68908 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_729
timestamp 1636993656
transform 1 0 69092 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_741
timestamp 1636993656
transform 1 0 70196 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_753
timestamp 1636993656
transform 1 0 71300 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_765
timestamp 1636993656
transform 1 0 72404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_777
timestamp 25201
transform 1 0 73508 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_783
timestamp 25201
transform 1 0 74060 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_785
timestamp 1636993656
transform 1 0 74244 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_797
timestamp 1636993656
transform 1 0 75348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_809
timestamp 1636993656
transform 1 0 76452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_821
timestamp 25201
transform 1 0 77556 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636993656
transform 1 0 2300 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636993656
transform 1 0 3404 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 25201
transform 1 0 4508 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636993656
transform 1 0 4692 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636993656
transform 1 0 5796 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636993656
transform 1 0 6900 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1636993656
transform 1 0 8004 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 25201
transform 1 0 9108 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 25201
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1636993656
transform 1 0 9844 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1636993656
transform 1 0 10948 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1636993656
transform 1 0 12052 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1636993656
transform 1 0 13156 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 25201
transform 1 0 14260 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 25201
transform 1 0 14812 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1636993656
transform 1 0 14996 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1636993656
transform 1 0 16100 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1636993656
transform 1 0 17204 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1636993656
transform 1 0 18308 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 25201
transform 1 0 19412 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 25201
transform 1 0 19964 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1636993656
transform 1 0 20148 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1636993656
transform 1 0 21252 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1636993656
transform 1 0 22356 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1636993656
transform 1 0 23460 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 25201
transform 1 0 24564 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 25201
transform 1 0 25116 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1636993656
transform 1 0 25300 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1636993656
transform 1 0 26404 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1636993656
transform 1 0 27508 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1636993656
transform 1 0 28612 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 25201
transform 1 0 29716 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 25201
transform 1 0 30268 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1636993656
transform 1 0 30452 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1636993656
transform 1 0 31556 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1636993656
transform 1 0 32660 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1636993656
transform 1 0 33764 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 25201
transform 1 0 34868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 25201
transform 1 0 35420 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1636993656
transform 1 0 35604 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1636993656
transform 1 0 36708 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1636993656
transform 1 0 37812 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1636993656
transform 1 0 38916 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 25201
transform 1 0 40020 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 25201
transform 1 0 40572 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1636993656
transform 1 0 40756 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1636993656
transform 1 0 41860 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1636993656
transform 1 0 42964 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1636993656
transform 1 0 44068 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 25201
transform 1 0 45172 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 25201
transform 1 0 45724 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1636993656
transform 1 0 45908 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1636993656
transform 1 0 47012 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1636993656
transform 1 0 48116 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1636993656
transform 1 0 49220 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 25201
transform 1 0 50324 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 25201
transform 1 0 50876 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1636993656
transform 1 0 51060 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1636993656
transform 1 0 52164 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1636993656
transform 1 0 53268 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1636993656
transform 1 0 54372 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 25201
transform 1 0 55476 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 25201
transform 1 0 56028 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1636993656
transform 1 0 56212 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1636993656
transform 1 0 57316 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1636993656
transform 1 0 58420 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_625
timestamp 1636993656
transform 1 0 59524 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 25201
transform 1 0 60628 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 25201
transform 1 0 61180 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1636993656
transform 1 0 61364 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1636993656
transform 1 0 62468 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_669
timestamp 1636993656
transform 1 0 63572 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_681
timestamp 1636993656
transform 1 0 64676 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 25201
transform 1 0 65780 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 25201
transform 1 0 66332 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1636993656
transform 1 0 66516 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1636993656
transform 1 0 67620 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_725
timestamp 1636993656
transform 1 0 68724 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_737
timestamp 1636993656
transform 1 0 69828 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_749
timestamp 25201
transform 1 0 70932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_755
timestamp 25201
transform 1 0 71484 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_757
timestamp 1636993656
transform 1 0 71668 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_769
timestamp 1636993656
transform 1 0 72772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_781
timestamp 1636993656
transform 1 0 73876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_793
timestamp 1636993656
transform 1 0 74980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_805
timestamp 25201
transform 1 0 76084 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_811
timestamp 25201
transform 1 0 76636 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_813
timestamp 25201
transform 1 0 76820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_821
timestamp 25201
transform 1 0 77556 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636993656
transform 1 0 2300 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636993656
transform 1 0 3404 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636993656
transform 1 0 4508 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636993656
transform 1 0 5612 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 25201
transform 1 0 6716 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 25201
transform 1 0 7084 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636993656
transform 1 0 7268 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1636993656
transform 1 0 8372 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1636993656
transform 1 0 9476 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1636993656
transform 1 0 10580 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 25201
transform 1 0 11684 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 25201
transform 1 0 12236 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1636993656
transform 1 0 12420 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1636993656
transform 1 0 13524 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1636993656
transform 1 0 14628 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1636993656
transform 1 0 15732 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 25201
transform 1 0 16836 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 25201
transform 1 0 17388 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1636993656
transform 1 0 17572 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1636993656
transform 1 0 18676 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1636993656
transform 1 0 19780 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1636993656
transform 1 0 20884 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 25201
transform 1 0 21988 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 25201
transform 1 0 22540 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1636993656
transform 1 0 22724 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1636993656
transform 1 0 23828 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1636993656
transform 1 0 24932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1636993656
transform 1 0 26036 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 25201
transform 1 0 27140 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 25201
transform 1 0 27692 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1636993656
transform 1 0 27876 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1636993656
transform 1 0 28980 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1636993656
transform 1 0 30084 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1636993656
transform 1 0 31188 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 25201
transform 1 0 32292 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 25201
transform 1 0 32844 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1636993656
transform 1 0 33028 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1636993656
transform 1 0 34132 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1636993656
transform 1 0 35236 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1636993656
transform 1 0 36340 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 25201
transform 1 0 37444 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 25201
transform 1 0 37996 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1636993656
transform 1 0 38180 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1636993656
transform 1 0 39284 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1636993656
transform 1 0 40388 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1636993656
transform 1 0 41492 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 25201
transform 1 0 42596 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 25201
transform 1 0 43148 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1636993656
transform 1 0 43332 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1636993656
transform 1 0 44436 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1636993656
transform 1 0 45540 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1636993656
transform 1 0 46644 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 25201
transform 1 0 47748 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 25201
transform 1 0 48300 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1636993656
transform 1 0 48484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1636993656
transform 1 0 49588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1636993656
transform 1 0 50692 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1636993656
transform 1 0 51796 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 25201
transform 1 0 52900 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 25201
transform 1 0 53452 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1636993656
transform 1 0 53636 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1636993656
transform 1 0 54740 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1636993656
transform 1 0 55844 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1636993656
transform 1 0 56948 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 25201
transform 1 0 58052 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 25201
transform 1 0 58604 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1636993656
transform 1 0 58788 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1636993656
transform 1 0 59892 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1636993656
transform 1 0 60996 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1636993656
transform 1 0 62100 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 25201
transform 1 0 63204 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 25201
transform 1 0 63756 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1636993656
transform 1 0 63940 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1636993656
transform 1 0 65044 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1636993656
transform 1 0 66148 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1636993656
transform 1 0 67252 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 25201
transform 1 0 68356 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 25201
transform 1 0 68908 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_729
timestamp 1636993656
transform 1 0 69092 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_741
timestamp 1636993656
transform 1 0 70196 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_753
timestamp 1636993656
transform 1 0 71300 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_765
timestamp 1636993656
transform 1 0 72404 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_777
timestamp 25201
transform 1 0 73508 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_783
timestamp 25201
transform 1 0 74060 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_785
timestamp 1636993656
transform 1 0 74244 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_797
timestamp 1636993656
transform 1 0 75348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_809
timestamp 1636993656
transform 1 0 76452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_821
timestamp 25201
transform 1 0 77556 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636993656
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636993656
transform 1 0 3404 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 25201
transform 1 0 4508 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636993656
transform 1 0 4692 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636993656
transform 1 0 5796 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636993656
transform 1 0 6900 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1636993656
transform 1 0 8004 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 25201
transform 1 0 9108 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 25201
transform 1 0 9660 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1636993656
transform 1 0 9844 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1636993656
transform 1 0 10948 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1636993656
transform 1 0 12052 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1636993656
transform 1 0 13156 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 25201
transform 1 0 14260 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 25201
transform 1 0 14812 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1636993656
transform 1 0 14996 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1636993656
transform 1 0 16100 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1636993656
transform 1 0 17204 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1636993656
transform 1 0 18308 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 25201
transform 1 0 19412 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 25201
transform 1 0 19964 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1636993656
transform 1 0 20148 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1636993656
transform 1 0 21252 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1636993656
transform 1 0 22356 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1636993656
transform 1 0 23460 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 25201
transform 1 0 24564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 25201
transform 1 0 25116 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1636993656
transform 1 0 25300 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1636993656
transform 1 0 26404 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1636993656
transform 1 0 27508 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1636993656
transform 1 0 28612 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 25201
transform 1 0 29716 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 25201
transform 1 0 30268 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1636993656
transform 1 0 30452 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1636993656
transform 1 0 31556 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1636993656
transform 1 0 32660 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1636993656
transform 1 0 33764 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 25201
transform 1 0 34868 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 25201
transform 1 0 35420 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1636993656
transform 1 0 35604 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1636993656
transform 1 0 36708 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1636993656
transform 1 0 37812 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1636993656
transform 1 0 38916 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 25201
transform 1 0 40020 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 25201
transform 1 0 40572 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1636993656
transform 1 0 40756 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1636993656
transform 1 0 41860 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1636993656
transform 1 0 42964 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1636993656
transform 1 0 44068 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 25201
transform 1 0 45172 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 25201
transform 1 0 45724 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1636993656
transform 1 0 45908 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1636993656
transform 1 0 47012 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1636993656
transform 1 0 48116 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1636993656
transform 1 0 49220 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 25201
transform 1 0 50324 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 25201
transform 1 0 50876 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1636993656
transform 1 0 51060 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1636993656
transform 1 0 52164 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1636993656
transform 1 0 53268 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1636993656
transform 1 0 54372 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 25201
transform 1 0 55476 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 25201
transform 1 0 56028 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1636993656
transform 1 0 56212 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1636993656
transform 1 0 57316 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1636993656
transform 1 0 58420 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1636993656
transform 1 0 59524 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 25201
transform 1 0 60628 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 25201
transform 1 0 61180 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1636993656
transform 1 0 61364 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1636993656
transform 1 0 62468 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1636993656
transform 1 0 63572 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1636993656
transform 1 0 64676 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 25201
transform 1 0 65780 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 25201
transform 1 0 66332 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1636993656
transform 1 0 66516 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1636993656
transform 1 0 67620 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_725
timestamp 1636993656
transform 1 0 68724 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_737
timestamp 1636993656
transform 1 0 69828 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_749
timestamp 25201
transform 1 0 70932 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_755
timestamp 25201
transform 1 0 71484 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_757
timestamp 1636993656
transform 1 0 71668 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_769
timestamp 1636993656
transform 1 0 72772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_781
timestamp 1636993656
transform 1 0 73876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_793
timestamp 1636993656
transform 1 0 74980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_805
timestamp 25201
transform 1 0 76084 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_811
timestamp 25201
transform 1 0 76636 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_813
timestamp 25201
transform 1 0 76820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_821
timestamp 25201
transform 1 0 77556 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636993656
transform 1 0 2300 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636993656
transform 1 0 3404 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636993656
transform 1 0 4508 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1636993656
transform 1 0 5612 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 25201
transform 1 0 6716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 25201
transform 1 0 7084 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636993656
transform 1 0 7268 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1636993656
transform 1 0 8372 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1636993656
transform 1 0 9476 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1636993656
transform 1 0 10580 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 25201
transform 1 0 11684 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 25201
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1636993656
transform 1 0 12420 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1636993656
transform 1 0 13524 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1636993656
transform 1 0 14628 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1636993656
transform 1 0 15732 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 25201
transform 1 0 16836 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 25201
transform 1 0 17388 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1636993656
transform 1 0 17572 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1636993656
transform 1 0 18676 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1636993656
transform 1 0 19780 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1636993656
transform 1 0 20884 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 25201
transform 1 0 21988 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 25201
transform 1 0 22540 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1636993656
transform 1 0 22724 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1636993656
transform 1 0 23828 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1636993656
transform 1 0 24932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1636993656
transform 1 0 26036 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 25201
transform 1 0 27140 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 25201
transform 1 0 27692 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1636993656
transform 1 0 27876 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1636993656
transform 1 0 28980 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1636993656
transform 1 0 30084 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1636993656
transform 1 0 31188 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 25201
transform 1 0 32292 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 25201
transform 1 0 32844 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1636993656
transform 1 0 33028 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1636993656
transform 1 0 34132 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1636993656
transform 1 0 35236 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1636993656
transform 1 0 36340 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 25201
transform 1 0 37444 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 25201
transform 1 0 37996 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1636993656
transform 1 0 38180 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1636993656
transform 1 0 39284 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1636993656
transform 1 0 40388 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1636993656
transform 1 0 41492 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 25201
transform 1 0 42596 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 25201
transform 1 0 43148 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1636993656
transform 1 0 43332 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1636993656
transform 1 0 44436 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1636993656
transform 1 0 45540 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1636993656
transform 1 0 46644 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 25201
transform 1 0 47748 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 25201
transform 1 0 48300 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1636993656
transform 1 0 48484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1636993656
transform 1 0 49588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1636993656
transform 1 0 50692 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1636993656
transform 1 0 51796 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 25201
transform 1 0 52900 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 25201
transform 1 0 53452 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1636993656
transform 1 0 53636 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1636993656
transform 1 0 54740 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1636993656
transform 1 0 55844 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1636993656
transform 1 0 56948 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 25201
transform 1 0 58052 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 25201
transform 1 0 58604 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1636993656
transform 1 0 58788 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1636993656
transform 1 0 59892 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1636993656
transform 1 0 60996 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1636993656
transform 1 0 62100 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 25201
transform 1 0 63204 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 25201
transform 1 0 63756 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1636993656
transform 1 0 63940 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1636993656
transform 1 0 65044 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1636993656
transform 1 0 66148 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1636993656
transform 1 0 67252 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 25201
transform 1 0 68356 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 25201
transform 1 0 68908 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_729
timestamp 1636993656
transform 1 0 69092 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_741
timestamp 1636993656
transform 1 0 70196 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_753
timestamp 1636993656
transform 1 0 71300 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_765
timestamp 1636993656
transform 1 0 72404 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_777
timestamp 25201
transform 1 0 73508 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_783
timestamp 25201
transform 1 0 74060 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_785
timestamp 1636993656
transform 1 0 74244 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_797
timestamp 1636993656
transform 1 0 75348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_809
timestamp 1636993656
transform 1 0 76452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_821
timestamp 25201
transform 1 0 77556 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636993656
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636993656
transform 1 0 3404 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 25201
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636993656
transform 1 0 4692 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636993656
transform 1 0 5796 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636993656
transform 1 0 6900 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1636993656
transform 1 0 8004 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 25201
transform 1 0 9108 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 25201
transform 1 0 9660 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1636993656
transform 1 0 9844 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1636993656
transform 1 0 10948 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1636993656
transform 1 0 12052 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1636993656
transform 1 0 13156 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 25201
transform 1 0 14260 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 25201
transform 1 0 14812 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1636993656
transform 1 0 14996 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1636993656
transform 1 0 16100 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1636993656
transform 1 0 17204 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1636993656
transform 1 0 18308 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 25201
transform 1 0 19412 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 25201
transform 1 0 19964 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1636993656
transform 1 0 20148 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1636993656
transform 1 0 21252 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1636993656
transform 1 0 22356 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1636993656
transform 1 0 23460 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 25201
transform 1 0 24564 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 25201
transform 1 0 25116 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1636993656
transform 1 0 25300 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1636993656
transform 1 0 26404 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1636993656
transform 1 0 27508 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1636993656
transform 1 0 28612 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 25201
transform 1 0 29716 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 25201
transform 1 0 30268 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1636993656
transform 1 0 30452 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1636993656
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1636993656
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1636993656
transform 1 0 33764 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 25201
transform 1 0 34868 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 25201
transform 1 0 35420 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1636993656
transform 1 0 35604 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1636993656
transform 1 0 36708 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1636993656
transform 1 0 37812 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1636993656
transform 1 0 38916 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 25201
transform 1 0 40020 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 25201
transform 1 0 40572 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1636993656
transform 1 0 40756 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1636993656
transform 1 0 41860 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1636993656
transform 1 0 42964 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1636993656
transform 1 0 44068 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 25201
transform 1 0 45172 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 25201
transform 1 0 45724 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1636993656
transform 1 0 45908 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1636993656
transform 1 0 47012 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1636993656
transform 1 0 48116 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1636993656
transform 1 0 49220 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 25201
transform 1 0 50324 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 25201
transform 1 0 50876 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1636993656
transform 1 0 51060 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1636993656
transform 1 0 52164 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1636993656
transform 1 0 53268 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1636993656
transform 1 0 54372 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 25201
transform 1 0 55476 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 25201
transform 1 0 56028 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1636993656
transform 1 0 56212 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1636993656
transform 1 0 57316 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1636993656
transform 1 0 58420 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1636993656
transform 1 0 59524 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 25201
transform 1 0 60628 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 25201
transform 1 0 61180 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1636993656
transform 1 0 61364 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1636993656
transform 1 0 62468 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1636993656
transform 1 0 63572 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1636993656
transform 1 0 64676 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 25201
transform 1 0 65780 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 25201
transform 1 0 66332 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1636993656
transform 1 0 66516 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1636993656
transform 1 0 67620 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_725
timestamp 1636993656
transform 1 0 68724 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_737
timestamp 1636993656
transform 1 0 69828 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_749
timestamp 25201
transform 1 0 70932 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_755
timestamp 25201
transform 1 0 71484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_757
timestamp 1636993656
transform 1 0 71668 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_769
timestamp 1636993656
transform 1 0 72772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_781
timestamp 1636993656
transform 1 0 73876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_793
timestamp 1636993656
transform 1 0 74980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_805
timestamp 25201
transform 1 0 76084 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_811
timestamp 25201
transform 1 0 76636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_813
timestamp 25201
transform 1 0 76820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_821
timestamp 25201
transform 1 0 77556 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636993656
transform 1 0 2300 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636993656
transform 1 0 3404 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636993656
transform 1 0 4508 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1636993656
transform 1 0 5612 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 25201
transform 1 0 6716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 25201
transform 1 0 7084 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636993656
transform 1 0 7268 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1636993656
transform 1 0 8372 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1636993656
transform 1 0 9476 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1636993656
transform 1 0 10580 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 25201
transform 1 0 11684 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 25201
transform 1 0 12236 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1636993656
transform 1 0 12420 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1636993656
transform 1 0 13524 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1636993656
transform 1 0 14628 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1636993656
transform 1 0 15732 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 25201
transform 1 0 16836 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 25201
transform 1 0 17388 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1636993656
transform 1 0 17572 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1636993656
transform 1 0 18676 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1636993656
transform 1 0 19780 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1636993656
transform 1 0 20884 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 25201
transform 1 0 21988 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 25201
transform 1 0 22540 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1636993656
transform 1 0 22724 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1636993656
transform 1 0 23828 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1636993656
transform 1 0 24932 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1636993656
transform 1 0 26036 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 25201
transform 1 0 27140 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 25201
transform 1 0 27692 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1636993656
transform 1 0 27876 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1636993656
transform 1 0 28980 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1636993656
transform 1 0 30084 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1636993656
transform 1 0 31188 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 25201
transform 1 0 32292 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 25201
transform 1 0 32844 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1636993656
transform 1 0 33028 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1636993656
transform 1 0 34132 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1636993656
transform 1 0 35236 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1636993656
transform 1 0 36340 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 25201
transform 1 0 37444 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 25201
transform 1 0 37996 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1636993656
transform 1 0 38180 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1636993656
transform 1 0 39284 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1636993656
transform 1 0 40388 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1636993656
transform 1 0 41492 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 25201
transform 1 0 42596 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 25201
transform 1 0 43148 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1636993656
transform 1 0 43332 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1636993656
transform 1 0 44436 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1636993656
transform 1 0 45540 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1636993656
transform 1 0 46644 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 25201
transform 1 0 47748 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 25201
transform 1 0 48300 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1636993656
transform 1 0 48484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1636993656
transform 1 0 49588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1636993656
transform 1 0 50692 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1636993656
transform 1 0 51796 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 25201
transform 1 0 52900 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 25201
transform 1 0 53452 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1636993656
transform 1 0 53636 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1636993656
transform 1 0 54740 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1636993656
transform 1 0 55844 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1636993656
transform 1 0 56948 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 25201
transform 1 0 58052 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 25201
transform 1 0 58604 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1636993656
transform 1 0 58788 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1636993656
transform 1 0 59892 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1636993656
transform 1 0 60996 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1636993656
transform 1 0 62100 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 25201
transform 1 0 63204 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 25201
transform 1 0 63756 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1636993656
transform 1 0 63940 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1636993656
transform 1 0 65044 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1636993656
transform 1 0 66148 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1636993656
transform 1 0 67252 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 25201
transform 1 0 68356 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 25201
transform 1 0 68908 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_729
timestamp 1636993656
transform 1 0 69092 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_741
timestamp 1636993656
transform 1 0 70196 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_753
timestamp 1636993656
transform 1 0 71300 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_765
timestamp 1636993656
transform 1 0 72404 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_777
timestamp 25201
transform 1 0 73508 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_783
timestamp 25201
transform 1 0 74060 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_785
timestamp 1636993656
transform 1 0 74244 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_797
timestamp 1636993656
transform 1 0 75348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_809
timestamp 1636993656
transform 1 0 76452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_821
timestamp 25201
transform 1 0 77556 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636993656
transform 1 0 2300 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636993656
transform 1 0 3404 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 25201
transform 1 0 4508 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636993656
transform 1 0 4692 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1636993656
transform 1 0 5796 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1636993656
transform 1 0 6900 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1636993656
transform 1 0 8004 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 25201
transform 1 0 9108 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 25201
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1636993656
transform 1 0 9844 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1636993656
transform 1 0 10948 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1636993656
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1636993656
transform 1 0 13156 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 25201
transform 1 0 14260 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 25201
transform 1 0 14812 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1636993656
transform 1 0 14996 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1636993656
transform 1 0 16100 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1636993656
transform 1 0 17204 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1636993656
transform 1 0 18308 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 25201
transform 1 0 19412 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 25201
transform 1 0 19964 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1636993656
transform 1 0 20148 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1636993656
transform 1 0 21252 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1636993656
transform 1 0 22356 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1636993656
transform 1 0 23460 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 25201
transform 1 0 24564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 25201
transform 1 0 25116 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1636993656
transform 1 0 25300 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1636993656
transform 1 0 26404 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1636993656
transform 1 0 27508 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1636993656
transform 1 0 28612 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 25201
transform 1 0 29716 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 25201
transform 1 0 30268 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1636993656
transform 1 0 30452 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1636993656
transform 1 0 31556 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1636993656
transform 1 0 32660 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1636993656
transform 1 0 33764 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 25201
transform 1 0 34868 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 25201
transform 1 0 35420 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1636993656
transform 1 0 35604 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1636993656
transform 1 0 36708 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1636993656
transform 1 0 37812 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1636993656
transform 1 0 38916 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 25201
transform 1 0 40020 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 25201
transform 1 0 40572 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1636993656
transform 1 0 40756 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1636993656
transform 1 0 41860 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1636993656
transform 1 0 42964 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1636993656
transform 1 0 44068 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 25201
transform 1 0 45172 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 25201
transform 1 0 45724 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1636993656
transform 1 0 45908 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1636993656
transform 1 0 47012 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1636993656
transform 1 0 48116 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1636993656
transform 1 0 49220 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 25201
transform 1 0 50324 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 25201
transform 1 0 50876 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1636993656
transform 1 0 51060 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1636993656
transform 1 0 52164 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1636993656
transform 1 0 53268 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1636993656
transform 1 0 54372 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 25201
transform 1 0 55476 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 25201
transform 1 0 56028 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1636993656
transform 1 0 56212 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1636993656
transform 1 0 57316 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1636993656
transform 1 0 58420 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1636993656
transform 1 0 59524 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 25201
transform 1 0 60628 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 25201
transform 1 0 61180 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1636993656
transform 1 0 61364 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1636993656
transform 1 0 62468 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1636993656
transform 1 0 63572 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1636993656
transform 1 0 64676 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 25201
transform 1 0 65780 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 25201
transform 1 0 66332 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1636993656
transform 1 0 66516 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1636993656
transform 1 0 67620 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_725
timestamp 1636993656
transform 1 0 68724 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_737
timestamp 1636993656
transform 1 0 69828 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_749
timestamp 25201
transform 1 0 70932 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_755
timestamp 25201
transform 1 0 71484 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_757
timestamp 1636993656
transform 1 0 71668 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_769
timestamp 1636993656
transform 1 0 72772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_781
timestamp 1636993656
transform 1 0 73876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_793
timestamp 1636993656
transform 1 0 74980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_805
timestamp 25201
transform 1 0 76084 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_811
timestamp 25201
transform 1 0 76636 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_813
timestamp 25201
transform 1 0 76820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_821
timestamp 25201
transform 1 0 77556 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636993656
transform 1 0 2300 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636993656
transform 1 0 3404 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1636993656
transform 1 0 4508 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1636993656
transform 1 0 5612 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 25201
transform 1 0 6716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 25201
transform 1 0 7084 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636993656
transform 1 0 7268 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1636993656
transform 1 0 8372 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1636993656
transform 1 0 9476 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1636993656
transform 1 0 10580 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 25201
transform 1 0 11684 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 25201
transform 1 0 12236 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1636993656
transform 1 0 12420 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1636993656
transform 1 0 13524 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1636993656
transform 1 0 14628 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1636993656
transform 1 0 15732 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 25201
transform 1 0 16836 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 25201
transform 1 0 17388 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1636993656
transform 1 0 17572 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1636993656
transform 1 0 18676 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1636993656
transform 1 0 19780 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1636993656
transform 1 0 20884 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 25201
transform 1 0 21988 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 25201
transform 1 0 22540 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1636993656
transform 1 0 22724 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1636993656
transform 1 0 23828 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1636993656
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1636993656
transform 1 0 26036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 25201
transform 1 0 27140 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 25201
transform 1 0 27692 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1636993656
transform 1 0 27876 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1636993656
transform 1 0 28980 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1636993656
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1636993656
transform 1 0 31188 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 25201
transform 1 0 32292 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 25201
transform 1 0 32844 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1636993656
transform 1 0 33028 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1636993656
transform 1 0 34132 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1636993656
transform 1 0 35236 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1636993656
transform 1 0 36340 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 25201
transform 1 0 37444 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 25201
transform 1 0 37996 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1636993656
transform 1 0 38180 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1636993656
transform 1 0 39284 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1636993656
transform 1 0 40388 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1636993656
transform 1 0 41492 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 25201
transform 1 0 42596 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 25201
transform 1 0 43148 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1636993656
transform 1 0 43332 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1636993656
transform 1 0 44436 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1636993656
transform 1 0 45540 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1636993656
transform 1 0 46644 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 25201
transform 1 0 47748 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 25201
transform 1 0 48300 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1636993656
transform 1 0 48484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1636993656
transform 1 0 49588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1636993656
transform 1 0 50692 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1636993656
transform 1 0 51796 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 25201
transform 1 0 52900 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 25201
transform 1 0 53452 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1636993656
transform 1 0 53636 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1636993656
transform 1 0 54740 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1636993656
transform 1 0 55844 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1636993656
transform 1 0 56948 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 25201
transform 1 0 58052 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 25201
transform 1 0 58604 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1636993656
transform 1 0 58788 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1636993656
transform 1 0 59892 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1636993656
transform 1 0 60996 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1636993656
transform 1 0 62100 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 25201
transform 1 0 63204 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 25201
transform 1 0 63756 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1636993656
transform 1 0 63940 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1636993656
transform 1 0 65044 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1636993656
transform 1 0 66148 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1636993656
transform 1 0 67252 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 25201
transform 1 0 68356 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 25201
transform 1 0 68908 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_729
timestamp 1636993656
transform 1 0 69092 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_741
timestamp 1636993656
transform 1 0 70196 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_753
timestamp 1636993656
transform 1 0 71300 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_765
timestamp 1636993656
transform 1 0 72404 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_777
timestamp 25201
transform 1 0 73508 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_783
timestamp 25201
transform 1 0 74060 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_785
timestamp 1636993656
transform 1 0 74244 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_797
timestamp 1636993656
transform 1 0 75348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_809
timestamp 1636993656
transform 1 0 76452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_821
timestamp 25201
transform 1 0 77556 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636993656
transform 1 0 2300 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636993656
transform 1 0 3404 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 25201
transform 1 0 4508 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636993656
transform 1 0 4692 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1636993656
transform 1 0 5796 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1636993656
transform 1 0 6900 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1636993656
transform 1 0 8004 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 25201
transform 1 0 9108 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 25201
transform 1 0 9660 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1636993656
transform 1 0 9844 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1636993656
transform 1 0 10948 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1636993656
transform 1 0 12052 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1636993656
transform 1 0 13156 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 25201
transform 1 0 14260 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 25201
transform 1 0 14812 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1636993656
transform 1 0 14996 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1636993656
transform 1 0 16100 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1636993656
transform 1 0 17204 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1636993656
transform 1 0 18308 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 25201
transform 1 0 19412 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 25201
transform 1 0 19964 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1636993656
transform 1 0 20148 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1636993656
transform 1 0 21252 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1636993656
transform 1 0 22356 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1636993656
transform 1 0 23460 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 25201
transform 1 0 24564 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 25201
transform 1 0 25116 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1636993656
transform 1 0 25300 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1636993656
transform 1 0 26404 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1636993656
transform 1 0 27508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1636993656
transform 1 0 28612 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 25201
transform 1 0 29716 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 25201
transform 1 0 30268 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1636993656
transform 1 0 30452 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1636993656
transform 1 0 31556 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1636993656
transform 1 0 32660 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1636993656
transform 1 0 33764 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 25201
transform 1 0 34868 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 25201
transform 1 0 35420 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1636993656
transform 1 0 35604 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1636993656
transform 1 0 36708 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1636993656
transform 1 0 37812 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1636993656
transform 1 0 38916 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 25201
transform 1 0 40020 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 25201
transform 1 0 40572 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1636993656
transform 1 0 40756 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1636993656
transform 1 0 41860 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1636993656
transform 1 0 42964 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1636993656
transform 1 0 44068 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 25201
transform 1 0 45172 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 25201
transform 1 0 45724 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1636993656
transform 1 0 45908 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1636993656
transform 1 0 47012 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1636993656
transform 1 0 48116 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1636993656
transform 1 0 49220 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 25201
transform 1 0 50324 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 25201
transform 1 0 50876 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1636993656
transform 1 0 51060 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1636993656
transform 1 0 52164 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1636993656
transform 1 0 53268 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1636993656
transform 1 0 54372 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 25201
transform 1 0 55476 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 25201
transform 1 0 56028 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1636993656
transform 1 0 56212 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1636993656
transform 1 0 57316 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1636993656
transform 1 0 58420 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1636993656
transform 1 0 59524 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 25201
transform 1 0 60628 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 25201
transform 1 0 61180 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1636993656
transform 1 0 61364 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1636993656
transform 1 0 62468 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1636993656
transform 1 0 63572 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1636993656
transform 1 0 64676 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 25201
transform 1 0 65780 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 25201
transform 1 0 66332 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1636993656
transform 1 0 66516 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1636993656
transform 1 0 67620 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_725
timestamp 1636993656
transform 1 0 68724 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_737
timestamp 1636993656
transform 1 0 69828 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_749
timestamp 25201
transform 1 0 70932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_755
timestamp 25201
transform 1 0 71484 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_757
timestamp 1636993656
transform 1 0 71668 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_769
timestamp 1636993656
transform 1 0 72772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_781
timestamp 1636993656
transform 1 0 73876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_793
timestamp 1636993656
transform 1 0 74980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_805
timestamp 25201
transform 1 0 76084 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_811
timestamp 25201
transform 1 0 76636 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_813
timestamp 25201
transform 1 0 76820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_821
timestamp 25201
transform 1 0 77556 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1636993656
transform 1 0 2300 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1636993656
transform 1 0 3404 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1636993656
transform 1 0 4508 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1636993656
transform 1 0 5612 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 25201
transform 1 0 6716 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 25201
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636993656
transform 1 0 7268 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1636993656
transform 1 0 8372 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1636993656
transform 1 0 9476 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1636993656
transform 1 0 10580 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 25201
transform 1 0 11684 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 25201
transform 1 0 12236 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1636993656
transform 1 0 12420 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1636993656
transform 1 0 13524 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1636993656
transform 1 0 14628 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1636993656
transform 1 0 15732 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 25201
transform 1 0 16836 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 25201
transform 1 0 17388 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1636993656
transform 1 0 17572 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1636993656
transform 1 0 18676 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1636993656
transform 1 0 19780 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1636993656
transform 1 0 20884 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 25201
transform 1 0 21988 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 25201
transform 1 0 22540 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1636993656
transform 1 0 22724 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1636993656
transform 1 0 23828 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1636993656
transform 1 0 24932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1636993656
transform 1 0 26036 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 25201
transform 1 0 27140 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 25201
transform 1 0 27692 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1636993656
transform 1 0 27876 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1636993656
transform 1 0 28980 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1636993656
transform 1 0 30084 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1636993656
transform 1 0 31188 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 25201
transform 1 0 32292 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 25201
transform 1 0 32844 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1636993656
transform 1 0 33028 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1636993656
transform 1 0 34132 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1636993656
transform 1 0 35236 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1636993656
transform 1 0 36340 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 25201
transform 1 0 37444 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 25201
transform 1 0 37996 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1636993656
transform 1 0 38180 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1636993656
transform 1 0 39284 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1636993656
transform 1 0 40388 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1636993656
transform 1 0 41492 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 25201
transform 1 0 42596 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 25201
transform 1 0 43148 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1636993656
transform 1 0 43332 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1636993656
transform 1 0 44436 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1636993656
transform 1 0 45540 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1636993656
transform 1 0 46644 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 25201
transform 1 0 47748 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 25201
transform 1 0 48300 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1636993656
transform 1 0 48484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1636993656
transform 1 0 49588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1636993656
transform 1 0 50692 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1636993656
transform 1 0 51796 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 25201
transform 1 0 52900 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 25201
transform 1 0 53452 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1636993656
transform 1 0 53636 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1636993656
transform 1 0 54740 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1636993656
transform 1 0 55844 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1636993656
transform 1 0 56948 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 25201
transform 1 0 58052 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 25201
transform 1 0 58604 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1636993656
transform 1 0 58788 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1636993656
transform 1 0 59892 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1636993656
transform 1 0 60996 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1636993656
transform 1 0 62100 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 25201
transform 1 0 63204 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 25201
transform 1 0 63756 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1636993656
transform 1 0 63940 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1636993656
transform 1 0 65044 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1636993656
transform 1 0 66148 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1636993656
transform 1 0 67252 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 25201
transform 1 0 68356 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 25201
transform 1 0 68908 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_729
timestamp 1636993656
transform 1 0 69092 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_741
timestamp 1636993656
transform 1 0 70196 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_753
timestamp 1636993656
transform 1 0 71300 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_765
timestamp 1636993656
transform 1 0 72404 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_777
timestamp 25201
transform 1 0 73508 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_783
timestamp 25201
transform 1 0 74060 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_785
timestamp 1636993656
transform 1 0 74244 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_797
timestamp 1636993656
transform 1 0 75348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_809
timestamp 1636993656
transform 1 0 76452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_821
timestamp 25201
transform 1 0 77556 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636993656
transform 1 0 2300 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636993656
transform 1 0 3404 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 25201
transform 1 0 4508 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636993656
transform 1 0 4692 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636993656
transform 1 0 5796 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636993656
transform 1 0 6900 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1636993656
transform 1 0 8004 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 25201
transform 1 0 9108 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 25201
transform 1 0 9660 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1636993656
transform 1 0 9844 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1636993656
transform 1 0 10948 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1636993656
transform 1 0 12052 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1636993656
transform 1 0 13156 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 25201
transform 1 0 14260 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 25201
transform 1 0 14812 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1636993656
transform 1 0 14996 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1636993656
transform 1 0 16100 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1636993656
transform 1 0 17204 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1636993656
transform 1 0 18308 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 25201
transform 1 0 19412 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 25201
transform 1 0 19964 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1636993656
transform 1 0 20148 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1636993656
transform 1 0 21252 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1636993656
transform 1 0 22356 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1636993656
transform 1 0 23460 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 25201
transform 1 0 24564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 25201
transform 1 0 25116 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1636993656
transform 1 0 25300 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1636993656
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1636993656
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1636993656
transform 1 0 28612 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 25201
transform 1 0 29716 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 25201
transform 1 0 30268 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1636993656
transform 1 0 30452 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1636993656
transform 1 0 31556 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1636993656
transform 1 0 32660 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1636993656
transform 1 0 33764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 25201
transform 1 0 34868 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 25201
transform 1 0 35420 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1636993656
transform 1 0 35604 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1636993656
transform 1 0 36708 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1636993656
transform 1 0 37812 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1636993656
transform 1 0 38916 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 25201
transform 1 0 40020 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 25201
transform 1 0 40572 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1636993656
transform 1 0 40756 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1636993656
transform 1 0 41860 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1636993656
transform 1 0 42964 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1636993656
transform 1 0 44068 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 25201
transform 1 0 45172 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 25201
transform 1 0 45724 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1636993656
transform 1 0 45908 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1636993656
transform 1 0 47012 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1636993656
transform 1 0 48116 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1636993656
transform 1 0 49220 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 25201
transform 1 0 50324 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 25201
transform 1 0 50876 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1636993656
transform 1 0 51060 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1636993656
transform 1 0 52164 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1636993656
transform 1 0 53268 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1636993656
transform 1 0 54372 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 25201
transform 1 0 55476 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 25201
transform 1 0 56028 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1636993656
transform 1 0 56212 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1636993656
transform 1 0 57316 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1636993656
transform 1 0 58420 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1636993656
transform 1 0 59524 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 25201
transform 1 0 60628 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 25201
transform 1 0 61180 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1636993656
transform 1 0 61364 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1636993656
transform 1 0 62468 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1636993656
transform 1 0 63572 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1636993656
transform 1 0 64676 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 25201
transform 1 0 65780 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 25201
transform 1 0 66332 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1636993656
transform 1 0 66516 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1636993656
transform 1 0 67620 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_725
timestamp 1636993656
transform 1 0 68724 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_737
timestamp 1636993656
transform 1 0 69828 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_749
timestamp 25201
transform 1 0 70932 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_755
timestamp 25201
transform 1 0 71484 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_757
timestamp 1636993656
transform 1 0 71668 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_769
timestamp 1636993656
transform 1 0 72772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_781
timestamp 1636993656
transform 1 0 73876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_793
timestamp 1636993656
transform 1 0 74980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_805
timestamp 25201
transform 1 0 76084 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_811
timestamp 25201
transform 1 0 76636 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_813
timestamp 25201
transform 1 0 76820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_821
timestamp 25201
transform 1 0 77556 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636993656
transform 1 0 2300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636993656
transform 1 0 3404 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636993656
transform 1 0 4508 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1636993656
transform 1 0 5612 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 25201
transform 1 0 6716 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 25201
transform 1 0 7084 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636993656
transform 1 0 7268 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1636993656
transform 1 0 8372 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1636993656
transform 1 0 9476 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1636993656
transform 1 0 10580 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 25201
transform 1 0 11684 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 25201
transform 1 0 12236 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1636993656
transform 1 0 12420 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1636993656
transform 1 0 13524 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1636993656
transform 1 0 14628 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1636993656
transform 1 0 15732 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 25201
transform 1 0 16836 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 25201
transform 1 0 17388 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1636993656
transform 1 0 17572 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1636993656
transform 1 0 18676 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1636993656
transform 1 0 19780 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1636993656
transform 1 0 20884 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 25201
transform 1 0 21988 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 25201
transform 1 0 22540 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1636993656
transform 1 0 22724 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1636993656
transform 1 0 23828 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1636993656
transform 1 0 24932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1636993656
transform 1 0 26036 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 25201
transform 1 0 27140 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 25201
transform 1 0 27692 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1636993656
transform 1 0 27876 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1636993656
transform 1 0 28980 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1636993656
transform 1 0 30084 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1636993656
transform 1 0 31188 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 25201
transform 1 0 32292 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 25201
transform 1 0 32844 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1636993656
transform 1 0 33028 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1636993656
transform 1 0 34132 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1636993656
transform 1 0 35236 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1636993656
transform 1 0 36340 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 25201
transform 1 0 37444 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 25201
transform 1 0 37996 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1636993656
transform 1 0 38180 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1636993656
transform 1 0 39284 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1636993656
transform 1 0 40388 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1636993656
transform 1 0 41492 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 25201
transform 1 0 42596 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 25201
transform 1 0 43148 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1636993656
transform 1 0 43332 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1636993656
transform 1 0 44436 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1636993656
transform 1 0 45540 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1636993656
transform 1 0 46644 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 25201
transform 1 0 47748 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 25201
transform 1 0 48300 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1636993656
transform 1 0 48484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1636993656
transform 1 0 49588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1636993656
transform 1 0 50692 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1636993656
transform 1 0 51796 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 25201
transform 1 0 52900 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 25201
transform 1 0 53452 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1636993656
transform 1 0 53636 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1636993656
transform 1 0 54740 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1636993656
transform 1 0 55844 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1636993656
transform 1 0 56948 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 25201
transform 1 0 58052 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 25201
transform 1 0 58604 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1636993656
transform 1 0 58788 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1636993656
transform 1 0 59892 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1636993656
transform 1 0 60996 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1636993656
transform 1 0 62100 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 25201
transform 1 0 63204 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 25201
transform 1 0 63756 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1636993656
transform 1 0 63940 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1636993656
transform 1 0 65044 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1636993656
transform 1 0 66148 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1636993656
transform 1 0 67252 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 25201
transform 1 0 68356 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 25201
transform 1 0 68908 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_729
timestamp 1636993656
transform 1 0 69092 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_741
timestamp 1636993656
transform 1 0 70196 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_753
timestamp 1636993656
transform 1 0 71300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_765
timestamp 1636993656
transform 1 0 72404 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_777
timestamp 25201
transform 1 0 73508 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_783
timestamp 25201
transform 1 0 74060 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_785
timestamp 1636993656
transform 1 0 74244 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_797
timestamp 1636993656
transform 1 0 75348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_809
timestamp 1636993656
transform 1 0 76452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_821
timestamp 25201
transform 1 0 77556 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636993656
transform 1 0 2300 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636993656
transform 1 0 3404 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 25201
transform 1 0 4508 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636993656
transform 1 0 4692 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636993656
transform 1 0 5796 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1636993656
transform 1 0 6900 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1636993656
transform 1 0 8004 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 25201
transform 1 0 9108 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 25201
transform 1 0 9660 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1636993656
transform 1 0 9844 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1636993656
transform 1 0 10948 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1636993656
transform 1 0 12052 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1636993656
transform 1 0 13156 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 25201
transform 1 0 14260 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 25201
transform 1 0 14812 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1636993656
transform 1 0 14996 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1636993656
transform 1 0 16100 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1636993656
transform 1 0 17204 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1636993656
transform 1 0 18308 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 25201
transform 1 0 19412 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 25201
transform 1 0 19964 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1636993656
transform 1 0 20148 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1636993656
transform 1 0 21252 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1636993656
transform 1 0 22356 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1636993656
transform 1 0 23460 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 25201
transform 1 0 24564 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 25201
transform 1 0 25116 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1636993656
transform 1 0 25300 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1636993656
transform 1 0 26404 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1636993656
transform 1 0 27508 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1636993656
transform 1 0 28612 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 25201
transform 1 0 29716 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 25201
transform 1 0 30268 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1636993656
transform 1 0 30452 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1636993656
transform 1 0 31556 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1636993656
transform 1 0 32660 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1636993656
transform 1 0 33764 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 25201
transform 1 0 34868 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 25201
transform 1 0 35420 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1636993656
transform 1 0 35604 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1636993656
transform 1 0 36708 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1636993656
transform 1 0 37812 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1636993656
transform 1 0 38916 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 25201
transform 1 0 40020 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 25201
transform 1 0 40572 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1636993656
transform 1 0 40756 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1636993656
transform 1 0 41860 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1636993656
transform 1 0 42964 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1636993656
transform 1 0 44068 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 25201
transform 1 0 45172 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 25201
transform 1 0 45724 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1636993656
transform 1 0 45908 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1636993656
transform 1 0 47012 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1636993656
transform 1 0 48116 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1636993656
transform 1 0 49220 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 25201
transform 1 0 50324 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 25201
transform 1 0 50876 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1636993656
transform 1 0 51060 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1636993656
transform 1 0 52164 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1636993656
transform 1 0 53268 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1636993656
transform 1 0 54372 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 25201
transform 1 0 55476 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 25201
transform 1 0 56028 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1636993656
transform 1 0 56212 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1636993656
transform 1 0 57316 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1636993656
transform 1 0 58420 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1636993656
transform 1 0 59524 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 25201
transform 1 0 60628 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 25201
transform 1 0 61180 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1636993656
transform 1 0 61364 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1636993656
transform 1 0 62468 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1636993656
transform 1 0 63572 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1636993656
transform 1 0 64676 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 25201
transform 1 0 65780 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 25201
transform 1 0 66332 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1636993656
transform 1 0 66516 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1636993656
transform 1 0 67620 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_725
timestamp 1636993656
transform 1 0 68724 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_737
timestamp 1636993656
transform 1 0 69828 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_749
timestamp 25201
transform 1 0 70932 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_755
timestamp 25201
transform 1 0 71484 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_757
timestamp 1636993656
transform 1 0 71668 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_769
timestamp 1636993656
transform 1 0 72772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_781
timestamp 1636993656
transform 1 0 73876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_793
timestamp 1636993656
transform 1 0 74980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_805
timestamp 25201
transform 1 0 76084 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_811
timestamp 25201
transform 1 0 76636 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_813
timestamp 25201
transform 1 0 76820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_821
timestamp 25201
transform 1 0 77556 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636993656
transform 1 0 2300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636993656
transform 1 0 3404 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1636993656
transform 1 0 4508 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1636993656
transform 1 0 5612 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 25201
transform 1 0 6716 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 25201
transform 1 0 7084 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636993656
transform 1 0 7268 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1636993656
transform 1 0 8372 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1636993656
transform 1 0 9476 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1636993656
transform 1 0 10580 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 25201
transform 1 0 11684 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 25201
transform 1 0 12236 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1636993656
transform 1 0 12420 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1636993656
transform 1 0 13524 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1636993656
transform 1 0 14628 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1636993656
transform 1 0 15732 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 25201
transform 1 0 16836 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 25201
transform 1 0 17388 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1636993656
transform 1 0 17572 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1636993656
transform 1 0 18676 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1636993656
transform 1 0 19780 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1636993656
transform 1 0 20884 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 25201
transform 1 0 21988 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 25201
transform 1 0 22540 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1636993656
transform 1 0 22724 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1636993656
transform 1 0 23828 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1636993656
transform 1 0 24932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1636993656
transform 1 0 26036 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 25201
transform 1 0 27140 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 25201
transform 1 0 27692 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1636993656
transform 1 0 27876 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1636993656
transform 1 0 28980 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1636993656
transform 1 0 30084 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1636993656
transform 1 0 31188 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 25201
transform 1 0 32292 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 25201
transform 1 0 32844 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1636993656
transform 1 0 33028 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1636993656
transform 1 0 34132 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1636993656
transform 1 0 35236 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1636993656
transform 1 0 36340 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 25201
transform 1 0 37444 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 25201
transform 1 0 37996 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1636993656
transform 1 0 38180 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1636993656
transform 1 0 39284 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1636993656
transform 1 0 40388 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1636993656
transform 1 0 41492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 25201
transform 1 0 42596 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 25201
transform 1 0 43148 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1636993656
transform 1 0 43332 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1636993656
transform 1 0 44436 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1636993656
transform 1 0 45540 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1636993656
transform 1 0 46644 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 25201
transform 1 0 47748 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 25201
transform 1 0 48300 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1636993656
transform 1 0 48484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1636993656
transform 1 0 49588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1636993656
transform 1 0 50692 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1636993656
transform 1 0 51796 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 25201
transform 1 0 52900 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 25201
transform 1 0 53452 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1636993656
transform 1 0 53636 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1636993656
transform 1 0 54740 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1636993656
transform 1 0 55844 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1636993656
transform 1 0 56948 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 25201
transform 1 0 58052 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 25201
transform 1 0 58604 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1636993656
transform 1 0 58788 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1636993656
transform 1 0 59892 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1636993656
transform 1 0 60996 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1636993656
transform 1 0 62100 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 25201
transform 1 0 63204 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 25201
transform 1 0 63756 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1636993656
transform 1 0 63940 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1636993656
transform 1 0 65044 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1636993656
transform 1 0 66148 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1636993656
transform 1 0 67252 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 25201
transform 1 0 68356 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 25201
transform 1 0 68908 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_729
timestamp 1636993656
transform 1 0 69092 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_741
timestamp 1636993656
transform 1 0 70196 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_753
timestamp 1636993656
transform 1 0 71300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_765
timestamp 1636993656
transform 1 0 72404 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_777
timestamp 25201
transform 1 0 73508 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_783
timestamp 25201
transform 1 0 74060 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_785
timestamp 1636993656
transform 1 0 74244 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_797
timestamp 1636993656
transform 1 0 75348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_809
timestamp 1636993656
transform 1 0 76452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_821
timestamp 25201
transform 1 0 77556 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636993656
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636993656
transform 1 0 3404 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 25201
transform 1 0 4508 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636993656
transform 1 0 4692 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636993656
transform 1 0 5796 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636993656
transform 1 0 6900 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1636993656
transform 1 0 8004 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 25201
transform 1 0 9108 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 25201
transform 1 0 9660 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1636993656
transform 1 0 9844 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1636993656
transform 1 0 10948 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1636993656
transform 1 0 12052 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1636993656
transform 1 0 13156 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 25201
transform 1 0 14260 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 25201
transform 1 0 14812 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1636993656
transform 1 0 14996 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1636993656
transform 1 0 16100 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1636993656
transform 1 0 17204 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1636993656
transform 1 0 18308 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 25201
transform 1 0 19412 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 25201
transform 1 0 19964 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1636993656
transform 1 0 20148 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1636993656
transform 1 0 21252 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1636993656
transform 1 0 22356 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1636993656
transform 1 0 23460 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 25201
transform 1 0 24564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 25201
transform 1 0 25116 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1636993656
transform 1 0 25300 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1636993656
transform 1 0 26404 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1636993656
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1636993656
transform 1 0 28612 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 25201
transform 1 0 29716 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 25201
transform 1 0 30268 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1636993656
transform 1 0 30452 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1636993656
transform 1 0 31556 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1636993656
transform 1 0 32660 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1636993656
transform 1 0 33764 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 25201
transform 1 0 34868 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 25201
transform 1 0 35420 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1636993656
transform 1 0 35604 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1636993656
transform 1 0 36708 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1636993656
transform 1 0 37812 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1636993656
transform 1 0 38916 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 25201
transform 1 0 40020 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 25201
transform 1 0 40572 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1636993656
transform 1 0 40756 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1636993656
transform 1 0 41860 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1636993656
transform 1 0 42964 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1636993656
transform 1 0 44068 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 25201
transform 1 0 45172 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 25201
transform 1 0 45724 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1636993656
transform 1 0 45908 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1636993656
transform 1 0 47012 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1636993656
transform 1 0 48116 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1636993656
transform 1 0 49220 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 25201
transform 1 0 50324 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 25201
transform 1 0 50876 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1636993656
transform 1 0 51060 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1636993656
transform 1 0 52164 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1636993656
transform 1 0 53268 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1636993656
transform 1 0 54372 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 25201
transform 1 0 55476 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 25201
transform 1 0 56028 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1636993656
transform 1 0 56212 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1636993656
transform 1 0 57316 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1636993656
transform 1 0 58420 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1636993656
transform 1 0 59524 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 25201
transform 1 0 60628 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 25201
transform 1 0 61180 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1636993656
transform 1 0 61364 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1636993656
transform 1 0 62468 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1636993656
transform 1 0 63572 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_681
timestamp 1636993656
transform 1 0 64676 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 25201
transform 1 0 65780 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 25201
transform 1 0 66332 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1636993656
transform 1 0 66516 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1636993656
transform 1 0 67620 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_725
timestamp 1636993656
transform 1 0 68724 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_737
timestamp 1636993656
transform 1 0 69828 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_749
timestamp 25201
transform 1 0 70932 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_755
timestamp 25201
transform 1 0 71484 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_757
timestamp 1636993656
transform 1 0 71668 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_769
timestamp 1636993656
transform 1 0 72772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_781
timestamp 1636993656
transform 1 0 73876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_793
timestamp 1636993656
transform 1 0 74980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_805
timestamp 25201
transform 1 0 76084 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_811
timestamp 25201
transform 1 0 76636 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_813
timestamp 25201
transform 1 0 76820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_821
timestamp 25201
transform 1 0 77556 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636993656
transform 1 0 2300 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636993656
transform 1 0 3404 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636993656
transform 1 0 4508 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636993656
transform 1 0 5612 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 25201
transform 1 0 6716 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 25201
transform 1 0 7084 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636993656
transform 1 0 7268 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1636993656
transform 1 0 8372 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1636993656
transform 1 0 9476 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1636993656
transform 1 0 10580 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 25201
transform 1 0 11684 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 25201
transform 1 0 12236 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1636993656
transform 1 0 12420 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1636993656
transform 1 0 13524 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1636993656
transform 1 0 14628 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1636993656
transform 1 0 15732 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 25201
transform 1 0 16836 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 25201
transform 1 0 17388 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1636993656
transform 1 0 17572 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1636993656
transform 1 0 18676 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1636993656
transform 1 0 19780 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1636993656
transform 1 0 20884 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 25201
transform 1 0 21988 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 25201
transform 1 0 22540 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1636993656
transform 1 0 22724 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1636993656
transform 1 0 23828 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1636993656
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1636993656
transform 1 0 26036 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 25201
transform 1 0 27140 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 25201
transform 1 0 27692 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1636993656
transform 1 0 27876 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1636993656
transform 1 0 28980 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1636993656
transform 1 0 30084 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1636993656
transform 1 0 31188 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 25201
transform 1 0 32292 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 25201
transform 1 0 32844 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1636993656
transform 1 0 33028 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1636993656
transform 1 0 34132 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1636993656
transform 1 0 35236 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1636993656
transform 1 0 36340 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 25201
transform 1 0 37444 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 25201
transform 1 0 37996 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1636993656
transform 1 0 38180 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1636993656
transform 1 0 39284 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1636993656
transform 1 0 40388 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1636993656
transform 1 0 41492 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 25201
transform 1 0 42596 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 25201
transform 1 0 43148 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1636993656
transform 1 0 43332 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1636993656
transform 1 0 44436 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1636993656
transform 1 0 45540 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1636993656
transform 1 0 46644 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 25201
transform 1 0 47748 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 25201
transform 1 0 48300 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1636993656
transform 1 0 48484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1636993656
transform 1 0 49588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1636993656
transform 1 0 50692 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1636993656
transform 1 0 51796 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 25201
transform 1 0 52900 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 25201
transform 1 0 53452 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1636993656
transform 1 0 53636 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1636993656
transform 1 0 54740 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1636993656
transform 1 0 55844 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1636993656
transform 1 0 56948 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 25201
transform 1 0 58052 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 25201
transform 1 0 58604 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1636993656
transform 1 0 58788 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1636993656
transform 1 0 59892 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1636993656
transform 1 0 60996 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1636993656
transform 1 0 62100 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 25201
transform 1 0 63204 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 25201
transform 1 0 63756 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1636993656
transform 1 0 63940 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1636993656
transform 1 0 65044 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1636993656
transform 1 0 66148 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1636993656
transform 1 0 67252 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 25201
transform 1 0 68356 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 25201
transform 1 0 68908 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_729
timestamp 1636993656
transform 1 0 69092 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_741
timestamp 1636993656
transform 1 0 70196 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_753
timestamp 1636993656
transform 1 0 71300 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_765
timestamp 1636993656
transform 1 0 72404 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_777
timestamp 25201
transform 1 0 73508 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_783
timestamp 25201
transform 1 0 74060 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_785
timestamp 1636993656
transform 1 0 74244 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_797
timestamp 1636993656
transform 1 0 75348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_809
timestamp 1636993656
transform 1 0 76452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_821
timestamp 25201
transform 1 0 77556 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636993656
transform 1 0 2300 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636993656
transform 1 0 3404 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 25201
transform 1 0 4508 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636993656
transform 1 0 4692 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636993656
transform 1 0 5796 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636993656
transform 1 0 6900 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1636993656
transform 1 0 8004 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 25201
transform 1 0 9108 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 25201
transform 1 0 9660 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1636993656
transform 1 0 9844 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1636993656
transform 1 0 10948 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1636993656
transform 1 0 12052 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1636993656
transform 1 0 13156 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 25201
transform 1 0 14260 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 25201
transform 1 0 14812 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1636993656
transform 1 0 14996 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1636993656
transform 1 0 16100 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1636993656
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1636993656
transform 1 0 18308 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 25201
transform 1 0 19412 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 25201
transform 1 0 19964 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1636993656
transform 1 0 20148 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1636993656
transform 1 0 21252 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1636993656
transform 1 0 22356 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1636993656
transform 1 0 23460 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 25201
transform 1 0 24564 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 25201
transform 1 0 25116 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1636993656
transform 1 0 25300 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1636993656
transform 1 0 26404 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1636993656
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1636993656
transform 1 0 28612 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 25201
transform 1 0 29716 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 25201
transform 1 0 30268 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1636993656
transform 1 0 30452 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1636993656
transform 1 0 31556 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1636993656
transform 1 0 32660 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1636993656
transform 1 0 33764 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 25201
transform 1 0 34868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 25201
transform 1 0 35420 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1636993656
transform 1 0 35604 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1636993656
transform 1 0 36708 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1636993656
transform 1 0 37812 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1636993656
transform 1 0 38916 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 25201
transform 1 0 40020 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 25201
transform 1 0 40572 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1636993656
transform 1 0 40756 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1636993656
transform 1 0 41860 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1636993656
transform 1 0 42964 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1636993656
transform 1 0 44068 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 25201
transform 1 0 45172 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 25201
transform 1 0 45724 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1636993656
transform 1 0 45908 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1636993656
transform 1 0 47012 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1636993656
transform 1 0 48116 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1636993656
transform 1 0 49220 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 25201
transform 1 0 50324 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 25201
transform 1 0 50876 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1636993656
transform 1 0 51060 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1636993656
transform 1 0 52164 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1636993656
transform 1 0 53268 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1636993656
transform 1 0 54372 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 25201
transform 1 0 55476 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 25201
transform 1 0 56028 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1636993656
transform 1 0 56212 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1636993656
transform 1 0 57316 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1636993656
transform 1 0 58420 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1636993656
transform 1 0 59524 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 25201
transform 1 0 60628 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 25201
transform 1 0 61180 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1636993656
transform 1 0 61364 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1636993656
transform 1 0 62468 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1636993656
transform 1 0 63572 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1636993656
transform 1 0 64676 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 25201
transform 1 0 65780 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 25201
transform 1 0 66332 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1636993656
transform 1 0 66516 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1636993656
transform 1 0 67620 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_725
timestamp 1636993656
transform 1 0 68724 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_737
timestamp 1636993656
transform 1 0 69828 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_749
timestamp 25201
transform 1 0 70932 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_755
timestamp 25201
transform 1 0 71484 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_757
timestamp 1636993656
transform 1 0 71668 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_769
timestamp 1636993656
transform 1 0 72772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_781
timestamp 1636993656
transform 1 0 73876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_793
timestamp 1636993656
transform 1 0 74980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_805
timestamp 25201
transform 1 0 76084 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_811
timestamp 25201
transform 1 0 76636 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_813
timestamp 25201
transform 1 0 76820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_821
timestamp 25201
transform 1 0 77556 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636993656
transform 1 0 2300 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636993656
transform 1 0 3404 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636993656
transform 1 0 4508 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636993656
transform 1 0 5612 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 25201
transform 1 0 6716 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 25201
transform 1 0 7084 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636993656
transform 1 0 7268 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1636993656
transform 1 0 8372 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1636993656
transform 1 0 9476 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1636993656
transform 1 0 10580 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 25201
transform 1 0 11684 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 25201
transform 1 0 12236 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1636993656
transform 1 0 12420 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1636993656
transform 1 0 13524 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1636993656
transform 1 0 14628 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1636993656
transform 1 0 15732 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 25201
transform 1 0 16836 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 25201
transform 1 0 17388 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636993656
transform 1 0 17572 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1636993656
transform 1 0 18676 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1636993656
transform 1 0 19780 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1636993656
transform 1 0 20884 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 25201
transform 1 0 21988 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 25201
transform 1 0 22540 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1636993656
transform 1 0 22724 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1636993656
transform 1 0 23828 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1636993656
transform 1 0 24932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1636993656
transform 1 0 26036 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 25201
transform 1 0 27140 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 25201
transform 1 0 27692 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1636993656
transform 1 0 27876 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1636993656
transform 1 0 28980 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1636993656
transform 1 0 30084 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1636993656
transform 1 0 31188 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 25201
transform 1 0 32292 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 25201
transform 1 0 32844 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1636993656
transform 1 0 33028 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1636993656
transform 1 0 34132 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1636993656
transform 1 0 35236 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1636993656
transform 1 0 36340 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 25201
transform 1 0 37444 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 25201
transform 1 0 37996 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1636993656
transform 1 0 38180 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1636993656
transform 1 0 39284 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1636993656
transform 1 0 40388 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1636993656
transform 1 0 41492 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 25201
transform 1 0 42596 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 25201
transform 1 0 43148 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1636993656
transform 1 0 43332 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1636993656
transform 1 0 44436 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1636993656
transform 1 0 45540 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1636993656
transform 1 0 46644 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 25201
transform 1 0 47748 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 25201
transform 1 0 48300 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1636993656
transform 1 0 48484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1636993656
transform 1 0 49588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1636993656
transform 1 0 50692 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1636993656
transform 1 0 51796 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 25201
transform 1 0 52900 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 25201
transform 1 0 53452 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1636993656
transform 1 0 53636 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1636993656
transform 1 0 54740 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1636993656
transform 1 0 55844 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1636993656
transform 1 0 56948 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 25201
transform 1 0 58052 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 25201
transform 1 0 58604 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_617
timestamp 1636993656
transform 1 0 58788 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_629
timestamp 1636993656
transform 1 0 59892 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_641
timestamp 1636993656
transform 1 0 60996 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_653
timestamp 1636993656
transform 1 0 62100 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 25201
transform 1 0 63204 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 25201
transform 1 0 63756 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1636993656
transform 1 0 63940 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_685
timestamp 1636993656
transform 1 0 65044 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_697
timestamp 1636993656
transform 1 0 66148 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_709
timestamp 1636993656
transform 1 0 67252 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 25201
transform 1 0 68356 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 25201
transform 1 0 68908 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_729
timestamp 1636993656
transform 1 0 69092 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_741
timestamp 1636993656
transform 1 0 70196 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_753
timestamp 1636993656
transform 1 0 71300 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_765
timestamp 1636993656
transform 1 0 72404 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_777
timestamp 25201
transform 1 0 73508 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_783
timestamp 25201
transform 1 0 74060 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_785
timestamp 1636993656
transform 1 0 74244 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_797
timestamp 1636993656
transform 1 0 75348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_809
timestamp 1636993656
transform 1 0 76452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_821
timestamp 25201
transform 1 0 77556 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636993656
transform 1 0 2300 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636993656
transform 1 0 3404 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 25201
transform 1 0 4508 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636993656
transform 1 0 4692 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636993656
transform 1 0 5796 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1636993656
transform 1 0 6900 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1636993656
transform 1 0 8004 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 25201
transform 1 0 9108 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 25201
transform 1 0 9660 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1636993656
transform 1 0 9844 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1636993656
transform 1 0 10948 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1636993656
transform 1 0 12052 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1636993656
transform 1 0 13156 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 25201
transform 1 0 14260 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 25201
transform 1 0 14812 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1636993656
transform 1 0 14996 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1636993656
transform 1 0 16100 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1636993656
transform 1 0 17204 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1636993656
transform 1 0 18308 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 25201
transform 1 0 19412 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 25201
transform 1 0 19964 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1636993656
transform 1 0 20148 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1636993656
transform 1 0 21252 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1636993656
transform 1 0 22356 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1636993656
transform 1 0 23460 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 25201
transform 1 0 24564 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 25201
transform 1 0 25116 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1636993656
transform 1 0 25300 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1636993656
transform 1 0 26404 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1636993656
transform 1 0 27508 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1636993656
transform 1 0 28612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 25201
transform 1 0 29716 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 25201
transform 1 0 30268 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1636993656
transform 1 0 30452 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1636993656
transform 1 0 31556 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1636993656
transform 1 0 32660 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1636993656
transform 1 0 33764 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 25201
transform 1 0 34868 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 25201
transform 1 0 35420 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1636993656
transform 1 0 35604 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1636993656
transform 1 0 36708 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1636993656
transform 1 0 37812 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1636993656
transform 1 0 38916 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 25201
transform 1 0 40020 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 25201
transform 1 0 40572 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1636993656
transform 1 0 40756 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1636993656
transform 1 0 41860 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1636993656
transform 1 0 42964 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1636993656
transform 1 0 44068 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 25201
transform 1 0 45172 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 25201
transform 1 0 45724 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1636993656
transform 1 0 45908 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1636993656
transform 1 0 47012 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1636993656
transform 1 0 48116 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1636993656
transform 1 0 49220 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 25201
transform 1 0 50324 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 25201
transform 1 0 50876 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1636993656
transform 1 0 51060 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1636993656
transform 1 0 52164 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1636993656
transform 1 0 53268 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1636993656
transform 1 0 54372 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 25201
transform 1 0 55476 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 25201
transform 1 0 56028 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1636993656
transform 1 0 56212 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1636993656
transform 1 0 57316 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1636993656
transform 1 0 58420 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_625
timestamp 1636993656
transform 1 0 59524 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 25201
transform 1 0 60628 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 25201
transform 1 0 61180 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_645
timestamp 1636993656
transform 1 0 61364 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_657
timestamp 1636993656
transform 1 0 62468 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_669
timestamp 1636993656
transform 1 0 63572 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_681
timestamp 1636993656
transform 1 0 64676 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 25201
transform 1 0 65780 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 25201
transform 1 0 66332 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_701
timestamp 1636993656
transform 1 0 66516 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_713
timestamp 1636993656
transform 1 0 67620 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_725
timestamp 1636993656
transform 1 0 68724 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_737
timestamp 1636993656
transform 1 0 69828 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_749
timestamp 25201
transform 1 0 70932 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_755
timestamp 25201
transform 1 0 71484 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_757
timestamp 1636993656
transform 1 0 71668 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_769
timestamp 1636993656
transform 1 0 72772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_781
timestamp 1636993656
transform 1 0 73876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_793
timestamp 1636993656
transform 1 0 74980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_805
timestamp 25201
transform 1 0 76084 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_811
timestamp 25201
transform 1 0 76636 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_813
timestamp 25201
transform 1 0 76820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_821
timestamp 25201
transform 1 0 77556 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636993656
transform 1 0 2300 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636993656
transform 1 0 3404 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1636993656
transform 1 0 4508 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1636993656
transform 1 0 5612 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 25201
transform 1 0 6716 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 25201
transform 1 0 7084 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636993656
transform 1 0 7268 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1636993656
transform 1 0 8372 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1636993656
transform 1 0 9476 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1636993656
transform 1 0 10580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 25201
transform 1 0 11684 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 25201
transform 1 0 12236 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1636993656
transform 1 0 12420 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1636993656
transform 1 0 13524 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1636993656
transform 1 0 14628 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1636993656
transform 1 0 15732 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 25201
transform 1 0 16836 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 25201
transform 1 0 17388 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1636993656
transform 1 0 17572 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1636993656
transform 1 0 18676 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1636993656
transform 1 0 19780 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1636993656
transform 1 0 20884 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 25201
transform 1 0 21988 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 25201
transform 1 0 22540 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1636993656
transform 1 0 22724 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1636993656
transform 1 0 23828 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1636993656
transform 1 0 24932 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1636993656
transform 1 0 26036 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 25201
transform 1 0 27140 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 25201
transform 1 0 27692 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1636993656
transform 1 0 27876 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1636993656
transform 1 0 28980 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1636993656
transform 1 0 30084 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1636993656
transform 1 0 31188 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 25201
transform 1 0 32292 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 25201
transform 1 0 32844 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1636993656
transform 1 0 33028 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1636993656
transform 1 0 34132 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1636993656
transform 1 0 35236 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1636993656
transform 1 0 36340 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 25201
transform 1 0 37444 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 25201
transform 1 0 37996 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1636993656
transform 1 0 38180 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1636993656
transform 1 0 39284 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1636993656
transform 1 0 40388 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1636993656
transform 1 0 41492 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 25201
transform 1 0 42596 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 25201
transform 1 0 43148 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1636993656
transform 1 0 43332 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1636993656
transform 1 0 44436 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1636993656
transform 1 0 45540 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1636993656
transform 1 0 46644 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 25201
transform 1 0 47748 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 25201
transform 1 0 48300 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1636993656
transform 1 0 48484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1636993656
transform 1 0 49588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1636993656
transform 1 0 50692 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1636993656
transform 1 0 51796 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 25201
transform 1 0 52900 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 25201
transform 1 0 53452 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1636993656
transform 1 0 53636 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1636993656
transform 1 0 54740 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1636993656
transform 1 0 55844 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1636993656
transform 1 0 56948 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 25201
transform 1 0 58052 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 25201
transform 1 0 58604 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_617
timestamp 1636993656
transform 1 0 58788 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_629
timestamp 1636993656
transform 1 0 59892 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_641
timestamp 1636993656
transform 1 0 60996 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_653
timestamp 1636993656
transform 1 0 62100 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 25201
transform 1 0 63204 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 25201
transform 1 0 63756 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_673
timestamp 1636993656
transform 1 0 63940 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_685
timestamp 1636993656
transform 1 0 65044 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_697
timestamp 1636993656
transform 1 0 66148 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_709
timestamp 1636993656
transform 1 0 67252 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 25201
transform 1 0 68356 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 25201
transform 1 0 68908 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_729
timestamp 1636993656
transform 1 0 69092 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_741
timestamp 1636993656
transform 1 0 70196 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_753
timestamp 1636993656
transform 1 0 71300 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_765
timestamp 1636993656
transform 1 0 72404 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_777
timestamp 25201
transform 1 0 73508 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_783
timestamp 25201
transform 1 0 74060 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_785
timestamp 1636993656
transform 1 0 74244 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_797
timestamp 1636993656
transform 1 0 75348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_809
timestamp 1636993656
transform 1 0 76452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_821
timestamp 25201
transform 1 0 77556 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636993656
transform 1 0 2300 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636993656
transform 1 0 3404 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 25201
transform 1 0 4508 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636993656
transform 1 0 4692 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636993656
transform 1 0 5796 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1636993656
transform 1 0 6900 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1636993656
transform 1 0 8004 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 25201
transform 1 0 9108 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 25201
transform 1 0 9660 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1636993656
transform 1 0 9844 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1636993656
transform 1 0 10948 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1636993656
transform 1 0 12052 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1636993656
transform 1 0 13156 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 25201
transform 1 0 14260 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 25201
transform 1 0 14812 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1636993656
transform 1 0 14996 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1636993656
transform 1 0 16100 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1636993656
transform 1 0 17204 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1636993656
transform 1 0 18308 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 25201
transform 1 0 19412 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 25201
transform 1 0 19964 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1636993656
transform 1 0 20148 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1636993656
transform 1 0 21252 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1636993656
transform 1 0 22356 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1636993656
transform 1 0 23460 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 25201
transform 1 0 24564 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 25201
transform 1 0 25116 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1636993656
transform 1 0 25300 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1636993656
transform 1 0 26404 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1636993656
transform 1 0 27508 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1636993656
transform 1 0 28612 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 25201
transform 1 0 29716 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 25201
transform 1 0 30268 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1636993656
transform 1 0 30452 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1636993656
transform 1 0 31556 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1636993656
transform 1 0 32660 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1636993656
transform 1 0 33764 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 25201
transform 1 0 34868 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 25201
transform 1 0 35420 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1636993656
transform 1 0 35604 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1636993656
transform 1 0 36708 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1636993656
transform 1 0 37812 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1636993656
transform 1 0 38916 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 25201
transform 1 0 40020 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 25201
transform 1 0 40572 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1636993656
transform 1 0 40756 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1636993656
transform 1 0 41860 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1636993656
transform 1 0 42964 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1636993656
transform 1 0 44068 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 25201
transform 1 0 45172 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 25201
transform 1 0 45724 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1636993656
transform 1 0 45908 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1636993656
transform 1 0 47012 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1636993656
transform 1 0 48116 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1636993656
transform 1 0 49220 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 25201
transform 1 0 50324 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 25201
transform 1 0 50876 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1636993656
transform 1 0 51060 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1636993656
transform 1 0 52164 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1636993656
transform 1 0 53268 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1636993656
transform 1 0 54372 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 25201
transform 1 0 55476 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 25201
transform 1 0 56028 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1636993656
transform 1 0 56212 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1636993656
transform 1 0 57316 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1636993656
transform 1 0 58420 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_625
timestamp 1636993656
transform 1 0 59524 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 25201
transform 1 0 60628 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 25201
transform 1 0 61180 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_645
timestamp 1636993656
transform 1 0 61364 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_657
timestamp 1636993656
transform 1 0 62468 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_669
timestamp 1636993656
transform 1 0 63572 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_681
timestamp 1636993656
transform 1 0 64676 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 25201
transform 1 0 65780 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 25201
transform 1 0 66332 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_701
timestamp 1636993656
transform 1 0 66516 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_713
timestamp 1636993656
transform 1 0 67620 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_725
timestamp 1636993656
transform 1 0 68724 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_737
timestamp 1636993656
transform 1 0 69828 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_749
timestamp 25201
transform 1 0 70932 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_755
timestamp 25201
transform 1 0 71484 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_757
timestamp 1636993656
transform 1 0 71668 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_769
timestamp 1636993656
transform 1 0 72772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_781
timestamp 1636993656
transform 1 0 73876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_793
timestamp 1636993656
transform 1 0 74980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_805
timestamp 25201
transform 1 0 76084 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_811
timestamp 25201
transform 1 0 76636 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_813
timestamp 25201
transform 1 0 76820 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_821
timestamp 25201
transform 1 0 77556 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636993656
transform 1 0 2300 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1636993656
transform 1 0 3404 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1636993656
transform 1 0 4508 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1636993656
transform 1 0 5612 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 25201
transform 1 0 6716 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 25201
transform 1 0 7084 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1636993656
transform 1 0 7268 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1636993656
transform 1 0 8372 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1636993656
transform 1 0 9476 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1636993656
transform 1 0 10580 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 25201
transform 1 0 11684 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 25201
transform 1 0 12236 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1636993656
transform 1 0 12420 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1636993656
transform 1 0 13524 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1636993656
transform 1 0 14628 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1636993656
transform 1 0 15732 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 25201
transform 1 0 16836 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 25201
transform 1 0 17388 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1636993656
transform 1 0 17572 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1636993656
transform 1 0 18676 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1636993656
transform 1 0 19780 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1636993656
transform 1 0 20884 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 25201
transform 1 0 21988 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 25201
transform 1 0 22540 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1636993656
transform 1 0 22724 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1636993656
transform 1 0 23828 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1636993656
transform 1 0 24932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1636993656
transform 1 0 26036 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 25201
transform 1 0 27140 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 25201
transform 1 0 27692 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1636993656
transform 1 0 27876 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1636993656
transform 1 0 28980 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1636993656
transform 1 0 30084 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1636993656
transform 1 0 31188 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 25201
transform 1 0 32292 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 25201
transform 1 0 32844 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1636993656
transform 1 0 33028 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1636993656
transform 1 0 34132 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1636993656
transform 1 0 35236 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1636993656
transform 1 0 36340 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 25201
transform 1 0 37444 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 25201
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1636993656
transform 1 0 38180 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1636993656
transform 1 0 39284 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1636993656
transform 1 0 40388 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1636993656
transform 1 0 41492 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 25201
transform 1 0 42596 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 25201
transform 1 0 43148 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1636993656
transform 1 0 43332 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1636993656
transform 1 0 44436 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1636993656
transform 1 0 45540 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1636993656
transform 1 0 46644 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 25201
transform 1 0 47748 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 25201
transform 1 0 48300 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1636993656
transform 1 0 48484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1636993656
transform 1 0 49588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1636993656
transform 1 0 50692 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1636993656
transform 1 0 51796 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 25201
transform 1 0 52900 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 25201
transform 1 0 53452 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1636993656
transform 1 0 53636 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1636993656
transform 1 0 54740 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1636993656
transform 1 0 55844 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1636993656
transform 1 0 56948 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 25201
transform 1 0 58052 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 25201
transform 1 0 58604 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_617
timestamp 1636993656
transform 1 0 58788 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_629
timestamp 1636993656
transform 1 0 59892 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_641
timestamp 1636993656
transform 1 0 60996 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_653
timestamp 1636993656
transform 1 0 62100 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 25201
transform 1 0 63204 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 25201
transform 1 0 63756 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_673
timestamp 1636993656
transform 1 0 63940 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_685
timestamp 1636993656
transform 1 0 65044 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_697
timestamp 1636993656
transform 1 0 66148 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_709
timestamp 1636993656
transform 1 0 67252 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 25201
transform 1 0 68356 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 25201
transform 1 0 68908 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_729
timestamp 1636993656
transform 1 0 69092 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_741
timestamp 1636993656
transform 1 0 70196 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_753
timestamp 1636993656
transform 1 0 71300 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_765
timestamp 1636993656
transform 1 0 72404 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_777
timestamp 25201
transform 1 0 73508 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_783
timestamp 25201
transform 1 0 74060 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_785
timestamp 1636993656
transform 1 0 74244 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_797
timestamp 1636993656
transform 1 0 75348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_809
timestamp 1636993656
transform 1 0 76452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_821
timestamp 25201
transform 1 0 77556 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1636993656
transform 1 0 2300 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1636993656
transform 1 0 3404 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 25201
transform 1 0 4508 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636993656
transform 1 0 4692 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1636993656
transform 1 0 5796 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1636993656
transform 1 0 6900 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1636993656
transform 1 0 8004 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 25201
transform 1 0 9108 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 25201
transform 1 0 9660 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1636993656
transform 1 0 9844 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1636993656
transform 1 0 10948 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1636993656
transform 1 0 12052 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1636993656
transform 1 0 13156 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 25201
transform 1 0 14260 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 25201
transform 1 0 14812 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1636993656
transform 1 0 14996 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1636993656
transform 1 0 16100 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1636993656
transform 1 0 17204 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1636993656
transform 1 0 18308 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 25201
transform 1 0 19412 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 25201
transform 1 0 19964 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1636993656
transform 1 0 20148 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1636993656
transform 1 0 21252 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1636993656
transform 1 0 22356 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1636993656
transform 1 0 23460 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 25201
transform 1 0 24564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 25201
transform 1 0 25116 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1636993656
transform 1 0 25300 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1636993656
transform 1 0 26404 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1636993656
transform 1 0 27508 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1636993656
transform 1 0 28612 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 25201
transform 1 0 29716 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 25201
transform 1 0 30268 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1636993656
transform 1 0 30452 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1636993656
transform 1 0 31556 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1636993656
transform 1 0 32660 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1636993656
transform 1 0 33764 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 25201
transform 1 0 34868 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 25201
transform 1 0 35420 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1636993656
transform 1 0 35604 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1636993656
transform 1 0 36708 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1636993656
transform 1 0 37812 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1636993656
transform 1 0 38916 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 25201
transform 1 0 40020 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 25201
transform 1 0 40572 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1636993656
transform 1 0 40756 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1636993656
transform 1 0 41860 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1636993656
transform 1 0 42964 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1636993656
transform 1 0 44068 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 25201
transform 1 0 45172 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 25201
transform 1 0 45724 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1636993656
transform 1 0 45908 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1636993656
transform 1 0 47012 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1636993656
transform 1 0 48116 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1636993656
transform 1 0 49220 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 25201
transform 1 0 50324 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 25201
transform 1 0 50876 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1636993656
transform 1 0 51060 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1636993656
transform 1 0 52164 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1636993656
transform 1 0 53268 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1636993656
transform 1 0 54372 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 25201
transform 1 0 55476 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 25201
transform 1 0 56028 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1636993656
transform 1 0 56212 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1636993656
transform 1 0 57316 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1636993656
transform 1 0 58420 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_625
timestamp 1636993656
transform 1 0 59524 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 25201
transform 1 0 60628 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 25201
transform 1 0 61180 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_645
timestamp 1636993656
transform 1 0 61364 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_657
timestamp 1636993656
transform 1 0 62468 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_669
timestamp 1636993656
transform 1 0 63572 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_681
timestamp 1636993656
transform 1 0 64676 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 25201
transform 1 0 65780 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 25201
transform 1 0 66332 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_701
timestamp 1636993656
transform 1 0 66516 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_713
timestamp 1636993656
transform 1 0 67620 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_725
timestamp 1636993656
transform 1 0 68724 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_737
timestamp 1636993656
transform 1 0 69828 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_749
timestamp 25201
transform 1 0 70932 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_755
timestamp 25201
transform 1 0 71484 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_757
timestamp 1636993656
transform 1 0 71668 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_769
timestamp 1636993656
transform 1 0 72772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_781
timestamp 1636993656
transform 1 0 73876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_793
timestamp 1636993656
transform 1 0 74980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_805
timestamp 25201
transform 1 0 76084 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_811
timestamp 25201
transform 1 0 76636 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_813
timestamp 25201
transform 1 0 76820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_821
timestamp 25201
transform 1 0 77556 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636993656
transform 1 0 2300 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636993656
transform 1 0 3404 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1636993656
transform 1 0 4508 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1636993656
transform 1 0 5612 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 25201
transform 1 0 6716 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 25201
transform 1 0 7084 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1636993656
transform 1 0 7268 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1636993656
transform 1 0 8372 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1636993656
transform 1 0 9476 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1636993656
transform 1 0 10580 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 25201
transform 1 0 11684 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 25201
transform 1 0 12236 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1636993656
transform 1 0 12420 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1636993656
transform 1 0 13524 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1636993656
transform 1 0 14628 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1636993656
transform 1 0 15732 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 25201
transform 1 0 16836 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 25201
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1636993656
transform 1 0 17572 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1636993656
transform 1 0 18676 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1636993656
transform 1 0 19780 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1636993656
transform 1 0 20884 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 25201
transform 1 0 21988 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 25201
transform 1 0 22540 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1636993656
transform 1 0 22724 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1636993656
transform 1 0 23828 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1636993656
transform 1 0 24932 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1636993656
transform 1 0 26036 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 25201
transform 1 0 27140 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 25201
transform 1 0 27692 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1636993656
transform 1 0 27876 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1636993656
transform 1 0 28980 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1636993656
transform 1 0 30084 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1636993656
transform 1 0 31188 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 25201
transform 1 0 32292 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 25201
transform 1 0 32844 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1636993656
transform 1 0 33028 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1636993656
transform 1 0 34132 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1636993656
transform 1 0 35236 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1636993656
transform 1 0 36340 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 25201
transform 1 0 37444 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 25201
transform 1 0 37996 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1636993656
transform 1 0 38180 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1636993656
transform 1 0 39284 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1636993656
transform 1 0 40388 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1636993656
transform 1 0 41492 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 25201
transform 1 0 42596 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 25201
transform 1 0 43148 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1636993656
transform 1 0 43332 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1636993656
transform 1 0 44436 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1636993656
transform 1 0 45540 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1636993656
transform 1 0 46644 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 25201
transform 1 0 47748 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 25201
transform 1 0 48300 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1636993656
transform 1 0 48484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1636993656
transform 1 0 49588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1636993656
transform 1 0 50692 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1636993656
transform 1 0 51796 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 25201
transform 1 0 52900 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 25201
transform 1 0 53452 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1636993656
transform 1 0 53636 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1636993656
transform 1 0 54740 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1636993656
transform 1 0 55844 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1636993656
transform 1 0 56948 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 25201
transform 1 0 58052 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 25201
transform 1 0 58604 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_617
timestamp 1636993656
transform 1 0 58788 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_629
timestamp 1636993656
transform 1 0 59892 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_641
timestamp 1636993656
transform 1 0 60996 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_653
timestamp 1636993656
transform 1 0 62100 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 25201
transform 1 0 63204 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 25201
transform 1 0 63756 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_673
timestamp 1636993656
transform 1 0 63940 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_685
timestamp 1636993656
transform 1 0 65044 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_697
timestamp 1636993656
transform 1 0 66148 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_709
timestamp 1636993656
transform 1 0 67252 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 25201
transform 1 0 68356 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 25201
transform 1 0 68908 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_729
timestamp 1636993656
transform 1 0 69092 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_741
timestamp 1636993656
transform 1 0 70196 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_753
timestamp 1636993656
transform 1 0 71300 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_765
timestamp 1636993656
transform 1 0 72404 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_777
timestamp 25201
transform 1 0 73508 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_783
timestamp 25201
transform 1 0 74060 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_785
timestamp 1636993656
transform 1 0 74244 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_797
timestamp 1636993656
transform 1 0 75348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_809
timestamp 1636993656
transform 1 0 76452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_821
timestamp 25201
transform 1 0 77556 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636993656
transform 1 0 2300 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636993656
transform 1 0 3404 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 25201
transform 1 0 4508 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636993656
transform 1 0 4692 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1636993656
transform 1 0 5796 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1636993656
transform 1 0 6900 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1636993656
transform 1 0 8004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 25201
transform 1 0 9108 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 25201
transform 1 0 9660 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1636993656
transform 1 0 9844 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1636993656
transform 1 0 10948 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1636993656
transform 1 0 12052 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1636993656
transform 1 0 13156 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 25201
transform 1 0 14260 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 25201
transform 1 0 14812 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1636993656
transform 1 0 14996 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1636993656
transform 1 0 16100 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1636993656
transform 1 0 17204 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1636993656
transform 1 0 18308 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 25201
transform 1 0 19412 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 25201
transform 1 0 19964 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1636993656
transform 1 0 20148 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1636993656
transform 1 0 21252 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1636993656
transform 1 0 22356 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1636993656
transform 1 0 23460 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 25201
transform 1 0 24564 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 25201
transform 1 0 25116 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1636993656
transform 1 0 25300 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1636993656
transform 1 0 26404 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1636993656
transform 1 0 27508 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1636993656
transform 1 0 28612 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 25201
transform 1 0 29716 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 25201
transform 1 0 30268 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1636993656
transform 1 0 30452 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1636993656
transform 1 0 31556 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1636993656
transform 1 0 32660 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1636993656
transform 1 0 33764 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 25201
transform 1 0 34868 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 25201
transform 1 0 35420 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1636993656
transform 1 0 35604 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1636993656
transform 1 0 36708 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1636993656
transform 1 0 37812 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1636993656
transform 1 0 38916 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 25201
transform 1 0 40020 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 25201
transform 1 0 40572 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1636993656
transform 1 0 40756 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1636993656
transform 1 0 41860 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1636993656
transform 1 0 42964 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1636993656
transform 1 0 44068 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 25201
transform 1 0 45172 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 25201
transform 1 0 45724 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1636993656
transform 1 0 45908 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1636993656
transform 1 0 47012 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1636993656
transform 1 0 48116 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1636993656
transform 1 0 49220 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 25201
transform 1 0 50324 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 25201
transform 1 0 50876 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1636993656
transform 1 0 51060 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1636993656
transform 1 0 52164 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1636993656
transform 1 0 53268 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1636993656
transform 1 0 54372 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 25201
transform 1 0 55476 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 25201
transform 1 0 56028 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1636993656
transform 1 0 56212 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1636993656
transform 1 0 57316 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1636993656
transform 1 0 58420 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_625
timestamp 1636993656
transform 1 0 59524 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 25201
transform 1 0 60628 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 25201
transform 1 0 61180 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_645
timestamp 1636993656
transform 1 0 61364 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_657
timestamp 1636993656
transform 1 0 62468 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_669
timestamp 1636993656
transform 1 0 63572 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_681
timestamp 1636993656
transform 1 0 64676 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 25201
transform 1 0 65780 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 25201
transform 1 0 66332 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_701
timestamp 1636993656
transform 1 0 66516 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_713
timestamp 1636993656
transform 1 0 67620 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_725
timestamp 1636993656
transform 1 0 68724 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_737
timestamp 1636993656
transform 1 0 69828 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_749
timestamp 25201
transform 1 0 70932 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_755
timestamp 25201
transform 1 0 71484 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_757
timestamp 1636993656
transform 1 0 71668 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_769
timestamp 1636993656
transform 1 0 72772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_781
timestamp 1636993656
transform 1 0 73876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_793
timestamp 1636993656
transform 1 0 74980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_805
timestamp 25201
transform 1 0 76084 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_811
timestamp 25201
transform 1 0 76636 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_813
timestamp 25201
transform 1 0 76820 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_821
timestamp 25201
transform 1 0 77556 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636993656
transform 1 0 2300 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636993656
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636993656
transform 1 0 4508 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1636993656
transform 1 0 5612 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 25201
transform 1 0 6716 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 25201
transform 1 0 7084 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1636993656
transform 1 0 7268 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1636993656
transform 1 0 8372 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1636993656
transform 1 0 9476 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1636993656
transform 1 0 10580 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 25201
transform 1 0 11684 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 25201
transform 1 0 12236 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1636993656
transform 1 0 12420 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1636993656
transform 1 0 13524 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1636993656
transform 1 0 14628 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1636993656
transform 1 0 15732 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 25201
transform 1 0 16836 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 25201
transform 1 0 17388 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1636993656
transform 1 0 17572 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1636993656
transform 1 0 18676 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1636993656
transform 1 0 19780 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1636993656
transform 1 0 20884 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 25201
transform 1 0 21988 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 25201
transform 1 0 22540 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1636993656
transform 1 0 22724 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1636993656
transform 1 0 23828 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1636993656
transform 1 0 24932 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1636993656
transform 1 0 26036 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 25201
transform 1 0 27140 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 25201
transform 1 0 27692 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1636993656
transform 1 0 27876 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1636993656
transform 1 0 28980 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1636993656
transform 1 0 30084 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1636993656
transform 1 0 31188 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 25201
transform 1 0 32292 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 25201
transform 1 0 32844 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1636993656
transform 1 0 33028 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1636993656
transform 1 0 34132 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1636993656
transform 1 0 35236 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1636993656
transform 1 0 36340 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 25201
transform 1 0 37444 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 25201
transform 1 0 37996 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1636993656
transform 1 0 38180 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1636993656
transform 1 0 39284 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1636993656
transform 1 0 40388 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1636993656
transform 1 0 41492 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 25201
transform 1 0 42596 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 25201
transform 1 0 43148 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1636993656
transform 1 0 43332 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1636993656
transform 1 0 44436 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1636993656
transform 1 0 45540 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1636993656
transform 1 0 46644 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 25201
transform 1 0 47748 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 25201
transform 1 0 48300 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1636993656
transform 1 0 48484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1636993656
transform 1 0 49588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1636993656
transform 1 0 50692 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1636993656
transform 1 0 51796 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 25201
transform 1 0 52900 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 25201
transform 1 0 53452 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1636993656
transform 1 0 53636 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1636993656
transform 1 0 54740 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1636993656
transform 1 0 55844 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1636993656
transform 1 0 56948 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 25201
transform 1 0 58052 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 25201
transform 1 0 58604 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_617
timestamp 1636993656
transform 1 0 58788 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_629
timestamp 1636993656
transform 1 0 59892 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_641
timestamp 1636993656
transform 1 0 60996 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_653
timestamp 1636993656
transform 1 0 62100 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 25201
transform 1 0 63204 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 25201
transform 1 0 63756 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_673
timestamp 1636993656
transform 1 0 63940 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_685
timestamp 1636993656
transform 1 0 65044 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_697
timestamp 1636993656
transform 1 0 66148 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_709
timestamp 1636993656
transform 1 0 67252 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 25201
transform 1 0 68356 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 25201
transform 1 0 68908 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_729
timestamp 1636993656
transform 1 0 69092 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_741
timestamp 1636993656
transform 1 0 70196 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_753
timestamp 1636993656
transform 1 0 71300 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_765
timestamp 1636993656
transform 1 0 72404 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_777
timestamp 25201
transform 1 0 73508 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_783
timestamp 25201
transform 1 0 74060 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_785
timestamp 1636993656
transform 1 0 74244 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_797
timestamp 1636993656
transform 1 0 75348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_809
timestamp 1636993656
transform 1 0 76452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_821
timestamp 25201
transform 1 0 77556 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636993656
transform 1 0 2300 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636993656
transform 1 0 3404 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 25201
transform 1 0 4508 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1636993656
transform 1 0 4692 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1636993656
transform 1 0 5796 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1636993656
transform 1 0 6900 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1636993656
transform 1 0 8004 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 25201
transform 1 0 9108 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 25201
transform 1 0 9660 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1636993656
transform 1 0 9844 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1636993656
transform 1 0 10948 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1636993656
transform 1 0 12052 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1636993656
transform 1 0 13156 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 25201
transform 1 0 14260 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 25201
transform 1 0 14812 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1636993656
transform 1 0 14996 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1636993656
transform 1 0 16100 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1636993656
transform 1 0 17204 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1636993656
transform 1 0 18308 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 25201
transform 1 0 19412 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 25201
transform 1 0 19964 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1636993656
transform 1 0 20148 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1636993656
transform 1 0 21252 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1636993656
transform 1 0 22356 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1636993656
transform 1 0 23460 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 25201
transform 1 0 24564 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 25201
transform 1 0 25116 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1636993656
transform 1 0 25300 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1636993656
transform 1 0 26404 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1636993656
transform 1 0 27508 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1636993656
transform 1 0 28612 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 25201
transform 1 0 29716 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 25201
transform 1 0 30268 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1636993656
transform 1 0 30452 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1636993656
transform 1 0 31556 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1636993656
transform 1 0 32660 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1636993656
transform 1 0 33764 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 25201
transform 1 0 34868 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 25201
transform 1 0 35420 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1636993656
transform 1 0 35604 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1636993656
transform 1 0 36708 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1636993656
transform 1 0 37812 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1636993656
transform 1 0 38916 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 25201
transform 1 0 40020 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 25201
transform 1 0 40572 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1636993656
transform 1 0 40756 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1636993656
transform 1 0 41860 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1636993656
transform 1 0 42964 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1636993656
transform 1 0 44068 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 25201
transform 1 0 45172 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 25201
transform 1 0 45724 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1636993656
transform 1 0 45908 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1636993656
transform 1 0 47012 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1636993656
transform 1 0 48116 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1636993656
transform 1 0 49220 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 25201
transform 1 0 50324 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 25201
transform 1 0 50876 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1636993656
transform 1 0 51060 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1636993656
transform 1 0 52164 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1636993656
transform 1 0 53268 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1636993656
transform 1 0 54372 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 25201
transform 1 0 55476 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 25201
transform 1 0 56028 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1636993656
transform 1 0 56212 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1636993656
transform 1 0 57316 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1636993656
transform 1 0 58420 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_625
timestamp 1636993656
transform 1 0 59524 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 25201
transform 1 0 60628 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 25201
transform 1 0 61180 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_645
timestamp 1636993656
transform 1 0 61364 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_657
timestamp 1636993656
transform 1 0 62468 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_669
timestamp 1636993656
transform 1 0 63572 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_681
timestamp 1636993656
transform 1 0 64676 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 25201
transform 1 0 65780 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 25201
transform 1 0 66332 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_701
timestamp 1636993656
transform 1 0 66516 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_713
timestamp 1636993656
transform 1 0 67620 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_725
timestamp 1636993656
transform 1 0 68724 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_737
timestamp 1636993656
transform 1 0 69828 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_749
timestamp 25201
transform 1 0 70932 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_755
timestamp 25201
transform 1 0 71484 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_757
timestamp 1636993656
transform 1 0 71668 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_769
timestamp 1636993656
transform 1 0 72772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_781
timestamp 1636993656
transform 1 0 73876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_793
timestamp 1636993656
transform 1 0 74980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_805
timestamp 25201
transform 1 0 76084 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_811
timestamp 25201
transform 1 0 76636 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_813
timestamp 25201
transform 1 0 76820 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_821
timestamp 25201
transform 1 0 77556 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1636993656
transform 1 0 2300 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1636993656
transform 1 0 3404 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1636993656
transform 1 0 4508 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1636993656
transform 1 0 5612 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 25201
transform 1 0 6716 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 25201
transform 1 0 7084 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1636993656
transform 1 0 7268 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1636993656
transform 1 0 8372 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1636993656
transform 1 0 9476 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1636993656
transform 1 0 10580 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 25201
transform 1 0 11684 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 25201
transform 1 0 12236 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1636993656
transform 1 0 12420 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1636993656
transform 1 0 13524 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1636993656
transform 1 0 14628 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1636993656
transform 1 0 15732 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 25201
transform 1 0 16836 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 25201
transform 1 0 17388 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1636993656
transform 1 0 17572 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1636993656
transform 1 0 18676 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1636993656
transform 1 0 19780 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1636993656
transform 1 0 20884 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 25201
transform 1 0 21988 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 25201
transform 1 0 22540 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1636993656
transform 1 0 22724 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1636993656
transform 1 0 23828 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1636993656
transform 1 0 24932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1636993656
transform 1 0 26036 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 25201
transform 1 0 27140 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 25201
transform 1 0 27692 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1636993656
transform 1 0 27876 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1636993656
transform 1 0 28980 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1636993656
transform 1 0 30084 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1636993656
transform 1 0 31188 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 25201
transform 1 0 32292 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 25201
transform 1 0 32844 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1636993656
transform 1 0 33028 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1636993656
transform 1 0 34132 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1636993656
transform 1 0 35236 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1636993656
transform 1 0 36340 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 25201
transform 1 0 37444 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 25201
transform 1 0 37996 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1636993656
transform 1 0 38180 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1636993656
transform 1 0 39284 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1636993656
transform 1 0 40388 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1636993656
transform 1 0 41492 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 25201
transform 1 0 42596 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 25201
transform 1 0 43148 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1636993656
transform 1 0 43332 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1636993656
transform 1 0 44436 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1636993656
transform 1 0 45540 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1636993656
transform 1 0 46644 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 25201
transform 1 0 47748 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 25201
transform 1 0 48300 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1636993656
transform 1 0 48484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1636993656
transform 1 0 49588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1636993656
transform 1 0 50692 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1636993656
transform 1 0 51796 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 25201
transform 1 0 52900 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 25201
transform 1 0 53452 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1636993656
transform 1 0 53636 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1636993656
transform 1 0 54740 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1636993656
transform 1 0 55844 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1636993656
transform 1 0 56948 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 25201
transform 1 0 58052 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 25201
transform 1 0 58604 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_617
timestamp 1636993656
transform 1 0 58788 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_629
timestamp 1636993656
transform 1 0 59892 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_641
timestamp 1636993656
transform 1 0 60996 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_653
timestamp 1636993656
transform 1 0 62100 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 25201
transform 1 0 63204 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 25201
transform 1 0 63756 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_673
timestamp 1636993656
transform 1 0 63940 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_685
timestamp 1636993656
transform 1 0 65044 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_697
timestamp 1636993656
transform 1 0 66148 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_709
timestamp 1636993656
transform 1 0 67252 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_721
timestamp 25201
transform 1 0 68356 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_727
timestamp 25201
transform 1 0 68908 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_729
timestamp 1636993656
transform 1 0 69092 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_741
timestamp 1636993656
transform 1 0 70196 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_753
timestamp 1636993656
transform 1 0 71300 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_765
timestamp 1636993656
transform 1 0 72404 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_777
timestamp 25201
transform 1 0 73508 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_783
timestamp 25201
transform 1 0 74060 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_785
timestamp 1636993656
transform 1 0 74244 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_797
timestamp 1636993656
transform 1 0 75348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_809
timestamp 1636993656
transform 1 0 76452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_821
timestamp 25201
transform 1 0 77556 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636993656
transform 1 0 2300 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636993656
transform 1 0 3404 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 25201
transform 1 0 4508 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636993656
transform 1 0 4692 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1636993656
transform 1 0 5796 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1636993656
transform 1 0 6900 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1636993656
transform 1 0 8004 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 25201
transform 1 0 9108 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 25201
transform 1 0 9660 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1636993656
transform 1 0 9844 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1636993656
transform 1 0 10948 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1636993656
transform 1 0 12052 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1636993656
transform 1 0 13156 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 25201
transform 1 0 14260 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 25201
transform 1 0 14812 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1636993656
transform 1 0 14996 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1636993656
transform 1 0 16100 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1636993656
transform 1 0 17204 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1636993656
transform 1 0 18308 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 25201
transform 1 0 19412 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 25201
transform 1 0 19964 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1636993656
transform 1 0 20148 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1636993656
transform 1 0 21252 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1636993656
transform 1 0 22356 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1636993656
transform 1 0 23460 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 25201
transform 1 0 24564 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 25201
transform 1 0 25116 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1636993656
transform 1 0 25300 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1636993656
transform 1 0 26404 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1636993656
transform 1 0 27508 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1636993656
transform 1 0 28612 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 25201
transform 1 0 29716 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 25201
transform 1 0 30268 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1636993656
transform 1 0 30452 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1636993656
transform 1 0 31556 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1636993656
transform 1 0 32660 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1636993656
transform 1 0 33764 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 25201
transform 1 0 34868 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 25201
transform 1 0 35420 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1636993656
transform 1 0 35604 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1636993656
transform 1 0 36708 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1636993656
transform 1 0 37812 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1636993656
transform 1 0 38916 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 25201
transform 1 0 40020 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 25201
transform 1 0 40572 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1636993656
transform 1 0 40756 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1636993656
transform 1 0 41860 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1636993656
transform 1 0 42964 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1636993656
transform 1 0 44068 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 25201
transform 1 0 45172 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 25201
transform 1 0 45724 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1636993656
transform 1 0 45908 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1636993656
transform 1 0 47012 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1636993656
transform 1 0 48116 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1636993656
transform 1 0 49220 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 25201
transform 1 0 50324 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 25201
transform 1 0 50876 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1636993656
transform 1 0 51060 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1636993656
transform 1 0 52164 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1636993656
transform 1 0 53268 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1636993656
transform 1 0 54372 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 25201
transform 1 0 55476 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 25201
transform 1 0 56028 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1636993656
transform 1 0 56212 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1636993656
transform 1 0 57316 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1636993656
transform 1 0 58420 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_625
timestamp 1636993656
transform 1 0 59524 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 25201
transform 1 0 60628 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 25201
transform 1 0 61180 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_645
timestamp 1636993656
transform 1 0 61364 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_657
timestamp 1636993656
transform 1 0 62468 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_669
timestamp 1636993656
transform 1 0 63572 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_681
timestamp 1636993656
transform 1 0 64676 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 25201
transform 1 0 65780 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 25201
transform 1 0 66332 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_701
timestamp 1636993656
transform 1 0 66516 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_713
timestamp 1636993656
transform 1 0 67620 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_725
timestamp 1636993656
transform 1 0 68724 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_737
timestamp 1636993656
transform 1 0 69828 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_749
timestamp 25201
transform 1 0 70932 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_755
timestamp 25201
transform 1 0 71484 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_757
timestamp 1636993656
transform 1 0 71668 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_769
timestamp 1636993656
transform 1 0 72772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_781
timestamp 1636993656
transform 1 0 73876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_793
timestamp 1636993656
transform 1 0 74980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_805
timestamp 25201
transform 1 0 76084 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_811
timestamp 25201
transform 1 0 76636 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_813
timestamp 25201
transform 1 0 76820 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_821
timestamp 25201
transform 1 0 77556 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1636993656
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1636993656
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1636993656
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1636993656
transform 1 0 5612 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 25201
transform 1 0 6716 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 25201
transform 1 0 7084 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1636993656
transform 1 0 7268 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1636993656
transform 1 0 8372 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1636993656
transform 1 0 9476 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1636993656
transform 1 0 10580 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 25201
transform 1 0 11684 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 25201
transform 1 0 12236 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1636993656
transform 1 0 12420 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1636993656
transform 1 0 13524 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1636993656
transform 1 0 14628 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1636993656
transform 1 0 15732 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 25201
transform 1 0 16836 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 25201
transform 1 0 17388 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1636993656
transform 1 0 17572 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1636993656
transform 1 0 18676 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1636993656
transform 1 0 19780 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1636993656
transform 1 0 20884 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 25201
transform 1 0 21988 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 25201
transform 1 0 22540 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1636993656
transform 1 0 22724 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1636993656
transform 1 0 23828 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1636993656
transform 1 0 24932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1636993656
transform 1 0 26036 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 25201
transform 1 0 27140 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 25201
transform 1 0 27692 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1636993656
transform 1 0 27876 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1636993656
transform 1 0 28980 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1636993656
transform 1 0 30084 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1636993656
transform 1 0 31188 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 25201
transform 1 0 32292 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 25201
transform 1 0 32844 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1636993656
transform 1 0 33028 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1636993656
transform 1 0 34132 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1636993656
transform 1 0 35236 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1636993656
transform 1 0 36340 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 25201
transform 1 0 37444 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 25201
transform 1 0 37996 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1636993656
transform 1 0 38180 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1636993656
transform 1 0 39284 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1636993656
transform 1 0 40388 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1636993656
transform 1 0 41492 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 25201
transform 1 0 42596 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 25201
transform 1 0 43148 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1636993656
transform 1 0 43332 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1636993656
transform 1 0 44436 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1636993656
transform 1 0 45540 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1636993656
transform 1 0 46644 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 25201
transform 1 0 47748 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 25201
transform 1 0 48300 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1636993656
transform 1 0 48484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1636993656
transform 1 0 49588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1636993656
transform 1 0 50692 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1636993656
transform 1 0 51796 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 25201
transform 1 0 52900 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 25201
transform 1 0 53452 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1636993656
transform 1 0 53636 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1636993656
transform 1 0 54740 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1636993656
transform 1 0 55844 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1636993656
transform 1 0 56948 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 25201
transform 1 0 58052 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 25201
transform 1 0 58604 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_617
timestamp 1636993656
transform 1 0 58788 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_629
timestamp 1636993656
transform 1 0 59892 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_641
timestamp 1636993656
transform 1 0 60996 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_653
timestamp 1636993656
transform 1 0 62100 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 25201
transform 1 0 63204 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 25201
transform 1 0 63756 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_673
timestamp 1636993656
transform 1 0 63940 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_685
timestamp 1636993656
transform 1 0 65044 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_697
timestamp 1636993656
transform 1 0 66148 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_709
timestamp 1636993656
transform 1 0 67252 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 25201
transform 1 0 68356 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 25201
transform 1 0 68908 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_729
timestamp 1636993656
transform 1 0 69092 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_741
timestamp 1636993656
transform 1 0 70196 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_753
timestamp 1636993656
transform 1 0 71300 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_765
timestamp 1636993656
transform 1 0 72404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_777
timestamp 25201
transform 1 0 73508 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_783
timestamp 25201
transform 1 0 74060 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_785
timestamp 1636993656
transform 1 0 74244 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_797
timestamp 1636993656
transform 1 0 75348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_809
timestamp 1636993656
transform 1 0 76452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_821
timestamp 25201
transform 1 0 77556 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636993656
transform 1 0 2300 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636993656
transform 1 0 3404 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 25201
transform 1 0 4508 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636993656
transform 1 0 4692 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1636993656
transform 1 0 5796 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1636993656
transform 1 0 6900 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1636993656
transform 1 0 8004 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 25201
transform 1 0 9108 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 25201
transform 1 0 9660 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1636993656
transform 1 0 9844 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1636993656
transform 1 0 10948 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1636993656
transform 1 0 12052 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1636993656
transform 1 0 13156 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 25201
transform 1 0 14260 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 25201
transform 1 0 14812 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1636993656
transform 1 0 14996 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1636993656
transform 1 0 16100 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1636993656
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1636993656
transform 1 0 18308 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 25201
transform 1 0 19412 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 25201
transform 1 0 19964 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1636993656
transform 1 0 20148 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1636993656
transform 1 0 21252 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1636993656
transform 1 0 22356 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1636993656
transform 1 0 23460 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 25201
transform 1 0 24564 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 25201
transform 1 0 25116 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1636993656
transform 1 0 25300 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1636993656
transform 1 0 26404 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1636993656
transform 1 0 27508 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1636993656
transform 1 0 28612 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 25201
transform 1 0 29716 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 25201
transform 1 0 30268 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1636993656
transform 1 0 30452 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1636993656
transform 1 0 31556 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1636993656
transform 1 0 32660 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1636993656
transform 1 0 33764 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 25201
transform 1 0 34868 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 25201
transform 1 0 35420 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1636993656
transform 1 0 35604 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1636993656
transform 1 0 36708 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1636993656
transform 1 0 37812 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1636993656
transform 1 0 38916 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 25201
transform 1 0 40020 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 25201
transform 1 0 40572 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1636993656
transform 1 0 40756 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1636993656
transform 1 0 41860 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1636993656
transform 1 0 42964 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1636993656
transform 1 0 44068 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 25201
transform 1 0 45172 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 25201
transform 1 0 45724 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1636993656
transform 1 0 45908 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1636993656
transform 1 0 47012 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1636993656
transform 1 0 48116 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1636993656
transform 1 0 49220 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 25201
transform 1 0 50324 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 25201
transform 1 0 50876 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1636993656
transform 1 0 51060 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1636993656
transform 1 0 52164 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1636993656
transform 1 0 53268 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1636993656
transform 1 0 54372 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 25201
transform 1 0 55476 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 25201
transform 1 0 56028 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1636993656
transform 1 0 56212 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1636993656
transform 1 0 57316 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1636993656
transform 1 0 58420 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_625
timestamp 1636993656
transform 1 0 59524 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 25201
transform 1 0 60628 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 25201
transform 1 0 61180 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_645
timestamp 1636993656
transform 1 0 61364 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_657
timestamp 1636993656
transform 1 0 62468 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_669
timestamp 1636993656
transform 1 0 63572 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_681
timestamp 1636993656
transform 1 0 64676 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 25201
transform 1 0 65780 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 25201
transform 1 0 66332 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_701
timestamp 1636993656
transform 1 0 66516 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_713
timestamp 1636993656
transform 1 0 67620 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_725
timestamp 1636993656
transform 1 0 68724 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_737
timestamp 1636993656
transform 1 0 69828 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_749
timestamp 25201
transform 1 0 70932 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_755
timestamp 25201
transform 1 0 71484 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_757
timestamp 1636993656
transform 1 0 71668 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_769
timestamp 1636993656
transform 1 0 72772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_781
timestamp 1636993656
transform 1 0 73876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_793
timestamp 1636993656
transform 1 0 74980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_805
timestamp 25201
transform 1 0 76084 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_811
timestamp 25201
transform 1 0 76636 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_813
timestamp 25201
transform 1 0 76820 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_821
timestamp 25201
transform 1 0 77556 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636993656
transform 1 0 2300 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636993656
transform 1 0 3404 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1636993656
transform 1 0 4508 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1636993656
transform 1 0 5612 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 25201
transform 1 0 6716 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 25201
transform 1 0 7084 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1636993656
transform 1 0 7268 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1636993656
transform 1 0 8372 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1636993656
transform 1 0 9476 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1636993656
transform 1 0 10580 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 25201
transform 1 0 11684 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 25201
transform 1 0 12236 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1636993656
transform 1 0 12420 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1636993656
transform 1 0 13524 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1636993656
transform 1 0 14628 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1636993656
transform 1 0 15732 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 25201
transform 1 0 16836 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 25201
transform 1 0 17388 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1636993656
transform 1 0 17572 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1636993656
transform 1 0 18676 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1636993656
transform 1 0 19780 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1636993656
transform 1 0 20884 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 25201
transform 1 0 21988 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 25201
transform 1 0 22540 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1636993656
transform 1 0 22724 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1636993656
transform 1 0 23828 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1636993656
transform 1 0 24932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1636993656
transform 1 0 26036 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 25201
transform 1 0 27140 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 25201
transform 1 0 27692 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1636993656
transform 1 0 27876 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1636993656
transform 1 0 28980 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1636993656
transform 1 0 30084 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1636993656
transform 1 0 31188 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 25201
transform 1 0 32292 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 25201
transform 1 0 32844 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1636993656
transform 1 0 33028 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1636993656
transform 1 0 34132 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1636993656
transform 1 0 35236 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1636993656
transform 1 0 36340 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 25201
transform 1 0 37444 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 25201
transform 1 0 37996 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1636993656
transform 1 0 38180 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1636993656
transform 1 0 39284 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1636993656
transform 1 0 40388 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1636993656
transform 1 0 41492 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 25201
transform 1 0 42596 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 25201
transform 1 0 43148 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1636993656
transform 1 0 43332 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1636993656
transform 1 0 44436 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1636993656
transform 1 0 45540 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1636993656
transform 1 0 46644 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 25201
transform 1 0 47748 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 25201
transform 1 0 48300 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1636993656
transform 1 0 48484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1636993656
transform 1 0 49588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1636993656
transform 1 0 50692 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1636993656
transform 1 0 51796 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 25201
transform 1 0 52900 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 25201
transform 1 0 53452 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1636993656
transform 1 0 53636 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1636993656
transform 1 0 54740 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1636993656
transform 1 0 55844 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1636993656
transform 1 0 56948 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 25201
transform 1 0 58052 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 25201
transform 1 0 58604 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_617
timestamp 1636993656
transform 1 0 58788 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_629
timestamp 1636993656
transform 1 0 59892 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_641
timestamp 1636993656
transform 1 0 60996 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_653
timestamp 1636993656
transform 1 0 62100 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 25201
transform 1 0 63204 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 25201
transform 1 0 63756 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_673
timestamp 1636993656
transform 1 0 63940 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_685
timestamp 1636993656
transform 1 0 65044 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_697
timestamp 1636993656
transform 1 0 66148 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_709
timestamp 1636993656
transform 1 0 67252 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 25201
transform 1 0 68356 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 25201
transform 1 0 68908 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_729
timestamp 1636993656
transform 1 0 69092 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_741
timestamp 1636993656
transform 1 0 70196 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_753
timestamp 1636993656
transform 1 0 71300 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_765
timestamp 1636993656
transform 1 0 72404 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_777
timestamp 25201
transform 1 0 73508 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_783
timestamp 25201
transform 1 0 74060 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_785
timestamp 1636993656
transform 1 0 74244 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_797
timestamp 1636993656
transform 1 0 75348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_809
timestamp 1636993656
transform 1 0 76452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_821
timestamp 25201
transform 1 0 77556 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1636993656
transform 1 0 2300 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1636993656
transform 1 0 3404 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 25201
transform 1 0 4508 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636993656
transform 1 0 4692 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1636993656
transform 1 0 5796 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1636993656
transform 1 0 6900 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1636993656
transform 1 0 8004 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 25201
transform 1 0 9108 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 25201
transform 1 0 9660 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1636993656
transform 1 0 9844 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1636993656
transform 1 0 10948 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1636993656
transform 1 0 12052 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1636993656
transform 1 0 13156 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 25201
transform 1 0 14260 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 25201
transform 1 0 14812 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1636993656
transform 1 0 14996 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1636993656
transform 1 0 16100 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1636993656
transform 1 0 17204 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1636993656
transform 1 0 18308 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 25201
transform 1 0 19412 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 25201
transform 1 0 19964 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1636993656
transform 1 0 20148 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1636993656
transform 1 0 21252 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1636993656
transform 1 0 22356 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1636993656
transform 1 0 23460 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 25201
transform 1 0 24564 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 25201
transform 1 0 25116 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1636993656
transform 1 0 25300 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1636993656
transform 1 0 26404 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1636993656
transform 1 0 27508 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1636993656
transform 1 0 28612 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 25201
transform 1 0 29716 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 25201
transform 1 0 30268 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1636993656
transform 1 0 30452 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1636993656
transform 1 0 31556 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1636993656
transform 1 0 32660 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1636993656
transform 1 0 33764 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 25201
transform 1 0 34868 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 25201
transform 1 0 35420 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1636993656
transform 1 0 35604 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1636993656
transform 1 0 36708 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1636993656
transform 1 0 37812 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1636993656
transform 1 0 38916 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 25201
transform 1 0 40020 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 25201
transform 1 0 40572 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1636993656
transform 1 0 40756 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1636993656
transform 1 0 41860 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1636993656
transform 1 0 42964 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1636993656
transform 1 0 44068 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 25201
transform 1 0 45172 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 25201
transform 1 0 45724 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1636993656
transform 1 0 45908 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1636993656
transform 1 0 47012 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1636993656
transform 1 0 48116 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1636993656
transform 1 0 49220 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 25201
transform 1 0 50324 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 25201
transform 1 0 50876 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1636993656
transform 1 0 51060 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1636993656
transform 1 0 52164 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1636993656
transform 1 0 53268 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1636993656
transform 1 0 54372 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 25201
transform 1 0 55476 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 25201
transform 1 0 56028 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1636993656
transform 1 0 56212 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1636993656
transform 1 0 57316 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1636993656
transform 1 0 58420 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_625
timestamp 1636993656
transform 1 0 59524 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 25201
transform 1 0 60628 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 25201
transform 1 0 61180 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_645
timestamp 1636993656
transform 1 0 61364 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_657
timestamp 1636993656
transform 1 0 62468 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_669
timestamp 1636993656
transform 1 0 63572 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_681
timestamp 1636993656
transform 1 0 64676 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 25201
transform 1 0 65780 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 25201
transform 1 0 66332 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_701
timestamp 1636993656
transform 1 0 66516 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_713
timestamp 1636993656
transform 1 0 67620 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_725
timestamp 1636993656
transform 1 0 68724 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_737
timestamp 1636993656
transform 1 0 69828 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_749
timestamp 25201
transform 1 0 70932 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_755
timestamp 25201
transform 1 0 71484 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_757
timestamp 1636993656
transform 1 0 71668 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_769
timestamp 1636993656
transform 1 0 72772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_781
timestamp 1636993656
transform 1 0 73876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_793
timestamp 1636993656
transform 1 0 74980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_805
timestamp 25201
transform 1 0 76084 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_811
timestamp 25201
transform 1 0 76636 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_813
timestamp 25201
transform 1 0 76820 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_821
timestamp 25201
transform 1 0 77556 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1636993656
transform 1 0 2300 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1636993656
transform 1 0 3404 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1636993656
transform 1 0 4508 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1636993656
transform 1 0 5612 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 25201
transform 1 0 6716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 25201
transform 1 0 7084 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1636993656
transform 1 0 7268 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1636993656
transform 1 0 8372 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1636993656
transform 1 0 9476 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1636993656
transform 1 0 10580 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 25201
transform 1 0 11684 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 25201
transform 1 0 12236 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1636993656
transform 1 0 12420 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1636993656
transform 1 0 13524 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1636993656
transform 1 0 14628 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1636993656
transform 1 0 15732 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 25201
transform 1 0 16836 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 25201
transform 1 0 17388 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1636993656
transform 1 0 17572 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1636993656
transform 1 0 18676 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1636993656
transform 1 0 19780 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1636993656
transform 1 0 20884 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 25201
transform 1 0 21988 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 25201
transform 1 0 22540 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1636993656
transform 1 0 22724 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1636993656
transform 1 0 23828 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1636993656
transform 1 0 24932 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1636993656
transform 1 0 26036 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 25201
transform 1 0 27140 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 25201
transform 1 0 27692 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1636993656
transform 1 0 27876 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1636993656
transform 1 0 28980 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1636993656
transform 1 0 30084 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1636993656
transform 1 0 31188 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 25201
transform 1 0 32292 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 25201
transform 1 0 32844 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1636993656
transform 1 0 33028 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1636993656
transform 1 0 34132 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1636993656
transform 1 0 35236 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1636993656
transform 1 0 36340 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 25201
transform 1 0 37444 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 25201
transform 1 0 37996 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1636993656
transform 1 0 38180 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1636993656
transform 1 0 39284 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1636993656
transform 1 0 40388 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1636993656
transform 1 0 41492 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 25201
transform 1 0 42596 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 25201
transform 1 0 43148 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1636993656
transform 1 0 43332 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1636993656
transform 1 0 44436 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1636993656
transform 1 0 45540 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1636993656
transform 1 0 46644 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 25201
transform 1 0 47748 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 25201
transform 1 0 48300 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1636993656
transform 1 0 48484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1636993656
transform 1 0 49588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1636993656
transform 1 0 50692 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1636993656
transform 1 0 51796 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 25201
transform 1 0 52900 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 25201
transform 1 0 53452 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1636993656
transform 1 0 53636 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1636993656
transform 1 0 54740 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1636993656
transform 1 0 55844 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1636993656
transform 1 0 56948 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 25201
transform 1 0 58052 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 25201
transform 1 0 58604 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_617
timestamp 1636993656
transform 1 0 58788 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_629
timestamp 1636993656
transform 1 0 59892 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_641
timestamp 1636993656
transform 1 0 60996 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_653
timestamp 1636993656
transform 1 0 62100 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 25201
transform 1 0 63204 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 25201
transform 1 0 63756 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_673
timestamp 1636993656
transform 1 0 63940 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_685
timestamp 1636993656
transform 1 0 65044 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_697
timestamp 1636993656
transform 1 0 66148 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_709
timestamp 1636993656
transform 1 0 67252 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 25201
transform 1 0 68356 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 25201
transform 1 0 68908 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_729
timestamp 1636993656
transform 1 0 69092 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_741
timestamp 1636993656
transform 1 0 70196 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_753
timestamp 1636993656
transform 1 0 71300 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_765
timestamp 1636993656
transform 1 0 72404 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_777
timestamp 25201
transform 1 0 73508 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_783
timestamp 25201
transform 1 0 74060 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_785
timestamp 1636993656
transform 1 0 74244 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_797
timestamp 1636993656
transform 1 0 75348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_809
timestamp 1636993656
transform 1 0 76452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_821
timestamp 25201
transform 1 0 77556 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636993656
transform 1 0 2300 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636993656
transform 1 0 3404 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 25201
transform 1 0 4508 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1636993656
transform 1 0 4692 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1636993656
transform 1 0 5796 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1636993656
transform 1 0 6900 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1636993656
transform 1 0 8004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 25201
transform 1 0 9108 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 25201
transform 1 0 9660 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1636993656
transform 1 0 9844 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1636993656
transform 1 0 10948 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1636993656
transform 1 0 12052 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1636993656
transform 1 0 13156 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 25201
transform 1 0 14260 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 25201
transform 1 0 14812 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1636993656
transform 1 0 14996 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1636993656
transform 1 0 16100 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1636993656
transform 1 0 17204 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1636993656
transform 1 0 18308 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 25201
transform 1 0 19412 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 25201
transform 1 0 19964 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1636993656
transform 1 0 20148 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1636993656
transform 1 0 21252 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1636993656
transform 1 0 22356 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1636993656
transform 1 0 23460 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 25201
transform 1 0 24564 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 25201
transform 1 0 25116 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1636993656
transform 1 0 25300 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1636993656
transform 1 0 26404 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1636993656
transform 1 0 27508 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1636993656
transform 1 0 28612 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 25201
transform 1 0 29716 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 25201
transform 1 0 30268 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1636993656
transform 1 0 30452 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1636993656
transform 1 0 31556 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1636993656
transform 1 0 32660 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1636993656
transform 1 0 33764 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 25201
transform 1 0 34868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 25201
transform 1 0 35420 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1636993656
transform 1 0 35604 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1636993656
transform 1 0 36708 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1636993656
transform 1 0 37812 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1636993656
transform 1 0 38916 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 25201
transform 1 0 40020 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 25201
transform 1 0 40572 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1636993656
transform 1 0 40756 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1636993656
transform 1 0 41860 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1636993656
transform 1 0 42964 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1636993656
transform 1 0 44068 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 25201
transform 1 0 45172 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 25201
transform 1 0 45724 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1636993656
transform 1 0 45908 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1636993656
transform 1 0 47012 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1636993656
transform 1 0 48116 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1636993656
transform 1 0 49220 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 25201
transform 1 0 50324 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 25201
transform 1 0 50876 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1636993656
transform 1 0 51060 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1636993656
transform 1 0 52164 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1636993656
transform 1 0 53268 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1636993656
transform 1 0 54372 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 25201
transform 1 0 55476 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 25201
transform 1 0 56028 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1636993656
transform 1 0 56212 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1636993656
transform 1 0 57316 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1636993656
transform 1 0 58420 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_625
timestamp 1636993656
transform 1 0 59524 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 25201
transform 1 0 60628 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 25201
transform 1 0 61180 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_645
timestamp 1636993656
transform 1 0 61364 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_657
timestamp 1636993656
transform 1 0 62468 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_669
timestamp 1636993656
transform 1 0 63572 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_681
timestamp 1636993656
transform 1 0 64676 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 25201
transform 1 0 65780 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 25201
transform 1 0 66332 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_701
timestamp 1636993656
transform 1 0 66516 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_713
timestamp 1636993656
transform 1 0 67620 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_725
timestamp 1636993656
transform 1 0 68724 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_737
timestamp 1636993656
transform 1 0 69828 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_749
timestamp 25201
transform 1 0 70932 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_755
timestamp 25201
transform 1 0 71484 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_757
timestamp 1636993656
transform 1 0 71668 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_769
timestamp 1636993656
transform 1 0 72772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_781
timestamp 1636993656
transform 1 0 73876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_793
timestamp 1636993656
transform 1 0 74980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_805
timestamp 25201
transform 1 0 76084 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_811
timestamp 25201
transform 1 0 76636 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_813
timestamp 25201
transform 1 0 76820 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_821
timestamp 25201
transform 1 0 77556 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636993656
transform 1 0 2300 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_15
timestamp 25201
transform 1 0 3404 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1636993656
transform 1 0 5612 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 25201
transform 1 0 6716 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 25201
transform 1 0 7084 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_57
timestamp 25201
transform 1 0 7268 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_63
timestamp 1636993656
transform 1 0 7820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_75
timestamp 25201
transform 1 0 8924 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_99
timestamp 25201
transform 1 0 11132 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 25201
transform 1 0 12144 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1636993656
transform 1 0 12420 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1636993656
transform 1 0 13524 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_137
timestamp 25201
transform 1 0 14628 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_143
timestamp 1636993656
transform 1 0 15180 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_155
timestamp 1636993656
transform 1 0 16284 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 25201
transform 1 0 17388 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_188
timestamp 1636993656
transform 1 0 19320 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_200
timestamp 1636993656
transform 1 0 20424 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_212
timestamp 25201
transform 1 0 21528 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 25201
transform 1 0 22540 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1636993656
transform 1 0 22724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_237
timestamp 25201
transform 1 0 23828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_259
timestamp 25201
transform 1 0 25852 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_263
timestamp 1636993656
transform 1 0 26220 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_275
timestamp 25201
transform 1 0 27324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 25201
transform 1 0 27692 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1636993656
transform 1 0 27876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_293
timestamp 25201
transform 1 0 28980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_299
timestamp 25201
transform 1 0 29532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_319
timestamp 1636993656
transform 1 0 31372 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_331
timestamp 25201
transform 1 0 32476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 25201
transform 1 0 32844 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 25201
transform 1 0 33028 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_348
timestamp 1636993656
transform 1 0 34040 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_360
timestamp 25201
transform 1 0 35144 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_379
timestamp 25201
transform 1 0 36892 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_383
timestamp 25201
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 25201
transform 1 0 37996 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1636993656
transform 1 0 38180 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1636993656
transform 1 0 39284 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_417
timestamp 25201
transform 1 0 40388 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_423
timestamp 1636993656
transform 1 0 40940 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_435
timestamp 1636993656
transform 1 0 42044 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 25201
transform 1 0 43148 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_449
timestamp 25201
transform 1 0 43332 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_457
timestamp 25201
transform 1 0 44068 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_479
timestamp 1636993656
transform 1 0 46092 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_491
timestamp 25201
transform 1 0 47196 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_499
timestamp 25201
transform 1 0 47932 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 25201
transform 1 0 48300 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1636993656
transform 1 0 48484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_517
timestamp 25201
transform 1 0 49588 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_539
timestamp 25201
transform 1 0 51612 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_543
timestamp 1636993656
transform 1 0 51980 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_555
timestamp 25201
transform 1 0 53084 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 25201
transform 1 0 53452 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1636993656
transform 1 0 53636 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_573
timestamp 25201
transform 1 0 54740 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_579
timestamp 25201
transform 1 0 55292 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_583
timestamp 1636993656
transform 1 0 55660 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_595
timestamp 1636993656
transform 1 0 56764 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_607
timestamp 25201
transform 1 0 57868 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_617
timestamp 25201
transform 1 0 58788 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_639
timestamp 1636993656
transform 1 0 60812 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_651
timestamp 1636993656
transform 1 0 61916 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_663
timestamp 25201
transform 1 0 63020 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 25201
transform 1 0 63756 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_673
timestamp 1636993656
transform 1 0 63940 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_685
timestamp 1636993656
transform 1 0 65044 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_697
timestamp 1636993656
transform 1 0 66148 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_709
timestamp 1636993656
transform 1 0 67252 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 25201
transform 1 0 68356 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 25201
transform 1 0 68908 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_729
timestamp 1636993656
transform 1 0 69092 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_741
timestamp 1636993656
transform 1 0 70196 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_753
timestamp 1636993656
transform 1 0 71300 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_765
timestamp 1636993656
transform 1 0 72404 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_777
timestamp 25201
transform 1 0 73508 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_783
timestamp 25201
transform 1 0 74060 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_785
timestamp 1636993656
transform 1 0 74244 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_797
timestamp 1636993656
transform 1 0 75348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_809
timestamp 1636993656
transform 1 0 76452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_821
timestamp 25201
transform 1 0 77556 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_19
timestamp 25201
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 25201
transform 1 0 4508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_29
timestamp 25201
transform 1 0 4692 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_37
timestamp 25201
transform 1 0 5428 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_57
timestamp 25201
transform 1 0 7268 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_79
timestamp 25201
transform 1 0 9292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 25201
transform 1 0 9660 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 25201
transform 1 0 9844 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_93
timestamp 25201
transform 1 0 10580 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_113
timestamp 25201
transform 1 0 12420 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_121
timestamp 25201
transform 1 0 13156 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 25201
transform 1 0 14812 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 25201
transform 1 0 14996 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_159
timestamp 25201
transform 1 0 16652 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 25201
transform 1 0 17388 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_169
timestamp 25201
transform 1 0 17572 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_177
timestamp 25201
transform 1 0 18308 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_197
timestamp 25201
transform 1 0 20148 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_219
timestamp 25201
transform 1 0 22172 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 25201
transform 1 0 22540 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_241
timestamp 25201
transform 1 0 24196 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 25201
transform 1 0 24932 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_253
timestamp 25201
transform 1 0 25300 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_261
timestamp 25201
transform 1 0 26036 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 25201
transform 1 0 27692 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 25201
transform 1 0 27876 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_299
timestamp 25201
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 25201
transform 1 0 30268 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 25201
transform 1 0 30452 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_317
timestamp 25201
transform 1 0 31188 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_337
timestamp 25201
transform 1 0 33028 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_359
timestamp 25201
transform 1 0 35052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 25201
transform 1 0 35420 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_365
timestamp 25201
transform 1 0 35604 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_373
timestamp 25201
transform 1 0 36340 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_393
timestamp 25201
transform 1 0 38180 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_401
timestamp 25201
transform 1 0 38916 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 25201
transform 1 0 40572 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_421
timestamp 25201
transform 1 0 40756 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_439
timestamp 25201
transform 1 0 42412 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_447
timestamp 25201
transform 1 0 43148 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_465
timestamp 25201
transform 1 0 44804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_473
timestamp 25201
transform 1 0 45540 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_477
timestamp 25201
transform 1 0 45908 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_499
timestamp 25201
transform 1 0 47932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_503
timestamp 25201
transform 1 0 48300 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_521
timestamp 25201
transform 1 0 49956 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_529
timestamp 25201
transform 1 0 50692 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_533
timestamp 25201
transform 1 0 51060 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_541
timestamp 25201
transform 1 0 51796 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_559
timestamp 25201
transform 1 0 53452 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_561
timestamp 25201
transform 1 0 53636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_579
timestamp 25201
transform 1 0 55292 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 25201
transform 1 0 56028 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_605
timestamp 25201
transform 1 0 57684 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_613
timestamp 25201
transform 1 0 58420 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_633
timestamp 25201
transform 1 0 60260 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_641
timestamp 25201
transform 1 0 60996 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_645
timestamp 1636993656
transform 1 0 61364 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_657
timestamp 1636993656
transform 1 0 62468 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_669
timestamp 25201
transform 1 0 63572 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_673
timestamp 1636993656
transform 1 0 63940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_685
timestamp 1636993656
transform 1 0 65044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_697
timestamp 25201
transform 1 0 66148 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_701
timestamp 1636993656
transform 1 0 66516 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_713
timestamp 1636993656
transform 1 0 67620 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_725
timestamp 25201
transform 1 0 68724 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_729
timestamp 1636993656
transform 1 0 69092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_741
timestamp 1636993656
transform 1 0 70196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_753
timestamp 25201
transform 1 0 71300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_757
timestamp 1636993656
transform 1 0 71668 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_769
timestamp 1636993656
transform 1 0 72772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_781
timestamp 25201
transform 1 0 73876 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_785
timestamp 1636993656
transform 1 0 74244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_797
timestamp 1636993656
transform 1 0 75348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_809
timestamp 25201
transform 1 0 76452 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_813
timestamp 25201
transform 1 0 76820 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_821
timestamp 25201
transform 1 0 77556 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 25201
transform 1 0 12696 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 25201
transform -1 0 26864 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 25201
transform 1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 25201
transform -1 0 34960 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 25201
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 25201
transform 1 0 23000 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 25201
transform 1 0 9016 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 25201
transform 1 0 17848 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 25201
transform 1 0 10120 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 25201
transform 1 0 35604 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 25201
transform -1 0 36708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 25201
transform 1 0 34776 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 25201
transform -1 0 48116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 25201
transform -1 0 43700 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 25201
transform -1 0 42964 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 25201
transform -1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 25201
transform 1 0 18216 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 25201
transform 1 0 16376 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 25201
transform -1 0 28612 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 25201
transform 1 0 28060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 25201
transform 1 0 21896 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 25201
transform -1 0 19320 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 25201
transform 1 0 15272 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 25201
transform 1 0 8280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 25201
transform 1 0 24472 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 25201
transform 1 0 28888 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 25201
transform -1 0 38916 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 25201
transform 1 0 21436 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 25201
transform 1 0 20608 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 25201
transform 1 0 29624 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 25201
transform 1 0 44804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 25201
transform -1 0 49956 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 25201
transform -1 0 44804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 25201
transform 1 0 8280 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 25201
transform 1 0 6440 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 25201
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 25201
transform -1 0 46644 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 25201
transform -1 0 46644 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 25201
transform -1 0 47104 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 25201
transform -1 0 31924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 25201
transform 1 0 29624 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 25201
transform -1 0 31464 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 25201
transform 1 0 40204 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 25201
transform 1 0 30728 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 25201
transform 1 0 34040 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 25201
transform -1 0 12328 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 25201
transform -1 0 11592 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 25201
transform 1 0 7544 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 25201
transform -1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 25201
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 25201
transform 1 0 10488 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 25201
transform 1 0 10488 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 25201
transform -1 0 16744 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 25201
transform 1 0 7912 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 25201
transform 1 0 25300 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 25201
transform 1 0 18584 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 25201
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 25201
transform -1 0 17112 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 25201
transform 1 0 22724 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 25201
transform 1 0 25944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 25201
transform 1 0 18952 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 25201
transform 1 0 10120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 25201
transform 1 0 14168 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 25201
transform -1 0 42228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 25201
transform -1 0 39836 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 25201
transform 1 0 34776 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 25201
transform 1 0 20700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 25201
transform -1 0 32568 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 25201
transform 1 0 32200 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 25201
transform -1 0 38916 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 25201
transform 1 0 31096 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 25201
transform -1 0 36340 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 25201
transform 1 0 17572 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 25201
transform 1 0 28152 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 25201
transform 1 0 29624 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 25201
transform -1 0 12696 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 25201
transform 1 0 11224 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 25201
transform 1 0 24196 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 25201
transform -1 0 16192 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 25201
transform 1 0 14536 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 25201
transform 1 0 17848 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 25201
transform -1 0 9752 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 25201
transform 1 0 20516 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 25201
transform 1 0 21896 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 25201
transform 1 0 47380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 25201
transform -1 0 45632 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 25201
transform 1 0 36156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 25201
transform 1 0 32200 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 25201
transform -1 0 33212 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 25201
transform 1 0 26128 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 25201
transform 1 0 24472 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 25201
transform 1 0 46644 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 25201
transform -1 0 44068 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 25201
transform -1 0 30360 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 25201
transform 1 0 31096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 25201
transform 1 0 18584 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 25201
transform 1 0 23736 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 25201
transform 1 0 28888 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 25201
transform 1 0 28152 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 25201
transform 1 0 7544 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 25201
transform 1 0 3864 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 25201
transform -1 0 15272 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 25201
transform 1 0 20424 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 25201
transform -1 0 50784 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 25201
transform -1 0 44160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 25201
transform -1 0 38088 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 25201
transform 1 0 36616 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 25201
transform 1 0 10856 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold109
timestamp 25201
transform -1 0 16376 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_12  hold110
timestamp 25201
transform -1 0 14904 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 25201
transform -1 0 42964 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 25201
transform 1 0 33304 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 25201
transform -1 0 36616 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 25201
transform 1 0 36892 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 25201
transform 1 0 13064 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 25201
transform 1 0 10488 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 25201
transform 1 0 20792 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 25201
transform 1 0 29624 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold119
timestamp 25201
transform 1 0 45908 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 25201
transform 1 0 19320 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 25201
transform -1 0 45632 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 25201
transform 1 0 28888 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold123
timestamp 25201
transform -1 0 32936 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 25201
transform -1 0 28888 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 25201
transform 1 0 21528 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold126
timestamp 25201
transform -1 0 30360 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 25201
transform -1 0 29624 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 25201
transform -1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold129
timestamp 25201
transform 1 0 28888 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 25201
transform -1 0 37352 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 25201
transform 1 0 30728 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold132
timestamp 25201
transform 1 0 38548 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 25201
transform -1 0 36524 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 25201
transform 1 0 28888 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold135
timestamp 25201
transform 1 0 36616 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 25201
transform 1 0 22264 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 25201
transform 1 0 17848 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold138
timestamp 25201
transform 1 0 26312 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 25201
transform -1 0 34776 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 25201
transform -1 0 29624 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold141
timestamp 25201
transform -1 0 35512 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 25201
transform 1 0 15640 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 25201
transform -1 0 24288 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold144
timestamp 25201
transform 1 0 22816 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 25201
transform -1 0 41492 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 25201
transform 1 0 39928 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold147
timestamp 25201
transform 1 0 43332 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 25201
transform -1 0 26312 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 25201
transform 1 0 11592 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold150
timestamp 25201
transform -1 0 25208 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 25201
transform 1 0 41124 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 25201
transform 1 0 34776 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold153
timestamp 25201
transform -1 0 38088 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 25201
transform -1 0 21160 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 25201
transform 1 0 9752 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold156
timestamp 25201
transform 1 0 20332 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 25201
transform 1 0 38916 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 25201
transform 1 0 45632 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold159
timestamp 25201
transform 1 0 46276 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 25201
transform -1 0 23736 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 25201
transform -1 0 20056 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold162
timestamp 25201
transform 1 0 18216 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 25201
transform 1 0 17112 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 25201
transform 1 0 42688 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 25201
transform 1 0 41032 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold168
timestamp 25201
transform -1 0 76728 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 25201
transform -1 0 35144 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 25201
transform -1 0 22816 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 25201
transform 1 0 15272 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 25201
transform 1 0 74520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold175
timestamp 25201
transform -1 0 76728 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 25201
transform 1 0 5336 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 25201
transform 1 0 4968 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 25201
transform 1 0 24472 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 25201
transform 1 0 22172 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 25201
transform -1 0 17848 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  hold184
timestamp 25201
transform 1 0 35604 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 25201
transform 1 0 57408 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold186
timestamp 25201
transform 1 0 58788 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  hold191
timestamp 25201
transform 1 0 52532 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 25201
transform 1 0 64768 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold193
timestamp 25201
transform 1 0 65504 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 25201
transform -1 0 19136 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 25201
transform 1 0 51336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold200
timestamp 25201
transform 1 0 52072 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 25201
transform 1 0 54372 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold207
timestamp 25201
transform 1 0 54004 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 25201
transform -1 0 68632 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold214
timestamp 25201
transform 1 0 67528 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 25201
transform 1 0 60996 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold221
timestamp 25201
transform 1 0 61732 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 25201
transform 1 0 69828 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold228
timestamp 25201
transform 1 0 69460 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 25201
transform 1 0 71392 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold235
timestamp 25201
transform -1 0 73232 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 25201
transform 1 0 6808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 25201
transform 1 0 6072 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  hold238
timestamp 25201
transform 1 0 9936 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 25201
transform 1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 25201
transform 1 0 43424 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 25201
transform -1 0 50692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold247
timestamp 25201
transform -1 0 50048 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 25201
transform -1 0 77648 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold253
timestamp 25201
transform 1 0 74704 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 25201
transform -1 0 32200 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 25201
transform 1 0 31924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 25201
transform 1 0 32660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 25201
transform 1 0 34776 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 25201
transform 1 0 30360 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 25201
transform 1 0 27876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 25201
transform -1 0 25024 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 25201
transform 1 0 17112 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 25201
transform -1 0 25208 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 25201
transform 1 0 14168 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 25201
transform -1 0 30360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 25201
transform -1 0 75256 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 25201
transform -1 0 77464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 25201
transform -1 0 77556 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold272
timestamp 25201
transform -1 0 11408 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 25201
transform 1 0 5704 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 25201
transform 1 0 8280 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 25201
transform 1 0 7912 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 25201
transform -1 0 30360 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 25201
transform 1 0 23000 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 25201
transform -1 0 28888 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 25201
transform 1 0 22724 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 25201
transform 1 0 37352 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 25201
transform -1 0 36892 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 25201
transform -1 0 34040 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 25201
transform -1 0 31740 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 25201
transform 1 0 28152 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 25201
transform -1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 25201
transform 1 0 17848 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 25201
transform -1 0 27048 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 25201
transform -1 0 27784 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 25201
transform -1 0 26312 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 25201
transform -1 0 27784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold291
timestamp 25201
transform -1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 25201
transform -1 0 35512 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 25201
transform -1 0 37076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold294
timestamp 25201
transform -1 0 37444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 25201
transform -1 0 25392 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold296
timestamp 25201
transform -1 0 24472 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold297
timestamp 25201
transform 1 0 23460 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold298
timestamp 25201
transform 1 0 13432 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 25201
transform 1 0 33304 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 25201
transform 1 0 29624 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold301
timestamp 25201
transform 1 0 25576 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold302
timestamp 25201
transform 1 0 25392 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold303
timestamp 25201
transform -1 0 41952 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 25201
transform 1 0 40388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 25201
transform -1 0 41584 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold306
timestamp 25201
transform 1 0 38180 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold307
timestamp 25201
transform -1 0 42228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold308
timestamp 25201
transform -1 0 36984 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold309
timestamp 25201
transform -1 0 25208 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 25201
transform 1 0 19688 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 25201
transform -1 0 22632 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold313
timestamp 25201
transform 1 0 39008 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 25201
transform 1 0 39928 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold315
timestamp 25201
transform 1 0 42044 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold316
timestamp 25201
transform 1 0 22724 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold317
timestamp 25201
transform 1 0 16008 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 25201
transform 1 0 10856 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd1_1  hold320
timestamp 25201
transform -1 0 15640 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold321
timestamp 25201
transform -1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold322
timestamp 25201
transform 1 0 12696 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold323
timestamp 25201
transform 1 0 33672 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 25201
transform -1 0 32476 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold325
timestamp 25201
transform -1 0 25944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold326
timestamp 25201
transform -1 0 21988 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold327
timestamp 25201
transform 1 0 14536 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold328
timestamp 25201
transform 1 0 15272 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold329
timestamp 25201
transform -1 0 15916 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold330
timestamp 25201
transform 1 0 21896 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold331
timestamp 25201
transform 1 0 13064 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold332
timestamp 25201
transform 1 0 29624 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold333
timestamp 25201
transform -1 0 31188 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold334
timestamp 25201
transform -1 0 24472 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold335
timestamp 25201
transform -1 0 34960 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold336
timestamp 25201
transform -1 0 35972 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold337
timestamp 25201
transform 1 0 25576 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold338
timestamp 25201
transform 1 0 44160 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold339
timestamp 25201
transform 1 0 35880 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold340
timestamp 25201
transform 1 0 41952 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold341
timestamp 25201
transform -1 0 27232 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold342
timestamp 25201
transform 1 0 16376 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold343
timestamp 25201
transform 1 0 11960 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold344
timestamp 25201
transform 1 0 38088 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold345
timestamp 25201
transform -1 0 29624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold346
timestamp 25201
transform -1 0 38088 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold347
timestamp 25201
transform 1 0 43700 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold348
timestamp 25201
transform 1 0 45540 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold349
timestamp 25201
transform 1 0 44620 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold350
timestamp 25201
transform -1 0 17296 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold351
timestamp 25201
transform 1 0 5704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold352
timestamp 25201
transform 1 0 10120 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold353
timestamp 25201
transform 1 0 39284 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold354
timestamp 25201
transform -1 0 41492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold355
timestamp 25201
transform -1 0 40112 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold356
timestamp 25201
transform -1 0 14904 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold357
timestamp 25201
transform -1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold358
timestamp 25201
transform -1 0 11960 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold359
timestamp 25201
transform 1 0 21712 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold360
timestamp 25201
transform 1 0 16744 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold361
timestamp 25201
transform 1 0 24472 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold362
timestamp 25201
transform -1 0 9568 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold363
timestamp 25201
transform 1 0 4232 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold364
timestamp 25201
transform 1 0 6440 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold365
timestamp 25201
transform 1 0 48300 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold366
timestamp 25201
transform -1 0 47012 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold367
timestamp 25201
transform -1 0 49220 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold368
timestamp 25201
transform 1 0 26864 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold372
timestamp 25201
transform 1 0 53636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold373
timestamp 25201
transform -1 0 56212 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold374
timestamp 25201
transform -1 0 34408 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold378
timestamp 25201
transform -1 0 58144 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold379
timestamp 25201
transform 1 0 58144 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold380
timestamp 25201
transform 1 0 9016 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold384
timestamp 25201
transform -1 0 52440 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold385
timestamp 25201
transform 1 0 52440 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold386
timestamp 25201
transform -1 0 44896 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold390
timestamp 25201
transform -1 0 65872 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold391
timestamp 25201
transform 1 0 65504 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold394
timestamp 25201
transform 1 0 18584 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold395
timestamp 25201
transform -1 0 62100 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold396
timestamp 25201
transform 1 0 62100 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold397
timestamp 25201
transform -1 0 33120 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold398
timestamp 25201
transform -1 0 27048 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold400
timestamp 25201
transform 1 0 69092 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold401
timestamp 25201
transform -1 0 71668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold405
timestamp 25201
transform 1 0 67160 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold406
timestamp 25201
transform 1 0 67528 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold410
timestamp 25201
transform -1 0 72404 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold411
timestamp 25201
transform 1 0 72404 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold412
timestamp 25201
transform 1 0 8648 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold413
timestamp 25201
transform 1 0 17480 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold414
timestamp 25201
transform 1 0 13432 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold415
timestamp 25201
transform 1 0 12696 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold418
timestamp 25201
transform 1 0 8280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold419
timestamp 25201
transform -1 0 24288 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold420
timestamp 25201
transform -1 0 16744 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold421
timestamp 25201
transform 1 0 16744 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold422
timestamp 25201
transform 1 0 24472 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold423
timestamp 25201
transform -1 0 26128 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold424
timestamp 25201
transform 1 0 14168 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold425
timestamp 25201
transform 1 0 19872 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold426
timestamp 25201
transform -1 0 19872 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold427
timestamp 25201
transform 1 0 15272 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold428
timestamp 25201
transform -1 0 27048 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold429
timestamp 25201
transform 1 0 27048 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold430
timestamp 25201
transform -1 0 45816 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold431
timestamp 25201
transform 1 0 33304 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold432
timestamp 25201
transform -1 0 40756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold433
timestamp 25201
transform 1 0 35512 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold434
timestamp 25201
transform -1 0 29624 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold435
timestamp 25201
transform -1 0 29532 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold436
timestamp 25201
transform 1 0 19320 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold437
timestamp 25201
transform -1 0 29624 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold438
timestamp 25201
transform 1 0 9384 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold439
timestamp 25201
transform 1 0 9016 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold440
timestamp 25201
transform -1 0 12328 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold441
timestamp 25201
transform -1 0 23736 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold442
timestamp 25201
transform -1 0 34040 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold443
timestamp 25201
transform -1 0 27784 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold444
timestamp 25201
transform 1 0 26404 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold445
timestamp 25201
transform 1 0 31832 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold446
timestamp 25201
transform 1 0 36616 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold447
timestamp 25201
transform -1 0 24472 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold448
timestamp 25201
transform 1 0 27140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold449
timestamp 25201
transform 1 0 34040 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold450
timestamp 25201
transform 1 0 7544 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold451
timestamp 25201
transform 1 0 4968 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold452
timestamp 25201
transform 1 0 19780 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold453
timestamp 25201
transform -1 0 21896 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold454
timestamp 25201
transform 1 0 47104 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold455
timestamp 25201
transform -1 0 48116 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold456
timestamp 25201
transform 1 0 41952 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold460
timestamp 25201
transform 1 0 48852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold461
timestamp 25201
transform 1 0 21896 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold462
timestamp 25201
transform -1 0 34224 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold463
timestamp 25201
transform -1 0 30728 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold464
timestamp 25201
transform -1 0 26680 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold465
timestamp 25201
transform -1 0 50692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold466
timestamp 25201
transform 1 0 48116 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold467
timestamp 25201
transform 1 0 30636 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold468
timestamp 25201
transform 1 0 28152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold469
timestamp 25201
transform 1 0 49956 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold470
timestamp 25201
transform -1 0 49956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold471
timestamp 25201
transform -1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold472
timestamp 25201
transform -1 0 9752 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold474
timestamp 25201
transform -1 0 20424 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold477
timestamp 25201
transform 1 0 76912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold478
timestamp 25201
transform -1 0 77648 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold479
timestamp 25201
transform 1 0 73416 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold480
timestamp 25201
transform 1 0 33304 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold481
timestamp 25201
transform -1 0 35880 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold482
timestamp 25201
transform -1 0 33304 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold483
timestamp 25201
transform -1 0 34040 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold484
timestamp 25201
transform -1 0 17480 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold485
timestamp 25201
transform 1 0 15640 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold486
timestamp 25201
transform 1 0 26312 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold487
timestamp 25201
transform 1 0 40756 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold488
timestamp 25201
transform 1 0 40480 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold489
timestamp 25201
transform -1 0 42596 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold490
timestamp 25201
transform 1 0 39652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold491
timestamp 25201
transform -1 0 40204 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold492
timestamp 25201
transform -1 0 40480 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold531
timestamp 25201
transform 1 0 18216 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold532
timestamp 25201
transform 1 0 13800 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold553
timestamp 25201
transform -1 0 38824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold554
timestamp 25201
transform -1 0 38916 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold583
timestamp 25201
transform 1 0 17664 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold584
timestamp 25201
transform -1 0 19688 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold637
timestamp 25201
transform 1 0 18584 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold638
timestamp 25201
transform 1 0 13800 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold665
timestamp 25201
transform -1 0 18952 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold666
timestamp 25201
transform -1 0 21160 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold667
timestamp 25201
transform -1 0 17480 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold695
timestamp 25201
transform -1 0 20056 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold696
timestamp 25201
transform -1 0 21896 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold697
timestamp 25201
transform -1 0 21896 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 25201
transform 1 0 9476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 25201
transform -1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 25201
transform -1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 25201
transform -1 0 35880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 25201
transform -1 0 41032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 25201
transform 1 0 45632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 25201
transform -1 0 46184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 25201
transform -1 0 3864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 25201
transform 1 0 14628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 25201
transform 1 0 22264 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 25201
transform 1 0 23460 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 25201
transform -1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 25201
transform 1 0 28612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 25201
transform 1 0 27784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 25201
transform -1 0 23000 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 25201
transform -1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 25201
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 25201
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 25201
transform -1 0 4968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 25201
transform 1 0 18952 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 25201
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 25201
transform -1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 25201
transform 1 0 41584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 25201
transform -1 0 38456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 25201
transform 1 0 45356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 25201
transform -1 0 48392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 25201
transform 1 0 48116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 25201
transform -1 0 18952 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 25201
transform 1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 25201
transform 1 0 22724 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 25201
transform -1 0 5336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 25201
transform 1 0 27508 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 25201
transform 1 0 27600 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 25201
transform -1 0 14168 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 25201
transform -1 0 25300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 25201
transform -1 0 23736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 25201
transform 1 0 12236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap103
timestamp 25201
transform -1 0 21896 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  max_cap104
timestamp 25201
transform -1 0 26128 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  output38
timestamp 25201
transform -1 0 14904 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output39
timestamp 25201
transform 1 0 36156 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output40
timestamp 25201
transform 1 0 37720 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output41
timestamp 25201
transform 1 0 39192 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output42
timestamp 25201
transform 1 0 41768 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output43
timestamp 25201
transform 1 0 43884 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output44
timestamp 25201
transform 1 0 45908 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output45
timestamp 25201
transform -1 0 49956 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output46
timestamp 25201
transform -1 0 53084 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output47
timestamp 25201
transform -1 0 55108 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output48
timestamp 25201
transform -1 0 17480 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output49
timestamp 25201
transform -1 0 58696 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output50
timestamp 25201
transform -1 0 62836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output51
timestamp 25201
transform -1 0 66424 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output52
timestamp 25201
transform -1 0 68540 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output53
timestamp 25201
transform -1 0 70564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output54
timestamp 25201
transform -1 0 73140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output55
timestamp 25201
transform 1 0 16008 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output56
timestamp 25201
transform -1 0 76268 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output57
timestamp 25201
transform 1 0 76176 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output58
timestamp 25201
transform 1 0 21896 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output59
timestamp 25201
transform 1 0 18584 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output60
timestamp 25201
transform -1 0 25208 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output61
timestamp 25201
transform 1 0 28428 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output62
timestamp 25201
transform 1 0 30452 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output63
timestamp 25201
transform -1 0 32936 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 25201
transform 1 0 34040 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 25201
transform 1 0 59340 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 25201
transform 1 0 22724 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 25201
transform 1 0 18584 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 25201
transform 1 0 15180 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 25201
transform -1 0 12328 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 25201
transform 1 0 7820 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 25201
transform -1 0 5612 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 25201
transform 1 0 56212 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 25201
transform 1 0 51980 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 25201
transform 1 0 48484 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 25201
transform 1 0 44620 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 25201
transform 1 0 40940 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 25201
transform 1 0 36616 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 25201
transform 1 0 33580 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 25201
transform 1 0 29900 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 25201
transform 1 0 26220 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 25201
transform 1 0 58788 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 25201
transform -1 0 22172 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 25201
transform -1 0 19044 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 25201
transform -1 0 14812 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 25201
transform -1 0 11132 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 25201
transform -1 0 7176 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 25201
transform -1 0 3772 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 25201
transform 1 0 53820 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 25201
transform 1 0 50140 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 25201
transform 1 0 46460 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 25201
transform 1 0 43332 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 25201
transform 1 0 39100 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 25201
transform 1 0 35420 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 25201
transform -1 0 32936 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 25201
transform -1 0 29532 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 25201
transform -1 0 25852 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_65
timestamp 25201
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 25201
transform -1 0 77924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_66
timestamp 25201
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 25201
transform -1 0 77924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_67
timestamp 25201
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 25201
transform -1 0 77924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_68
timestamp 25201
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 25201
transform -1 0 77924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_69
timestamp 25201
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 25201
transform -1 0 77924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_70
timestamp 25201
transform 1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 25201
transform -1 0 77924 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_71
timestamp 25201
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 25201
transform -1 0 77924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_72
timestamp 25201
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 25201
transform -1 0 77924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_73
timestamp 25201
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 25201
transform -1 0 77924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_74
timestamp 25201
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 25201
transform -1 0 77924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_75
timestamp 25201
transform 1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 25201
transform -1 0 77924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_76
timestamp 25201
transform 1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 25201
transform -1 0 77924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_77
timestamp 25201
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 25201
transform -1 0 77924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_78
timestamp 25201
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 25201
transform -1 0 77924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_79
timestamp 25201
transform 1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 25201
transform -1 0 77924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_80
timestamp 25201
transform 1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 25201
transform -1 0 77924 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_81
timestamp 25201
transform 1 0 2024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 25201
transform -1 0 77924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_82
timestamp 25201
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 25201
transform -1 0 77924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_83
timestamp 25201
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 25201
transform -1 0 77924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_84
timestamp 25201
transform 1 0 2024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 25201
transform -1 0 77924 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_85
timestamp 25201
transform 1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 25201
transform -1 0 77924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_86
timestamp 25201
transform 1 0 2024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 25201
transform -1 0 77924 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_87
timestamp 25201
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 25201
transform -1 0 77924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_88
timestamp 25201
transform 1 0 2024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 25201
transform -1 0 77924 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_89
timestamp 25201
transform 1 0 2024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 25201
transform -1 0 77924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_90
timestamp 25201
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 25201
transform -1 0 77924 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_91
timestamp 25201
transform 1 0 2024 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 25201
transform -1 0 77924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_92
timestamp 25201
transform 1 0 2024 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 25201
transform -1 0 77924 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_93
timestamp 25201
transform 1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 25201
transform -1 0 77924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_94
timestamp 25201
transform 1 0 2024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 25201
transform -1 0 77924 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_95
timestamp 25201
transform 1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 25201
transform -1 0 77924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_96
timestamp 25201
transform 1 0 2024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 25201
transform -1 0 77924 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_97
timestamp 25201
transform 1 0 2024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 25201
transform -1 0 77924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_98
timestamp 25201
transform 1 0 2024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 25201
transform -1 0 77924 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_99
timestamp 25201
transform 1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 25201
transform -1 0 77924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_100
timestamp 25201
transform 1 0 2024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 25201
transform -1 0 77924 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_101
timestamp 25201
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 25201
transform -1 0 77924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_102
timestamp 25201
transform 1 0 2024 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 25201
transform -1 0 77924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_103
timestamp 25201
transform 1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 25201
transform -1 0 77924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_104
timestamp 25201
transform 1 0 2024 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 25201
transform -1 0 77924 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_105
timestamp 25201
transform 1 0 2024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 25201
transform -1 0 77924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_106
timestamp 25201
transform 1 0 2024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 25201
transform -1 0 77924 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_107
timestamp 25201
transform 1 0 2024 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 25201
transform -1 0 77924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_108
timestamp 25201
transform 1 0 2024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 25201
transform -1 0 77924 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_109
timestamp 25201
transform 1 0 2024 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 25201
transform -1 0 77924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_110
timestamp 25201
transform 1 0 2024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 25201
transform -1 0 77924 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_111
timestamp 25201
transform 1 0 2024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 25201
transform -1 0 77924 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_112
timestamp 25201
transform 1 0 2024 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 25201
transform -1 0 77924 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_113
timestamp 25201
transform 1 0 2024 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 25201
transform -1 0 77924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_114
timestamp 25201
transform 1 0 2024 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 25201
transform -1 0 77924 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_115
timestamp 25201
transform 1 0 2024 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 25201
transform -1 0 77924 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_116
timestamp 25201
transform 1 0 2024 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 25201
transform -1 0 77924 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_117
timestamp 25201
transform 1 0 2024 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 25201
transform -1 0 77924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_118
timestamp 25201
transform 1 0 2024 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 25201
transform -1 0 77924 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_119
timestamp 25201
transform 1 0 2024 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 25201
transform -1 0 77924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_120
timestamp 25201
transform 1 0 2024 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 25201
transform -1 0 77924 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_121
timestamp 25201
transform 1 0 2024 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 25201
transform -1 0 77924 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_122
timestamp 25201
transform 1 0 2024 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 25201
transform -1 0 77924 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_123
timestamp 25201
transform 1 0 2024 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 25201
transform -1 0 77924 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_124
timestamp 25201
transform 1 0 2024 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 25201
transform -1 0 77924 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_125
timestamp 25201
transform 1 0 2024 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 25201
transform -1 0 77924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_126
timestamp 25201
transform 1 0 2024 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 25201
transform -1 0 77924 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_127
timestamp 25201
transform 1 0 2024 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 25201
transform -1 0 77924 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_128
timestamp 25201
transform 1 0 2024 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 25201
transform -1 0 77924 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_129
timestamp 25201
transform 1 0 2024 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 25201
transform -1 0 77924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_130
timestamp 25201
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_131
timestamp 25201
transform 1 0 7176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp 25201
transform 1 0 9752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp 25201
transform 1 0 12328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp 25201
transform 1 0 14904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp 25201
transform 1 0 17480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp 25201
transform 1 0 20056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_137
timestamp 25201
transform 1 0 22632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138
timestamp 25201
transform 1 0 25208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 25201
transform 1 0 27784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 25201
transform 1 0 30360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 25201
transform 1 0 32936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 25201
transform 1 0 35512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_143
timestamp 25201
transform 1 0 38088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_144
timestamp 25201
transform 1 0 40664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_145
timestamp 25201
transform 1 0 43240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_146
timestamp 25201
transform 1 0 45816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_147
timestamp 25201
transform 1 0 48392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_148
timestamp 25201
transform 1 0 50968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_149
timestamp 25201
transform 1 0 53544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_150
timestamp 25201
transform 1 0 56120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_151
timestamp 25201
transform 1 0 58696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_152
timestamp 25201
transform 1 0 61272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_153
timestamp 25201
transform 1 0 63848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_154
timestamp 25201
transform 1 0 66424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_155
timestamp 25201
transform 1 0 69000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_156
timestamp 25201
transform 1 0 71576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_157
timestamp 25201
transform 1 0 74152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_158
timestamp 25201
transform 1 0 76728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_159
timestamp 25201
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_160
timestamp 25201
transform 1 0 12328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_161
timestamp 25201
transform 1 0 17480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_162
timestamp 25201
transform 1 0 22632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_163
timestamp 25201
transform 1 0 27784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_164
timestamp 25201
transform 1 0 32936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_165
timestamp 25201
transform 1 0 38088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_166
timestamp 25201
transform 1 0 43240 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_167
timestamp 25201
transform 1 0 48392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_168
timestamp 25201
transform 1 0 53544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_169
timestamp 25201
transform 1 0 58696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_170
timestamp 25201
transform 1 0 63848 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_171
timestamp 25201
transform 1 0 69000 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_172
timestamp 25201
transform 1 0 74152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_173
timestamp 25201
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_174
timestamp 25201
transform 1 0 9752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_175
timestamp 25201
transform 1 0 14904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_176
timestamp 25201
transform 1 0 20056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_177
timestamp 25201
transform 1 0 25208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_178
timestamp 25201
transform 1 0 30360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_179
timestamp 25201
transform 1 0 35512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_180
timestamp 25201
transform 1 0 40664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_181
timestamp 25201
transform 1 0 45816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_182
timestamp 25201
transform 1 0 50968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_183
timestamp 25201
transform 1 0 56120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_184
timestamp 25201
transform 1 0 61272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_185
timestamp 25201
transform 1 0 66424 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_186
timestamp 25201
transform 1 0 71576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_187
timestamp 25201
transform 1 0 76728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_188
timestamp 25201
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_189
timestamp 25201
transform 1 0 12328 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_190
timestamp 25201
transform 1 0 17480 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_191
timestamp 25201
transform 1 0 22632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_192
timestamp 25201
transform 1 0 27784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_193
timestamp 25201
transform 1 0 32936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_194
timestamp 25201
transform 1 0 38088 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_195
timestamp 25201
transform 1 0 43240 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_196
timestamp 25201
transform 1 0 48392 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_197
timestamp 25201
transform 1 0 53544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_198
timestamp 25201
transform 1 0 58696 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_199
timestamp 25201
transform 1 0 63848 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_200
timestamp 25201
transform 1 0 69000 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_201
timestamp 25201
transform 1 0 74152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_202
timestamp 25201
transform 1 0 4600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_203
timestamp 25201
transform 1 0 9752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_204
timestamp 25201
transform 1 0 14904 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_205
timestamp 25201
transform 1 0 20056 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_206
timestamp 25201
transform 1 0 25208 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_207
timestamp 25201
transform 1 0 30360 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_208
timestamp 25201
transform 1 0 35512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_209
timestamp 25201
transform 1 0 40664 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_210
timestamp 25201
transform 1 0 45816 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_211
timestamp 25201
transform 1 0 50968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_212
timestamp 25201
transform 1 0 56120 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_213
timestamp 25201
transform 1 0 61272 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_214
timestamp 25201
transform 1 0 66424 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_215
timestamp 25201
transform 1 0 71576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_216
timestamp 25201
transform 1 0 76728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_217
timestamp 25201
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_218
timestamp 25201
transform 1 0 12328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_219
timestamp 25201
transform 1 0 17480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_220
timestamp 25201
transform 1 0 22632 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_221
timestamp 25201
transform 1 0 27784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_222
timestamp 25201
transform 1 0 32936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_223
timestamp 25201
transform 1 0 38088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_224
timestamp 25201
transform 1 0 43240 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_225
timestamp 25201
transform 1 0 48392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_226
timestamp 25201
transform 1 0 53544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_227
timestamp 25201
transform 1 0 58696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_228
timestamp 25201
transform 1 0 63848 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_229
timestamp 25201
transform 1 0 69000 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_230
timestamp 25201
transform 1 0 74152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_231
timestamp 25201
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_232
timestamp 25201
transform 1 0 9752 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_233
timestamp 25201
transform 1 0 14904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_234
timestamp 25201
transform 1 0 20056 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_235
timestamp 25201
transform 1 0 25208 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_236
timestamp 25201
transform 1 0 30360 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_237
timestamp 25201
transform 1 0 35512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_238
timestamp 25201
transform 1 0 40664 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_239
timestamp 25201
transform 1 0 45816 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_240
timestamp 25201
transform 1 0 50968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_241
timestamp 25201
transform 1 0 56120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_242
timestamp 25201
transform 1 0 61272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_243
timestamp 25201
transform 1 0 66424 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_244
timestamp 25201
transform 1 0 71576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_245
timestamp 25201
transform 1 0 76728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_246
timestamp 25201
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_247
timestamp 25201
transform 1 0 12328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_248
timestamp 25201
transform 1 0 17480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_249
timestamp 25201
transform 1 0 22632 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_250
timestamp 25201
transform 1 0 27784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_251
timestamp 25201
transform 1 0 32936 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_252
timestamp 25201
transform 1 0 38088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_253
timestamp 25201
transform 1 0 43240 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_254
timestamp 25201
transform 1 0 48392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_255
timestamp 25201
transform 1 0 53544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_256
timestamp 25201
transform 1 0 58696 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_257
timestamp 25201
transform 1 0 63848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_258
timestamp 25201
transform 1 0 69000 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_259
timestamp 25201
transform 1 0 74152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_260
timestamp 25201
transform 1 0 4600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_261
timestamp 25201
transform 1 0 9752 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_262
timestamp 25201
transform 1 0 14904 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_263
timestamp 25201
transform 1 0 20056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_264
timestamp 25201
transform 1 0 25208 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_265
timestamp 25201
transform 1 0 30360 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_266
timestamp 25201
transform 1 0 35512 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_267
timestamp 25201
transform 1 0 40664 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_268
timestamp 25201
transform 1 0 45816 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_269
timestamp 25201
transform 1 0 50968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_270
timestamp 25201
transform 1 0 56120 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_271
timestamp 25201
transform 1 0 61272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_272
timestamp 25201
transform 1 0 66424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_273
timestamp 25201
transform 1 0 71576 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_274
timestamp 25201
transform 1 0 76728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_275
timestamp 25201
transform 1 0 7176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_276
timestamp 25201
transform 1 0 12328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_277
timestamp 25201
transform 1 0 17480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_278
timestamp 25201
transform 1 0 22632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_279
timestamp 25201
transform 1 0 27784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_280
timestamp 25201
transform 1 0 32936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_281
timestamp 25201
transform 1 0 38088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_282
timestamp 25201
transform 1 0 43240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_283
timestamp 25201
transform 1 0 48392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_284
timestamp 25201
transform 1 0 53544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_285
timestamp 25201
transform 1 0 58696 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_286
timestamp 25201
transform 1 0 63848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_287
timestamp 25201
transform 1 0 69000 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_288
timestamp 25201
transform 1 0 74152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_289
timestamp 25201
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_290
timestamp 25201
transform 1 0 9752 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_291
timestamp 25201
transform 1 0 14904 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_292
timestamp 25201
transform 1 0 20056 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_293
timestamp 25201
transform 1 0 25208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_294
timestamp 25201
transform 1 0 30360 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_295
timestamp 25201
transform 1 0 35512 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_296
timestamp 25201
transform 1 0 40664 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_297
timestamp 25201
transform 1 0 45816 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_298
timestamp 25201
transform 1 0 50968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_299
timestamp 25201
transform 1 0 56120 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_300
timestamp 25201
transform 1 0 61272 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_301
timestamp 25201
transform 1 0 66424 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_302
timestamp 25201
transform 1 0 71576 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_303
timestamp 25201
transform 1 0 76728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_304
timestamp 25201
transform 1 0 7176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_305
timestamp 25201
transform 1 0 12328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_306
timestamp 25201
transform 1 0 17480 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_307
timestamp 25201
transform 1 0 22632 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_308
timestamp 25201
transform 1 0 27784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_309
timestamp 25201
transform 1 0 32936 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_310
timestamp 25201
transform 1 0 38088 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_311
timestamp 25201
transform 1 0 43240 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_312
timestamp 25201
transform 1 0 48392 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_313
timestamp 25201
transform 1 0 53544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_314
timestamp 25201
transform 1 0 58696 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_315
timestamp 25201
transform 1 0 63848 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_316
timestamp 25201
transform 1 0 69000 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_317
timestamp 25201
transform 1 0 74152 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_318
timestamp 25201
transform 1 0 4600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_319
timestamp 25201
transform 1 0 9752 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_320
timestamp 25201
transform 1 0 14904 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_321
timestamp 25201
transform 1 0 20056 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_322
timestamp 25201
transform 1 0 25208 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_323
timestamp 25201
transform 1 0 30360 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_324
timestamp 25201
transform 1 0 35512 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_325
timestamp 25201
transform 1 0 40664 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_326
timestamp 25201
transform 1 0 45816 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_327
timestamp 25201
transform 1 0 50968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_328
timestamp 25201
transform 1 0 56120 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_329
timestamp 25201
transform 1 0 61272 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_330
timestamp 25201
transform 1 0 66424 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_331
timestamp 25201
transform 1 0 71576 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_332
timestamp 25201
transform 1 0 76728 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_333
timestamp 25201
transform 1 0 7176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_334
timestamp 25201
transform 1 0 12328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_335
timestamp 25201
transform 1 0 17480 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_336
timestamp 25201
transform 1 0 22632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_337
timestamp 25201
transform 1 0 27784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_338
timestamp 25201
transform 1 0 32936 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_339
timestamp 25201
transform 1 0 38088 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_340
timestamp 25201
transform 1 0 43240 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_341
timestamp 25201
transform 1 0 48392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_342
timestamp 25201
transform 1 0 53544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_343
timestamp 25201
transform 1 0 58696 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_344
timestamp 25201
transform 1 0 63848 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_345
timestamp 25201
transform 1 0 69000 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_346
timestamp 25201
transform 1 0 74152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_347
timestamp 25201
transform 1 0 4600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_348
timestamp 25201
transform 1 0 9752 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_349
timestamp 25201
transform 1 0 14904 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_350
timestamp 25201
transform 1 0 20056 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_351
timestamp 25201
transform 1 0 25208 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_352
timestamp 25201
transform 1 0 30360 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_353
timestamp 25201
transform 1 0 35512 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_354
timestamp 25201
transform 1 0 40664 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_355
timestamp 25201
transform 1 0 45816 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_356
timestamp 25201
transform 1 0 50968 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_357
timestamp 25201
transform 1 0 56120 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_358
timestamp 25201
transform 1 0 61272 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_359
timestamp 25201
transform 1 0 66424 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_360
timestamp 25201
transform 1 0 71576 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_361
timestamp 25201
transform 1 0 76728 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_362
timestamp 25201
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_363
timestamp 25201
transform 1 0 12328 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_364
timestamp 25201
transform 1 0 17480 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_365
timestamp 25201
transform 1 0 22632 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_366
timestamp 25201
transform 1 0 27784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_367
timestamp 25201
transform 1 0 32936 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_368
timestamp 25201
transform 1 0 38088 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_369
timestamp 25201
transform 1 0 43240 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_370
timestamp 25201
transform 1 0 48392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_371
timestamp 25201
transform 1 0 53544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_372
timestamp 25201
transform 1 0 58696 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_373
timestamp 25201
transform 1 0 63848 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_374
timestamp 25201
transform 1 0 69000 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_375
timestamp 25201
transform 1 0 74152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_376
timestamp 25201
transform 1 0 4600 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_377
timestamp 25201
transform 1 0 9752 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_378
timestamp 25201
transform 1 0 14904 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_379
timestamp 25201
transform 1 0 20056 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_380
timestamp 25201
transform 1 0 25208 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_381
timestamp 25201
transform 1 0 30360 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_382
timestamp 25201
transform 1 0 35512 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_383
timestamp 25201
transform 1 0 40664 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_384
timestamp 25201
transform 1 0 45816 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_385
timestamp 25201
transform 1 0 50968 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_386
timestamp 25201
transform 1 0 56120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_387
timestamp 25201
transform 1 0 61272 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_388
timestamp 25201
transform 1 0 66424 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_389
timestamp 25201
transform 1 0 71576 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_390
timestamp 25201
transform 1 0 76728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_391
timestamp 25201
transform 1 0 7176 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_392
timestamp 25201
transform 1 0 12328 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_393
timestamp 25201
transform 1 0 17480 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_394
timestamp 25201
transform 1 0 22632 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_395
timestamp 25201
transform 1 0 27784 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_396
timestamp 25201
transform 1 0 32936 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_397
timestamp 25201
transform 1 0 38088 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_398
timestamp 25201
transform 1 0 43240 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_399
timestamp 25201
transform 1 0 48392 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_400
timestamp 25201
transform 1 0 53544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_401
timestamp 25201
transform 1 0 58696 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_402
timestamp 25201
transform 1 0 63848 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_403
timestamp 25201
transform 1 0 69000 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_404
timestamp 25201
transform 1 0 74152 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_405
timestamp 25201
transform 1 0 4600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_406
timestamp 25201
transform 1 0 9752 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_407
timestamp 25201
transform 1 0 14904 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_408
timestamp 25201
transform 1 0 20056 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_409
timestamp 25201
transform 1 0 25208 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_410
timestamp 25201
transform 1 0 30360 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_411
timestamp 25201
transform 1 0 35512 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_412
timestamp 25201
transform 1 0 40664 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_413
timestamp 25201
transform 1 0 45816 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_414
timestamp 25201
transform 1 0 50968 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_415
timestamp 25201
transform 1 0 56120 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_416
timestamp 25201
transform 1 0 61272 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_417
timestamp 25201
transform 1 0 66424 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_418
timestamp 25201
transform 1 0 71576 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_419
timestamp 25201
transform 1 0 76728 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_420
timestamp 25201
transform 1 0 7176 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_421
timestamp 25201
transform 1 0 12328 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_422
timestamp 25201
transform 1 0 17480 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_423
timestamp 25201
transform 1 0 22632 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_424
timestamp 25201
transform 1 0 27784 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_425
timestamp 25201
transform 1 0 32936 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_426
timestamp 25201
transform 1 0 38088 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_427
timestamp 25201
transform 1 0 43240 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_428
timestamp 25201
transform 1 0 48392 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_429
timestamp 25201
transform 1 0 53544 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_430
timestamp 25201
transform 1 0 58696 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_431
timestamp 25201
transform 1 0 63848 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_432
timestamp 25201
transform 1 0 69000 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_433
timestamp 25201
transform 1 0 74152 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_434
timestamp 25201
transform 1 0 4600 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_435
timestamp 25201
transform 1 0 9752 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_436
timestamp 25201
transform 1 0 14904 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_437
timestamp 25201
transform 1 0 20056 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_438
timestamp 25201
transform 1 0 25208 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_439
timestamp 25201
transform 1 0 30360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_440
timestamp 25201
transform 1 0 35512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_441
timestamp 25201
transform 1 0 40664 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_442
timestamp 25201
transform 1 0 45816 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_443
timestamp 25201
transform 1 0 50968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_444
timestamp 25201
transform 1 0 56120 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_445
timestamp 25201
transform 1 0 61272 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_446
timestamp 25201
transform 1 0 66424 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_447
timestamp 25201
transform 1 0 71576 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_448
timestamp 25201
transform 1 0 76728 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_449
timestamp 25201
transform 1 0 7176 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_450
timestamp 25201
transform 1 0 12328 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_451
timestamp 25201
transform 1 0 17480 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_452
timestamp 25201
transform 1 0 22632 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_453
timestamp 25201
transform 1 0 27784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_454
timestamp 25201
transform 1 0 32936 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_455
timestamp 25201
transform 1 0 38088 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_456
timestamp 25201
transform 1 0 43240 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_457
timestamp 25201
transform 1 0 48392 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_458
timestamp 25201
transform 1 0 53544 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_459
timestamp 25201
transform 1 0 58696 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_460
timestamp 25201
transform 1 0 63848 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_461
timestamp 25201
transform 1 0 69000 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_462
timestamp 25201
transform 1 0 74152 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_463
timestamp 25201
transform 1 0 4600 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_464
timestamp 25201
transform 1 0 9752 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_465
timestamp 25201
transform 1 0 14904 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_466
timestamp 25201
transform 1 0 20056 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_467
timestamp 25201
transform 1 0 25208 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_468
timestamp 25201
transform 1 0 30360 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_469
timestamp 25201
transform 1 0 35512 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_470
timestamp 25201
transform 1 0 40664 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_471
timestamp 25201
transform 1 0 45816 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_472
timestamp 25201
transform 1 0 50968 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_473
timestamp 25201
transform 1 0 56120 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_474
timestamp 25201
transform 1 0 61272 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_475
timestamp 25201
transform 1 0 66424 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_476
timestamp 25201
transform 1 0 71576 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_477
timestamp 25201
transform 1 0 76728 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_478
timestamp 25201
transform 1 0 7176 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_479
timestamp 25201
transform 1 0 12328 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_480
timestamp 25201
transform 1 0 17480 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_481
timestamp 25201
transform 1 0 22632 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_482
timestamp 25201
transform 1 0 27784 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_483
timestamp 25201
transform 1 0 32936 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_484
timestamp 25201
transform 1 0 38088 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_485
timestamp 25201
transform 1 0 43240 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_486
timestamp 25201
transform 1 0 48392 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_487
timestamp 25201
transform 1 0 53544 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_488
timestamp 25201
transform 1 0 58696 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_489
timestamp 25201
transform 1 0 63848 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_490
timestamp 25201
transform 1 0 69000 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_491
timestamp 25201
transform 1 0 74152 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_492
timestamp 25201
transform 1 0 4600 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_493
timestamp 25201
transform 1 0 9752 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_494
timestamp 25201
transform 1 0 14904 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_495
timestamp 25201
transform 1 0 20056 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_496
timestamp 25201
transform 1 0 25208 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_497
timestamp 25201
transform 1 0 30360 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_498
timestamp 25201
transform 1 0 35512 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_499
timestamp 25201
transform 1 0 40664 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_500
timestamp 25201
transform 1 0 45816 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_501
timestamp 25201
transform 1 0 50968 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_502
timestamp 25201
transform 1 0 56120 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_503
timestamp 25201
transform 1 0 61272 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_504
timestamp 25201
transform 1 0 66424 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_505
timestamp 25201
transform 1 0 71576 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_506
timestamp 25201
transform 1 0 76728 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_507
timestamp 25201
transform 1 0 7176 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_508
timestamp 25201
transform 1 0 12328 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_509
timestamp 25201
transform 1 0 17480 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_510
timestamp 25201
transform 1 0 22632 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_511
timestamp 25201
transform 1 0 27784 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_512
timestamp 25201
transform 1 0 32936 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_513
timestamp 25201
transform 1 0 38088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_514
timestamp 25201
transform 1 0 43240 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_515
timestamp 25201
transform 1 0 48392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_516
timestamp 25201
transform 1 0 53544 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_517
timestamp 25201
transform 1 0 58696 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_518
timestamp 25201
transform 1 0 63848 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_519
timestamp 25201
transform 1 0 69000 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_520
timestamp 25201
transform 1 0 74152 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_521
timestamp 25201
transform 1 0 4600 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_522
timestamp 25201
transform 1 0 9752 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_523
timestamp 25201
transform 1 0 14904 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_524
timestamp 25201
transform 1 0 20056 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_525
timestamp 25201
transform 1 0 25208 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_526
timestamp 25201
transform 1 0 30360 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_527
timestamp 25201
transform 1 0 35512 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_528
timestamp 25201
transform 1 0 40664 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_529
timestamp 25201
transform 1 0 45816 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_530
timestamp 25201
transform 1 0 50968 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_531
timestamp 25201
transform 1 0 56120 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_532
timestamp 25201
transform 1 0 61272 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_533
timestamp 25201
transform 1 0 66424 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_534
timestamp 25201
transform 1 0 71576 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_535
timestamp 25201
transform 1 0 76728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_536
timestamp 25201
transform 1 0 7176 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_537
timestamp 25201
transform 1 0 12328 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_538
timestamp 25201
transform 1 0 17480 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_539
timestamp 25201
transform 1 0 22632 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_540
timestamp 25201
transform 1 0 27784 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_541
timestamp 25201
transform 1 0 32936 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_542
timestamp 25201
transform 1 0 38088 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_543
timestamp 25201
transform 1 0 43240 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_544
timestamp 25201
transform 1 0 48392 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_545
timestamp 25201
transform 1 0 53544 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_546
timestamp 25201
transform 1 0 58696 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_547
timestamp 25201
transform 1 0 63848 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_548
timestamp 25201
transform 1 0 69000 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_549
timestamp 25201
transform 1 0 74152 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_550
timestamp 25201
transform 1 0 4600 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_551
timestamp 25201
transform 1 0 9752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_552
timestamp 25201
transform 1 0 14904 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_553
timestamp 25201
transform 1 0 20056 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_554
timestamp 25201
transform 1 0 25208 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_555
timestamp 25201
transform 1 0 30360 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_556
timestamp 25201
transform 1 0 35512 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_557
timestamp 25201
transform 1 0 40664 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_558
timestamp 25201
transform 1 0 45816 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_559
timestamp 25201
transform 1 0 50968 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_560
timestamp 25201
transform 1 0 56120 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_561
timestamp 25201
transform 1 0 61272 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_562
timestamp 25201
transform 1 0 66424 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_563
timestamp 25201
transform 1 0 71576 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_564
timestamp 25201
transform 1 0 76728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_565
timestamp 25201
transform 1 0 7176 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_566
timestamp 25201
transform 1 0 12328 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_567
timestamp 25201
transform 1 0 17480 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_568
timestamp 25201
transform 1 0 22632 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_569
timestamp 25201
transform 1 0 27784 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_570
timestamp 25201
transform 1 0 32936 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_571
timestamp 25201
transform 1 0 38088 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_572
timestamp 25201
transform 1 0 43240 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_573
timestamp 25201
transform 1 0 48392 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_574
timestamp 25201
transform 1 0 53544 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_575
timestamp 25201
transform 1 0 58696 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_576
timestamp 25201
transform 1 0 63848 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_577
timestamp 25201
transform 1 0 69000 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_578
timestamp 25201
transform 1 0 74152 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_579
timestamp 25201
transform 1 0 4600 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_580
timestamp 25201
transform 1 0 9752 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_581
timestamp 25201
transform 1 0 14904 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_582
timestamp 25201
transform 1 0 20056 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_583
timestamp 25201
transform 1 0 25208 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_584
timestamp 25201
transform 1 0 30360 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_585
timestamp 25201
transform 1 0 35512 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_586
timestamp 25201
transform 1 0 40664 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_587
timestamp 25201
transform 1 0 45816 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_588
timestamp 25201
transform 1 0 50968 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_589
timestamp 25201
transform 1 0 56120 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_590
timestamp 25201
transform 1 0 61272 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_591
timestamp 25201
transform 1 0 66424 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_592
timestamp 25201
transform 1 0 71576 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_593
timestamp 25201
transform 1 0 76728 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_594
timestamp 25201
transform 1 0 7176 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_595
timestamp 25201
transform 1 0 12328 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_596
timestamp 25201
transform 1 0 17480 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_597
timestamp 25201
transform 1 0 22632 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_598
timestamp 25201
transform 1 0 27784 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_599
timestamp 25201
transform 1 0 32936 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_600
timestamp 25201
transform 1 0 38088 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_601
timestamp 25201
transform 1 0 43240 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_602
timestamp 25201
transform 1 0 48392 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_603
timestamp 25201
transform 1 0 53544 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_604
timestamp 25201
transform 1 0 58696 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_605
timestamp 25201
transform 1 0 63848 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_606
timestamp 25201
transform 1 0 69000 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_607
timestamp 25201
transform 1 0 74152 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_608
timestamp 25201
transform 1 0 4600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_609
timestamp 25201
transform 1 0 9752 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_610
timestamp 25201
transform 1 0 14904 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_611
timestamp 25201
transform 1 0 20056 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_612
timestamp 25201
transform 1 0 25208 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_613
timestamp 25201
transform 1 0 30360 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_614
timestamp 25201
transform 1 0 35512 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_615
timestamp 25201
transform 1 0 40664 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_616
timestamp 25201
transform 1 0 45816 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_617
timestamp 25201
transform 1 0 50968 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_618
timestamp 25201
transform 1 0 56120 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_619
timestamp 25201
transform 1 0 61272 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_620
timestamp 25201
transform 1 0 66424 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_621
timestamp 25201
transform 1 0 71576 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_622
timestamp 25201
transform 1 0 76728 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_623
timestamp 25201
transform 1 0 7176 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_624
timestamp 25201
transform 1 0 12328 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_625
timestamp 25201
transform 1 0 17480 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_626
timestamp 25201
transform 1 0 22632 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_627
timestamp 25201
transform 1 0 27784 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_628
timestamp 25201
transform 1 0 32936 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_629
timestamp 25201
transform 1 0 38088 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_630
timestamp 25201
transform 1 0 43240 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_631
timestamp 25201
transform 1 0 48392 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_632
timestamp 25201
transform 1 0 53544 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_633
timestamp 25201
transform 1 0 58696 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_634
timestamp 25201
transform 1 0 63848 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_635
timestamp 25201
transform 1 0 69000 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_636
timestamp 25201
transform 1 0 74152 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_637
timestamp 25201
transform 1 0 4600 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_638
timestamp 25201
transform 1 0 9752 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_639
timestamp 25201
transform 1 0 14904 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_640
timestamp 25201
transform 1 0 20056 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_641
timestamp 25201
transform 1 0 25208 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_642
timestamp 25201
transform 1 0 30360 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_643
timestamp 25201
transform 1 0 35512 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_644
timestamp 25201
transform 1 0 40664 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_645
timestamp 25201
transform 1 0 45816 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_646
timestamp 25201
transform 1 0 50968 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_647
timestamp 25201
transform 1 0 56120 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_648
timestamp 25201
transform 1 0 61272 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_649
timestamp 25201
transform 1 0 66424 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_650
timestamp 25201
transform 1 0 71576 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_651
timestamp 25201
transform 1 0 76728 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_652
timestamp 25201
transform 1 0 7176 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_653
timestamp 25201
transform 1 0 12328 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_654
timestamp 25201
transform 1 0 17480 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_655
timestamp 25201
transform 1 0 22632 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_656
timestamp 25201
transform 1 0 27784 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_657
timestamp 25201
transform 1 0 32936 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_658
timestamp 25201
transform 1 0 38088 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_659
timestamp 25201
transform 1 0 43240 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_660
timestamp 25201
transform 1 0 48392 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_661
timestamp 25201
transform 1 0 53544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_662
timestamp 25201
transform 1 0 58696 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_663
timestamp 25201
transform 1 0 63848 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_664
timestamp 25201
transform 1 0 69000 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_665
timestamp 25201
transform 1 0 74152 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_666
timestamp 25201
transform 1 0 4600 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_667
timestamp 25201
transform 1 0 9752 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_668
timestamp 25201
transform 1 0 14904 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_669
timestamp 25201
transform 1 0 20056 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_670
timestamp 25201
transform 1 0 25208 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_671
timestamp 25201
transform 1 0 30360 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_672
timestamp 25201
transform 1 0 35512 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_673
timestamp 25201
transform 1 0 40664 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_674
timestamp 25201
transform 1 0 45816 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_675
timestamp 25201
transform 1 0 50968 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_676
timestamp 25201
transform 1 0 56120 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_677
timestamp 25201
transform 1 0 61272 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_678
timestamp 25201
transform 1 0 66424 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_679
timestamp 25201
transform 1 0 71576 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_680
timestamp 25201
transform 1 0 76728 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_681
timestamp 25201
transform 1 0 7176 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_682
timestamp 25201
transform 1 0 12328 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_683
timestamp 25201
transform 1 0 17480 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_684
timestamp 25201
transform 1 0 22632 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_685
timestamp 25201
transform 1 0 27784 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_686
timestamp 25201
transform 1 0 32936 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_687
timestamp 25201
transform 1 0 38088 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_688
timestamp 25201
transform 1 0 43240 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_689
timestamp 25201
transform 1 0 48392 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_690
timestamp 25201
transform 1 0 53544 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_691
timestamp 25201
transform 1 0 58696 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_692
timestamp 25201
transform 1 0 63848 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_693
timestamp 25201
transform 1 0 69000 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_694
timestamp 25201
transform 1 0 74152 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_695
timestamp 25201
transform 1 0 4600 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_696
timestamp 25201
transform 1 0 9752 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_697
timestamp 25201
transform 1 0 14904 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_698
timestamp 25201
transform 1 0 20056 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_699
timestamp 25201
transform 1 0 25208 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_700
timestamp 25201
transform 1 0 30360 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_701
timestamp 25201
transform 1 0 35512 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_702
timestamp 25201
transform 1 0 40664 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_703
timestamp 25201
transform 1 0 45816 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_704
timestamp 25201
transform 1 0 50968 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_705
timestamp 25201
transform 1 0 56120 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_706
timestamp 25201
transform 1 0 61272 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_707
timestamp 25201
transform 1 0 66424 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_708
timestamp 25201
transform 1 0 71576 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_709
timestamp 25201
transform 1 0 76728 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_710
timestamp 25201
transform 1 0 7176 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_711
timestamp 25201
transform 1 0 12328 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_712
timestamp 25201
transform 1 0 17480 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_713
timestamp 25201
transform 1 0 22632 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_714
timestamp 25201
transform 1 0 27784 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_715
timestamp 25201
transform 1 0 32936 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_716
timestamp 25201
transform 1 0 38088 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_717
timestamp 25201
transform 1 0 43240 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_718
timestamp 25201
transform 1 0 48392 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_719
timestamp 25201
transform 1 0 53544 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_720
timestamp 25201
transform 1 0 58696 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_721
timestamp 25201
transform 1 0 63848 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_722
timestamp 25201
transform 1 0 69000 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_723
timestamp 25201
transform 1 0 74152 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_724
timestamp 25201
transform 1 0 4600 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_725
timestamp 25201
transform 1 0 9752 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_726
timestamp 25201
transform 1 0 14904 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_727
timestamp 25201
transform 1 0 20056 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_728
timestamp 25201
transform 1 0 25208 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_729
timestamp 25201
transform 1 0 30360 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_730
timestamp 25201
transform 1 0 35512 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_731
timestamp 25201
transform 1 0 40664 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_732
timestamp 25201
transform 1 0 45816 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_733
timestamp 25201
transform 1 0 50968 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_734
timestamp 25201
transform 1 0 56120 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_735
timestamp 25201
transform 1 0 61272 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_736
timestamp 25201
transform 1 0 66424 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_737
timestamp 25201
transform 1 0 71576 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_738
timestamp 25201
transform 1 0 76728 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_739
timestamp 25201
transform 1 0 7176 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_740
timestamp 25201
transform 1 0 12328 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_741
timestamp 25201
transform 1 0 17480 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_742
timestamp 25201
transform 1 0 22632 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_743
timestamp 25201
transform 1 0 27784 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_744
timestamp 25201
transform 1 0 32936 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_745
timestamp 25201
transform 1 0 38088 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_746
timestamp 25201
transform 1 0 43240 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_747
timestamp 25201
transform 1 0 48392 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_748
timestamp 25201
transform 1 0 53544 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_749
timestamp 25201
transform 1 0 58696 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_750
timestamp 25201
transform 1 0 63848 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_751
timestamp 25201
transform 1 0 69000 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_752
timestamp 25201
transform 1 0 74152 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_753
timestamp 25201
transform 1 0 4600 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_754
timestamp 25201
transform 1 0 9752 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_755
timestamp 25201
transform 1 0 14904 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_756
timestamp 25201
transform 1 0 20056 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_757
timestamp 25201
transform 1 0 25208 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_758
timestamp 25201
transform 1 0 30360 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_759
timestamp 25201
transform 1 0 35512 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_760
timestamp 25201
transform 1 0 40664 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_761
timestamp 25201
transform 1 0 45816 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_762
timestamp 25201
transform 1 0 50968 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_763
timestamp 25201
transform 1 0 56120 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_764
timestamp 25201
transform 1 0 61272 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_765
timestamp 25201
transform 1 0 66424 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_766
timestamp 25201
transform 1 0 71576 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_767
timestamp 25201
transform 1 0 76728 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_768
timestamp 25201
transform 1 0 7176 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_769
timestamp 25201
transform 1 0 12328 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_770
timestamp 25201
transform 1 0 17480 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_771
timestamp 25201
transform 1 0 22632 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_772
timestamp 25201
transform 1 0 27784 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_773
timestamp 25201
transform 1 0 32936 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_774
timestamp 25201
transform 1 0 38088 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_775
timestamp 25201
transform 1 0 43240 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_776
timestamp 25201
transform 1 0 48392 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_777
timestamp 25201
transform 1 0 53544 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_778
timestamp 25201
transform 1 0 58696 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_779
timestamp 25201
transform 1 0 63848 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_780
timestamp 25201
transform 1 0 69000 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_781
timestamp 25201
transform 1 0 74152 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_782
timestamp 25201
transform 1 0 4600 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_783
timestamp 25201
transform 1 0 9752 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_784
timestamp 25201
transform 1 0 14904 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_785
timestamp 25201
transform 1 0 20056 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_786
timestamp 25201
transform 1 0 25208 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_787
timestamp 25201
transform 1 0 30360 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_788
timestamp 25201
transform 1 0 35512 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_789
timestamp 25201
transform 1 0 40664 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_790
timestamp 25201
transform 1 0 45816 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_791
timestamp 25201
transform 1 0 50968 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_792
timestamp 25201
transform 1 0 56120 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_793
timestamp 25201
transform 1 0 61272 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_794
timestamp 25201
transform 1 0 66424 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_795
timestamp 25201
transform 1 0 71576 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_796
timestamp 25201
transform 1 0 76728 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_797
timestamp 25201
transform 1 0 7176 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_798
timestamp 25201
transform 1 0 12328 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_799
timestamp 25201
transform 1 0 17480 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_800
timestamp 25201
transform 1 0 22632 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_801
timestamp 25201
transform 1 0 27784 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_802
timestamp 25201
transform 1 0 32936 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_803
timestamp 25201
transform 1 0 38088 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_804
timestamp 25201
transform 1 0 43240 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_805
timestamp 25201
transform 1 0 48392 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_806
timestamp 25201
transform 1 0 53544 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_807
timestamp 25201
transform 1 0 58696 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_808
timestamp 25201
transform 1 0 63848 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_809
timestamp 25201
transform 1 0 69000 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_810
timestamp 25201
transform 1 0 74152 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_811
timestamp 25201
transform 1 0 4600 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_812
timestamp 25201
transform 1 0 9752 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_813
timestamp 25201
transform 1 0 14904 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_814
timestamp 25201
transform 1 0 20056 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_815
timestamp 25201
transform 1 0 25208 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_816
timestamp 25201
transform 1 0 30360 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_817
timestamp 25201
transform 1 0 35512 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_818
timestamp 25201
transform 1 0 40664 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_819
timestamp 25201
transform 1 0 45816 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_820
timestamp 25201
transform 1 0 50968 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_821
timestamp 25201
transform 1 0 56120 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_822
timestamp 25201
transform 1 0 61272 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_823
timestamp 25201
transform 1 0 66424 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_824
timestamp 25201
transform 1 0 71576 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_825
timestamp 25201
transform 1 0 76728 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_826
timestamp 25201
transform 1 0 7176 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_827
timestamp 25201
transform 1 0 12328 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_828
timestamp 25201
transform 1 0 17480 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_829
timestamp 25201
transform 1 0 22632 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_830
timestamp 25201
transform 1 0 27784 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_831
timestamp 25201
transform 1 0 32936 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_832
timestamp 25201
transform 1 0 38088 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_833
timestamp 25201
transform 1 0 43240 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_834
timestamp 25201
transform 1 0 48392 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_835
timestamp 25201
transform 1 0 53544 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_836
timestamp 25201
transform 1 0 58696 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_837
timestamp 25201
transform 1 0 63848 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_838
timestamp 25201
transform 1 0 69000 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_839
timestamp 25201
transform 1 0 74152 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_840
timestamp 25201
transform 1 0 4600 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_841
timestamp 25201
transform 1 0 9752 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_842
timestamp 25201
transform 1 0 14904 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_843
timestamp 25201
transform 1 0 20056 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_844
timestamp 25201
transform 1 0 25208 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_845
timestamp 25201
transform 1 0 30360 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_846
timestamp 25201
transform 1 0 35512 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_847
timestamp 25201
transform 1 0 40664 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_848
timestamp 25201
transform 1 0 45816 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_849
timestamp 25201
transform 1 0 50968 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_850
timestamp 25201
transform 1 0 56120 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_851
timestamp 25201
transform 1 0 61272 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_852
timestamp 25201
transform 1 0 66424 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_853
timestamp 25201
transform 1 0 71576 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_854
timestamp 25201
transform 1 0 76728 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_855
timestamp 25201
transform 1 0 7176 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_856
timestamp 25201
transform 1 0 12328 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_857
timestamp 25201
transform 1 0 17480 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_858
timestamp 25201
transform 1 0 22632 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_859
timestamp 25201
transform 1 0 27784 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_860
timestamp 25201
transform 1 0 32936 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_861
timestamp 25201
transform 1 0 38088 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_862
timestamp 25201
transform 1 0 43240 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_863
timestamp 25201
transform 1 0 48392 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_864
timestamp 25201
transform 1 0 53544 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_865
timestamp 25201
transform 1 0 58696 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_866
timestamp 25201
transform 1 0 63848 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_867
timestamp 25201
transform 1 0 69000 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_868
timestamp 25201
transform 1 0 74152 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_869
timestamp 25201
transform 1 0 4600 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_870
timestamp 25201
transform 1 0 9752 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_871
timestamp 25201
transform 1 0 14904 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_872
timestamp 25201
transform 1 0 20056 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_873
timestamp 25201
transform 1 0 25208 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_874
timestamp 25201
transform 1 0 30360 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_875
timestamp 25201
transform 1 0 35512 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_876
timestamp 25201
transform 1 0 40664 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_877
timestamp 25201
transform 1 0 45816 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_878
timestamp 25201
transform 1 0 50968 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_879
timestamp 25201
transform 1 0 56120 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_880
timestamp 25201
transform 1 0 61272 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_881
timestamp 25201
transform 1 0 66424 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_882
timestamp 25201
transform 1 0 71576 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_883
timestamp 25201
transform 1 0 76728 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_884
timestamp 25201
transform 1 0 7176 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_885
timestamp 25201
transform 1 0 12328 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_886
timestamp 25201
transform 1 0 17480 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_887
timestamp 25201
transform 1 0 22632 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_888
timestamp 25201
transform 1 0 27784 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_889
timestamp 25201
transform 1 0 32936 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_890
timestamp 25201
transform 1 0 38088 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_891
timestamp 25201
transform 1 0 43240 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_892
timestamp 25201
transform 1 0 48392 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_893
timestamp 25201
transform 1 0 53544 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_894
timestamp 25201
transform 1 0 58696 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_895
timestamp 25201
transform 1 0 63848 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_896
timestamp 25201
transform 1 0 69000 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_897
timestamp 25201
transform 1 0 74152 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_898
timestamp 25201
transform 1 0 4600 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_899
timestamp 25201
transform 1 0 9752 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_900
timestamp 25201
transform 1 0 14904 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_901
timestamp 25201
transform 1 0 20056 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_902
timestamp 25201
transform 1 0 25208 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_903
timestamp 25201
transform 1 0 30360 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_904
timestamp 25201
transform 1 0 35512 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_905
timestamp 25201
transform 1 0 40664 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_906
timestamp 25201
transform 1 0 45816 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_907
timestamp 25201
transform 1 0 50968 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_908
timestamp 25201
transform 1 0 56120 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_909
timestamp 25201
transform 1 0 61272 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_910
timestamp 25201
transform 1 0 66424 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_911
timestamp 25201
transform 1 0 71576 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_912
timestamp 25201
transform 1 0 76728 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_913
timestamp 25201
transform 1 0 7176 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_914
timestamp 25201
transform 1 0 12328 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_915
timestamp 25201
transform 1 0 17480 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_916
timestamp 25201
transform 1 0 22632 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_917
timestamp 25201
transform 1 0 27784 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_918
timestamp 25201
transform 1 0 32936 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_919
timestamp 25201
transform 1 0 38088 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_920
timestamp 25201
transform 1 0 43240 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_921
timestamp 25201
transform 1 0 48392 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_922
timestamp 25201
transform 1 0 53544 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_923
timestamp 25201
transform 1 0 58696 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_924
timestamp 25201
transform 1 0 63848 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_925
timestamp 25201
transform 1 0 69000 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_926
timestamp 25201
transform 1 0 74152 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_927
timestamp 25201
transform 1 0 4600 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_928
timestamp 25201
transform 1 0 9752 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_929
timestamp 25201
transform 1 0 14904 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_930
timestamp 25201
transform 1 0 20056 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_931
timestamp 25201
transform 1 0 25208 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_932
timestamp 25201
transform 1 0 30360 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_933
timestamp 25201
transform 1 0 35512 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_934
timestamp 25201
transform 1 0 40664 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_935
timestamp 25201
transform 1 0 45816 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_936
timestamp 25201
transform 1 0 50968 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_937
timestamp 25201
transform 1 0 56120 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_938
timestamp 25201
transform 1 0 61272 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_939
timestamp 25201
transform 1 0 66424 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_940
timestamp 25201
transform 1 0 71576 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_941
timestamp 25201
transform 1 0 76728 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_942
timestamp 25201
transform 1 0 7176 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_943
timestamp 25201
transform 1 0 12328 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_944
timestamp 25201
transform 1 0 17480 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_945
timestamp 25201
transform 1 0 22632 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_946
timestamp 25201
transform 1 0 27784 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_947
timestamp 25201
transform 1 0 32936 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_948
timestamp 25201
transform 1 0 38088 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_949
timestamp 25201
transform 1 0 43240 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_950
timestamp 25201
transform 1 0 48392 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_951
timestamp 25201
transform 1 0 53544 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_952
timestamp 25201
transform 1 0 58696 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_953
timestamp 25201
transform 1 0 63848 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_954
timestamp 25201
transform 1 0 69000 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_955
timestamp 25201
transform 1 0 74152 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_956
timestamp 25201
transform 1 0 4600 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_957
timestamp 25201
transform 1 0 9752 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_958
timestamp 25201
transform 1 0 14904 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_959
timestamp 25201
transform 1 0 20056 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_960
timestamp 25201
transform 1 0 25208 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_961
timestamp 25201
transform 1 0 30360 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_962
timestamp 25201
transform 1 0 35512 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_963
timestamp 25201
transform 1 0 40664 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_964
timestamp 25201
transform 1 0 45816 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_965
timestamp 25201
transform 1 0 50968 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_966
timestamp 25201
transform 1 0 56120 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_967
timestamp 25201
transform 1 0 61272 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_968
timestamp 25201
transform 1 0 66424 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_969
timestamp 25201
transform 1 0 71576 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_970
timestamp 25201
transform 1 0 76728 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_971
timestamp 25201
transform 1 0 7176 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_972
timestamp 25201
transform 1 0 12328 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_973
timestamp 25201
transform 1 0 17480 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_974
timestamp 25201
transform 1 0 22632 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_975
timestamp 25201
transform 1 0 27784 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_976
timestamp 25201
transform 1 0 32936 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_977
timestamp 25201
transform 1 0 38088 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_978
timestamp 25201
transform 1 0 43240 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_979
timestamp 25201
transform 1 0 48392 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_980
timestamp 25201
transform 1 0 53544 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_981
timestamp 25201
transform 1 0 58696 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_982
timestamp 25201
transform 1 0 63848 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_983
timestamp 25201
transform 1 0 69000 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_984
timestamp 25201
transform 1 0 74152 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_985
timestamp 25201
transform 1 0 4600 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_986
timestamp 25201
transform 1 0 9752 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_987
timestamp 25201
transform 1 0 14904 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_988
timestamp 25201
transform 1 0 20056 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_989
timestamp 25201
transform 1 0 25208 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_990
timestamp 25201
transform 1 0 30360 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_991
timestamp 25201
transform 1 0 35512 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_992
timestamp 25201
transform 1 0 40664 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_993
timestamp 25201
transform 1 0 45816 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_994
timestamp 25201
transform 1 0 50968 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_995
timestamp 25201
transform 1 0 56120 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_996
timestamp 25201
transform 1 0 61272 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_997
timestamp 25201
transform 1 0 66424 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_998
timestamp 25201
transform 1 0 71576 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_999
timestamp 25201
transform 1 0 76728 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1000
timestamp 25201
transform 1 0 7176 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1001
timestamp 25201
transform 1 0 12328 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1002
timestamp 25201
transform 1 0 17480 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1003
timestamp 25201
transform 1 0 22632 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1004
timestamp 25201
transform 1 0 27784 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1005
timestamp 25201
transform 1 0 32936 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1006
timestamp 25201
transform 1 0 38088 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1007
timestamp 25201
transform 1 0 43240 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1008
timestamp 25201
transform 1 0 48392 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1009
timestamp 25201
transform 1 0 53544 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1010
timestamp 25201
transform 1 0 58696 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1011
timestamp 25201
transform 1 0 63848 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1012
timestamp 25201
transform 1 0 69000 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1013
timestamp 25201
transform 1 0 74152 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1014
timestamp 25201
transform 1 0 4600 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1015
timestamp 25201
transform 1 0 9752 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1016
timestamp 25201
transform 1 0 14904 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1017
timestamp 25201
transform 1 0 20056 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1018
timestamp 25201
transform 1 0 25208 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1019
timestamp 25201
transform 1 0 30360 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1020
timestamp 25201
transform 1 0 35512 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1021
timestamp 25201
transform 1 0 40664 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1022
timestamp 25201
transform 1 0 45816 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1023
timestamp 25201
transform 1 0 50968 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1024
timestamp 25201
transform 1 0 56120 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1025
timestamp 25201
transform 1 0 61272 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1026
timestamp 25201
transform 1 0 66424 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1027
timestamp 25201
transform 1 0 71576 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1028
timestamp 25201
transform 1 0 76728 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1029
timestamp 25201
transform 1 0 7176 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1030
timestamp 25201
transform 1 0 12328 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1031
timestamp 25201
transform 1 0 17480 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1032
timestamp 25201
transform 1 0 22632 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1033
timestamp 25201
transform 1 0 27784 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1034
timestamp 25201
transform 1 0 32936 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1035
timestamp 25201
transform 1 0 38088 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1036
timestamp 25201
transform 1 0 43240 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1037
timestamp 25201
transform 1 0 48392 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1038
timestamp 25201
transform 1 0 53544 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1039
timestamp 25201
transform 1 0 58696 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1040
timestamp 25201
transform 1 0 63848 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1041
timestamp 25201
transform 1 0 69000 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1042
timestamp 25201
transform 1 0 74152 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1043
timestamp 25201
transform 1 0 4600 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1044
timestamp 25201
transform 1 0 9752 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1045
timestamp 25201
transform 1 0 14904 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1046
timestamp 25201
transform 1 0 20056 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1047
timestamp 25201
transform 1 0 25208 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1048
timestamp 25201
transform 1 0 30360 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1049
timestamp 25201
transform 1 0 35512 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1050
timestamp 25201
transform 1 0 40664 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1051
timestamp 25201
transform 1 0 45816 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1052
timestamp 25201
transform 1 0 50968 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1053
timestamp 25201
transform 1 0 56120 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1054
timestamp 25201
transform 1 0 61272 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1055
timestamp 25201
transform 1 0 66424 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1056
timestamp 25201
transform 1 0 71576 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1057
timestamp 25201
transform 1 0 76728 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1058
timestamp 25201
transform 1 0 7176 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1059
timestamp 25201
transform 1 0 12328 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1060
timestamp 25201
transform 1 0 17480 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1061
timestamp 25201
transform 1 0 22632 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1062
timestamp 25201
transform 1 0 27784 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1063
timestamp 25201
transform 1 0 32936 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1064
timestamp 25201
transform 1 0 38088 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1065
timestamp 25201
transform 1 0 43240 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1066
timestamp 25201
transform 1 0 48392 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1067
timestamp 25201
transform 1 0 53544 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1068
timestamp 25201
transform 1 0 58696 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1069
timestamp 25201
transform 1 0 63848 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1070
timestamp 25201
transform 1 0 69000 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1071
timestamp 25201
transform 1 0 74152 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1072
timestamp 25201
transform 1 0 4600 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1073
timestamp 25201
transform 1 0 7176 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1074
timestamp 25201
transform 1 0 9752 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1075
timestamp 25201
transform 1 0 12328 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1076
timestamp 25201
transform 1 0 14904 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1077
timestamp 25201
transform 1 0 17480 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1078
timestamp 25201
transform 1 0 20056 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1079
timestamp 25201
transform 1 0 22632 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1080
timestamp 25201
transform 1 0 25208 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1081
timestamp 25201
transform 1 0 27784 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1082
timestamp 25201
transform 1 0 30360 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1083
timestamp 25201
transform 1 0 32936 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1084
timestamp 25201
transform 1 0 35512 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1085
timestamp 25201
transform 1 0 38088 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1086
timestamp 25201
transform 1 0 40664 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1087
timestamp 25201
transform 1 0 43240 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1088
timestamp 25201
transform 1 0 45816 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1089
timestamp 25201
transform 1 0 48392 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1090
timestamp 25201
transform 1 0 50968 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1091
timestamp 25201
transform 1 0 53544 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1092
timestamp 25201
transform 1 0 56120 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1093
timestamp 25201
transform 1 0 58696 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1094
timestamp 25201
transform 1 0 61272 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1095
timestamp 25201
transform 1 0 63848 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1096
timestamp 25201
transform 1 0 66424 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1097
timestamp 25201
transform 1 0 69000 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1098
timestamp 25201
transform 1 0 71576 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1099
timestamp 25201
transform 1 0 74152 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1100
timestamp 25201
transform 1 0 76728 0 1 36992
box -38 -48 130 592
<< labels >>
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 HADDR[0]
port 0 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 HADDR[10]
port 1 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 HADDR[11]
port 2 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 HADDR[12]
port 3 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 HADDR[13]
port 4 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 HADDR[14]
port 5 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 HADDR[15]
port 6 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 HADDR[16]
port 7 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 HADDR[17]
port 8 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 HADDR[18]
port 9 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 HADDR[19]
port 10 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 HADDR[1]
port 11 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 HADDR[20]
port 12 nsew signal input
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 HADDR[21]
port 13 nsew signal input
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 HADDR[22]
port 14 nsew signal input
flabel metal2 s 60554 0 60610 800 0 FreeSans 224 90 0 0 HADDR[23]
port 15 nsew signal input
flabel metal2 s 62486 0 62542 800 0 FreeSans 224 90 0 0 HADDR[24]
port 16 nsew signal input
flabel metal2 s 64418 0 64474 800 0 FreeSans 224 90 0 0 HADDR[25]
port 17 nsew signal input
flabel metal2 s 66350 0 66406 800 0 FreeSans 224 90 0 0 HADDR[26]
port 18 nsew signal input
flabel metal2 s 68282 0 68338 800 0 FreeSans 224 90 0 0 HADDR[27]
port 19 nsew signal input
flabel metal2 s 70214 0 70270 800 0 FreeSans 224 90 0 0 HADDR[28]
port 20 nsew signal input
flabel metal2 s 72146 0 72202 800 0 FreeSans 224 90 0 0 HADDR[29]
port 21 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 HADDR[2]
port 22 nsew signal input
flabel metal2 s 74078 0 74134 800 0 FreeSans 224 90 0 0 HADDR[30]
port 23 nsew signal input
flabel metal2 s 76010 0 76066 800 0 FreeSans 224 90 0 0 HADDR[31]
port 24 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 HADDR[3]
port 25 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 HADDR[4]
port 26 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 HADDR[5]
port 27 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 HADDR[6]
port 28 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 HADDR[7]
port 29 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 HADDR[8]
port 30 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 HADDR[9]
port 31 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 HCLK
port 32 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 HRDATA[0]
port 33 nsew signal output
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 HRDATA[10]
port 34 nsew signal output
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 HRDATA[11]
port 35 nsew signal output
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 HRDATA[12]
port 36 nsew signal output
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 HRDATA[13]
port 37 nsew signal output
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 HRDATA[14]
port 38 nsew signal output
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 HRDATA[15]
port 39 nsew signal output
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 HRDATA[16]
port 40 nsew signal output
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 HRDATA[17]
port 41 nsew signal output
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 HRDATA[18]
port 42 nsew signal output
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 HRDATA[19]
port 43 nsew signal output
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 HRDATA[1]
port 44 nsew signal output
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 HRDATA[20]
port 45 nsew signal output
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 HRDATA[21]
port 46 nsew signal output
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 HRDATA[22]
port 47 nsew signal output
flabel metal2 s 61198 0 61254 800 0 FreeSans 224 90 0 0 HRDATA[23]
port 48 nsew signal output
flabel metal2 s 63130 0 63186 800 0 FreeSans 224 90 0 0 HRDATA[24]
port 49 nsew signal output
flabel metal2 s 65062 0 65118 800 0 FreeSans 224 90 0 0 HRDATA[25]
port 50 nsew signal output
flabel metal2 s 66994 0 67050 800 0 FreeSans 224 90 0 0 HRDATA[26]
port 51 nsew signal output
flabel metal2 s 68926 0 68982 800 0 FreeSans 224 90 0 0 HRDATA[27]
port 52 nsew signal output
flabel metal2 s 70858 0 70914 800 0 FreeSans 224 90 0 0 HRDATA[28]
port 53 nsew signal output
flabel metal2 s 72790 0 72846 800 0 FreeSans 224 90 0 0 HRDATA[29]
port 54 nsew signal output
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 HRDATA[2]
port 55 nsew signal output
flabel metal2 s 74722 0 74778 800 0 FreeSans 224 90 0 0 HRDATA[30]
port 56 nsew signal output
flabel metal2 s 76654 0 76710 800 0 FreeSans 224 90 0 0 HRDATA[31]
port 57 nsew signal output
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 HRDATA[3]
port 58 nsew signal output
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 HRDATA[4]
port 59 nsew signal output
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 HRDATA[5]
port 60 nsew signal output
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 HRDATA[6]
port 61 nsew signal output
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 HRDATA[7]
port 62 nsew signal output
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 HRDATA[8]
port 63 nsew signal output
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 HRDATA[9]
port 64 nsew signal output
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 HREADY
port 65 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 HREADYOUT
port 66 nsew signal output
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 HRESETn
port 67 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 HSEL
port 68 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 HSIZE[0]
port 69 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 HSIZE[1]
port 70 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 HSIZE[2]
port 71 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 HTRANS[0]
port 72 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 HTRANS[1]
port 73 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 HWDATA[0]
port 74 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 HWDATA[10]
port 75 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 HWDATA[11]
port 76 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 HWDATA[12]
port 77 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 HWDATA[13]
port 78 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 HWDATA[14]
port 79 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 HWDATA[15]
port 80 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 HWDATA[16]
port 81 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 HWDATA[17]
port 82 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 HWDATA[18]
port 83 nsew signal input
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 HWDATA[19]
port 84 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 HWDATA[1]
port 85 nsew signal input
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 HWDATA[20]
port 86 nsew signal input
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 HWDATA[21]
port 87 nsew signal input
flabel metal2 s 59910 0 59966 800 0 FreeSans 224 90 0 0 HWDATA[22]
port 88 nsew signal input
flabel metal2 s 61842 0 61898 800 0 FreeSans 224 90 0 0 HWDATA[23]
port 89 nsew signal input
flabel metal2 s 63774 0 63830 800 0 FreeSans 224 90 0 0 HWDATA[24]
port 90 nsew signal input
flabel metal2 s 65706 0 65762 800 0 FreeSans 224 90 0 0 HWDATA[25]
port 91 nsew signal input
flabel metal2 s 67638 0 67694 800 0 FreeSans 224 90 0 0 HWDATA[26]
port 92 nsew signal input
flabel metal2 s 69570 0 69626 800 0 FreeSans 224 90 0 0 HWDATA[27]
port 93 nsew signal input
flabel metal2 s 71502 0 71558 800 0 FreeSans 224 90 0 0 HWDATA[28]
port 94 nsew signal input
flabel metal2 s 73434 0 73490 800 0 FreeSans 224 90 0 0 HWDATA[29]
port 95 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 HWDATA[2]
port 96 nsew signal input
flabel metal2 s 75366 0 75422 800 0 FreeSans 224 90 0 0 HWDATA[30]
port 97 nsew signal input
flabel metal2 s 77298 0 77354 800 0 FreeSans 224 90 0 0 HWDATA[31]
port 98 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 HWDATA[3]
port 99 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 HWDATA[4]
port 100 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 HWDATA[5]
port 101 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 HWDATA[6]
port 102 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 HWDATA[7]
port 103 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 HWDATA[8]
port 104 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 HWDATA[9]
port 105 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 HWRITE
port 106 nsew signal input
flabel metal2 s 59266 39200 59322 40000 0 FreeSans 224 90 0 0 gpio_oeb[0]
port 107 nsew signal output
flabel metal2 s 22466 39200 22522 40000 0 FreeSans 224 90 0 0 gpio_oeb[10]
port 108 nsew signal output
flabel metal2 s 18786 39200 18842 40000 0 FreeSans 224 90 0 0 gpio_oeb[11]
port 109 nsew signal output
flabel metal2 s 15106 39200 15162 40000 0 FreeSans 224 90 0 0 gpio_oeb[12]
port 110 nsew signal output
flabel metal2 s 11426 39200 11482 40000 0 FreeSans 224 90 0 0 gpio_oeb[13]
port 111 nsew signal output
flabel metal2 s 7746 39200 7802 40000 0 FreeSans 224 90 0 0 gpio_oeb[14]
port 112 nsew signal output
flabel metal2 s 4066 39200 4122 40000 0 FreeSans 224 90 0 0 gpio_oeb[15]
port 113 nsew signal output
flabel metal2 s 55586 39200 55642 40000 0 FreeSans 224 90 0 0 gpio_oeb[1]
port 114 nsew signal output
flabel metal2 s 51906 39200 51962 40000 0 FreeSans 224 90 0 0 gpio_oeb[2]
port 115 nsew signal output
flabel metal2 s 48226 39200 48282 40000 0 FreeSans 224 90 0 0 gpio_oeb[3]
port 116 nsew signal output
flabel metal2 s 44546 39200 44602 40000 0 FreeSans 224 90 0 0 gpio_oeb[4]
port 117 nsew signal output
flabel metal2 s 40866 39200 40922 40000 0 FreeSans 224 90 0 0 gpio_oeb[5]
port 118 nsew signal output
flabel metal2 s 37186 39200 37242 40000 0 FreeSans 224 90 0 0 gpio_oeb[6]
port 119 nsew signal output
flabel metal2 s 33506 39200 33562 40000 0 FreeSans 224 90 0 0 gpio_oeb[7]
port 120 nsew signal output
flabel metal2 s 29826 39200 29882 40000 0 FreeSans 224 90 0 0 gpio_oeb[8]
port 121 nsew signal output
flabel metal2 s 26146 39200 26202 40000 0 FreeSans 224 90 0 0 gpio_oeb[9]
port 122 nsew signal output
flabel metal2 s 57426 39200 57482 40000 0 FreeSans 224 90 0 0 gpio_out[0]
port 123 nsew signal output
flabel metal2 s 20626 39200 20682 40000 0 FreeSans 224 90 0 0 gpio_out[10]
port 124 nsew signal output
flabel metal2 s 16946 39200 17002 40000 0 FreeSans 224 90 0 0 gpio_out[11]
port 125 nsew signal output
flabel metal2 s 13266 39200 13322 40000 0 FreeSans 224 90 0 0 gpio_out[12]
port 126 nsew signal output
flabel metal2 s 9586 39200 9642 40000 0 FreeSans 224 90 0 0 gpio_out[13]
port 127 nsew signal output
flabel metal2 s 5906 39200 5962 40000 0 FreeSans 224 90 0 0 gpio_out[14]
port 128 nsew signal output
flabel metal2 s 2226 39200 2282 40000 0 FreeSans 224 90 0 0 gpio_out[15]
port 129 nsew signal output
flabel metal2 s 53746 39200 53802 40000 0 FreeSans 224 90 0 0 gpio_out[1]
port 130 nsew signal output
flabel metal2 s 50066 39200 50122 40000 0 FreeSans 224 90 0 0 gpio_out[2]
port 131 nsew signal output
flabel metal2 s 46386 39200 46442 40000 0 FreeSans 224 90 0 0 gpio_out[3]
port 132 nsew signal output
flabel metal2 s 42706 39200 42762 40000 0 FreeSans 224 90 0 0 gpio_out[4]
port 133 nsew signal output
flabel metal2 s 39026 39200 39082 40000 0 FreeSans 224 90 0 0 gpio_out[5]
port 134 nsew signal output
flabel metal2 s 35346 39200 35402 40000 0 FreeSans 224 90 0 0 gpio_out[6]
port 135 nsew signal output
flabel metal2 s 31666 39200 31722 40000 0 FreeSans 224 90 0 0 gpio_out[7]
port 136 nsew signal output
flabel metal2 s 27986 39200 28042 40000 0 FreeSans 224 90 0 0 gpio_out[8]
port 137 nsew signal output
flabel metal2 s 24306 39200 24362 40000 0 FreeSans 224 90 0 0 gpio_out[9]
port 138 nsew signal output
flabel metal4 s 5128 2128 5448 37584 0 FreeSans 1920 90 0 0 vccd1
port 139 nsew power bidirectional
flabel metal4 s 35848 2128 36168 37584 0 FreeSans 1920 90 0 0 vccd1
port 139 nsew power bidirectional
flabel metal4 s 66568 2128 66888 37584 0 FreeSans 1920 90 0 0 vccd1
port 139 nsew power bidirectional
flabel metal4 s 5788 2128 6108 37584 0 FreeSans 1920 90 0 0 vssd1
port 140 nsew ground bidirectional
flabel metal4 s 36508 2128 36828 37584 0 FreeSans 1920 90 0 0 vssd1
port 140 nsew ground bidirectional
flabel metal4 s 67228 2128 67548 37584 0 FreeSans 1920 90 0 0 vssd1
port 140 nsew ground bidirectional
rlabel metal1 39974 37536 39974 37536 0 vccd1
rlabel metal1 39974 36992 39974 36992 0 vssd1
rlabel metal2 18814 7514 18814 7514 0 CTRL_REG
rlabel metal1 10350 5032 10350 5032 0 HADDR[0]
rlabel metal2 35466 1761 35466 1761 0 HADDR[10]
rlabel metal2 37444 7820 37444 7820 0 HADDR[11]
rlabel metal2 39330 4580 39330 4580 0 HADDR[12]
rlabel metal2 41262 959 41262 959 0 HADDR[13]
rlabel metal1 43470 5678 43470 5678 0 HADDR[14]
rlabel metal1 46046 3094 46046 3094 0 HADDR[15]
rlabel metal2 16146 1044 16146 1044 0 HADDR[1]
rlabel metal2 19366 1027 19366 1027 0 HADDR[2]
rlabel metal1 21620 9486 21620 9486 0 HADDR[3]
rlabel metal2 18630 1958 18630 1958 0 HADDR[4]
rlabel via2 16330 5763 16330 5763 0 HADDR[5]
rlabel metal3 27623 5508 27623 5508 0 HADDR[6]
rlabel metal2 29670 1761 29670 1761 0 HADDR[7]
rlabel metal2 21758 1533 21758 1533 0 HADDR[8]
rlabel metal2 33534 1761 33534 1761 0 HADDR[9]
rlabel metal2 9154 493 9154 493 0 HCLK
rlabel metal2 13570 1554 13570 1554 0 HRDATA[0]
rlabel metal2 36110 1095 36110 1095 0 HRDATA[10]
rlabel metal2 38042 1095 38042 1095 0 HRDATA[11]
rlabel metal2 39974 959 39974 959 0 HRDATA[12]
rlabel metal2 41906 1622 41906 1622 0 HRDATA[13]
rlabel metal2 43838 1554 43838 1554 0 HRDATA[14]
rlabel metal1 46276 3570 46276 3570 0 HRDATA[15]
rlabel metal1 48254 2958 48254 2958 0 HRDATA[16]
rlabel metal2 51566 1860 51566 1860 0 HRDATA[18]
rlabel metal2 53498 1860 53498 1860 0 HRDATA[19]
rlabel metal1 17756 3706 17756 3706 0 HRDATA[1]
rlabel metal2 57362 1554 57362 1554 0 HRDATA[21]
rlabel metal2 61226 1860 61226 1860 0 HRDATA[23]
rlabel metal2 65090 1860 65090 1860 0 HRDATA[25]
rlabel metal2 67022 1826 67022 1826 0 HRDATA[26]
rlabel metal2 68954 1860 68954 1860 0 HRDATA[27]
rlabel metal2 70886 1860 70886 1860 0 HRDATA[28]
rlabel metal2 20010 1095 20010 1095 0 HRDATA[2]
rlabel metal2 74750 1860 74750 1860 0 HRDATA[30]
rlabel metal2 76682 1435 76682 1435 0 HRDATA[31]
rlabel metal2 22586 1095 22586 1095 0 HRDATA[3]
rlabel metal1 24196 3366 24196 3366 0 HRDATA[4]
rlabel metal2 26450 1622 26450 1622 0 HRDATA[5]
rlabel metal1 28888 3570 28888 3570 0 HRDATA[6]
rlabel metal2 30314 1622 30314 1622 0 HRDATA[7]
rlabel metal2 32246 1622 32246 1622 0 HRDATA[8]
rlabel metal2 34178 1554 34178 1554 0 HRDATA[9]
rlabel metal2 9706 1554 9706 1554 0 HREADY
rlabel metal1 5474 3604 5474 3604 0 HRESETn
rlabel metal2 6302 2822 6302 2822 0 HSEL
rlabel metal1 8786 4012 8786 4012 0 HTRANS[1]
rlabel metal2 7682 3349 7682 3349 0 HWDATA[0]
rlabel metal2 36754 823 36754 823 0 HWDATA[10]
rlabel metal2 38686 2115 38686 2115 0 HWDATA[11]
rlabel metal2 40618 942 40618 942 0 HWDATA[12]
rlabel metal2 42550 1044 42550 1044 0 HWDATA[13]
rlabel metal2 44482 1384 44482 1384 0 HWDATA[14]
rlabel metal2 46414 823 46414 823 0 HWDATA[15]
rlabel metal2 7682 1360 7682 1360 0 HWDATA[1]
rlabel metal1 10120 3366 10120 3366 0 HWDATA[2]
rlabel metal2 8418 1292 8418 1292 0 HWDATA[3]
rlabel metal1 24886 10030 24886 10030 0 HWDATA[4]
rlabel metal1 20010 6222 20010 6222 0 HWDATA[5]
rlabel metal2 29026 9741 29026 9741 0 HWDATA[6]
rlabel metal2 30958 3475 30958 3475 0 HWDATA[7]
rlabel metal2 32798 561 32798 561 0 HWDATA[8]
rlabel metal2 34822 823 34822 823 0 HWDATA[9]
rlabel metal2 12282 3492 12282 3492 0 HWRITE
rlabel metal2 8602 2856 8602 2856 0 _000_
rlabel metal1 20700 5338 20700 5338 0 _001_
rlabel metal1 20509 6970 20509 6970 0 _002_
rlabel metal1 21528 8058 21528 8058 0 _003_
rlabel metal1 24242 6732 24242 6732 0 _004_
rlabel metal2 14306 3655 14306 3655 0 _005_
rlabel metal2 23506 7004 23506 7004 0 _006_
rlabel metal1 26496 6426 26496 6426 0 _007_
rlabel metal2 25898 7072 25898 7072 0 _008_
rlabel metal1 28520 7378 28520 7378 0 _009_
rlabel metal1 27186 2890 27186 2890 0 _010_
rlabel metal2 32246 7956 32246 7956 0 _011_
rlabel metal1 35834 9010 35834 9010 0 _012_
rlabel metal1 36938 8534 36938 8534 0 _013_
rlabel metal1 34914 5236 34914 5236 0 _014_
rlabel metal1 34960 4998 34960 4998 0 _015_
rlabel metal2 31142 6817 31142 6817 0 _016_
rlabel metal1 36478 6426 36478 6426 0 _017_
rlabel metal1 7682 4556 7682 4556 0 _018_
rlabel metal1 10166 2584 10166 2584 0 _019_
rlabel metal2 10626 6562 10626 6562 0 _020_
rlabel metal1 17388 2618 17388 2618 0 _021_
rlabel via2 8418 3043 8418 3043 0 _022_
rlabel via2 10258 3485 10258 3485 0 _023_
rlabel metal1 21298 5848 21298 5848 0 _024_
rlabel metal2 10626 2176 10626 2176 0 _025_
rlabel via2 22034 7293 22034 7293 0 _026_
rlabel metal1 29716 3978 29716 3978 0 _027_
rlabel metal1 31372 4794 31372 4794 0 _028_
rlabel via2 33074 2907 33074 2907 0 _029_
rlabel metal1 34776 3706 34776 3706 0 _030_
rlabel metal1 36892 3910 36892 3910 0 _031_
rlabel metal1 40388 3366 40388 3366 0 _032_
rlabel metal2 41722 3298 41722 3298 0 _033_
rlabel metal1 44804 2618 44804 2618 0 _034_
rlabel metal1 45908 3706 45908 3706 0 _035_
rlabel metal4 21804 7004 21804 7004 0 _036_
rlabel metal1 32430 6358 32430 6358 0 _037_
rlabel metal2 33166 6052 33166 6052 0 _038_
rlabel metal1 37582 5814 37582 5814 0 _039_
rlabel metal1 39698 2380 39698 2380 0 _040_
rlabel metal2 38962 2210 38962 2210 0 _041_
rlabel metal2 38870 7004 38870 7004 0 _042_
rlabel metal1 27830 12614 27830 12614 0 _043_
rlabel metal1 36662 2278 36662 2278 0 _044_
rlabel metal2 10626 4454 10626 4454 0 _045_
rlabel metal1 12604 4114 12604 4114 0 _046_
rlabel metal1 19274 9520 19274 9520 0 _047_
rlabel metal1 19182 6936 19182 6936 0 _048_
rlabel metal2 18630 5049 18630 5049 0 _049_
rlabel metal1 21390 5202 21390 5202 0 _050_
rlabel metal2 24242 10234 24242 10234 0 _051_
rlabel metal2 33718 7497 33718 7497 0 _052_
rlabel metal2 16698 4352 16698 4352 0 _053_
rlabel metal1 35834 6630 35834 6630 0 _054_
rlabel metal1 21068 6222 21068 6222 0 _055_
rlabel metal2 21758 5508 21758 5508 0 _056_
rlabel metal2 20930 8517 20930 8517 0 _057_
rlabel metal2 21390 7293 21390 7293 0 _058_
rlabel metal1 20654 7820 20654 7820 0 _059_
rlabel metal1 20470 7922 20470 7922 0 _060_
rlabel metal1 20470 5542 20470 5542 0 _061_
rlabel metal1 20792 3910 20792 3910 0 _062_
rlabel metal1 20976 5882 20976 5882 0 _063_
rlabel metal1 25300 9894 25300 9894 0 _064_
rlabel metal2 24794 11424 24794 11424 0 _065_
rlabel via2 26726 3995 26726 3995 0 _066_
rlabel metal1 24978 5338 24978 5338 0 _067_
rlabel metal1 24610 7990 24610 7990 0 _068_
rlabel metal1 24288 7310 24288 7310 0 _069_
rlabel metal1 28106 8432 28106 8432 0 _070_
rlabel metal2 22586 4250 22586 4250 0 _071_
rlabel metal1 27646 6426 27646 6426 0 _072_
rlabel metal1 28198 7990 28198 7990 0 _073_
rlabel metal1 22540 2278 22540 2278 0 _074_
rlabel metal2 28474 7820 28474 7820 0 _075_
rlabel metal1 28198 2992 28198 2992 0 _076_
rlabel metal1 33212 10574 33212 10574 0 _077_
rlabel metal2 28014 3196 28014 3196 0 _078_
rlabel metal1 30360 5542 30360 5542 0 _079_
rlabel metal1 26082 5678 26082 5678 0 _080_
rlabel metal1 32255 7310 32255 7310 0 _081_
rlabel metal2 32522 8908 32522 8908 0 _082_
rlabel metal1 35098 10744 35098 10744 0 _083_
rlabel metal1 33626 8534 33626 8534 0 _084_
rlabel metal1 35282 8058 35282 8058 0 _085_
rlabel metal1 28290 3060 28290 3060 0 _086_
rlabel metal1 39330 3536 39330 3536 0 _087_
rlabel metal1 35006 5882 35006 5882 0 _088_
rlabel metal1 40710 3604 40710 3604 0 _089_
rlabel metal1 34270 5236 34270 5236 0 _090_
rlabel metal1 31096 7854 31096 7854 0 _091_
rlabel metal1 36156 4250 36156 4250 0 _092_
rlabel metal1 30452 8058 30452 8058 0 _093_
rlabel metal2 30866 10030 30866 10030 0 _094_
rlabel metal2 34270 4386 34270 4386 0 _095_
rlabel metal1 35696 6290 35696 6290 0 _096_
rlabel metal2 40618 6528 40618 6528 0 _097_
rlabel metal2 36202 6511 36202 6511 0 _098_
rlabel metal1 22724 5270 22724 5270 0 clknet_0_HCLK
rlabel metal1 12006 3468 12006 3468 0 clknet_2_0__leaf_HCLK
rlabel metal2 18078 7854 18078 7854 0 clknet_2_1__leaf_HCLK
rlabel metal1 38686 3094 38686 3094 0 clknet_2_2__leaf_HCLK
rlabel metal2 34178 8126 34178 8126 0 clknet_2_3__leaf_HCLK
rlabel metal1 59846 36754 59846 36754 0 gpio_oeb[0]
rlabel metal1 23138 37162 23138 37162 0 gpio_oeb[10]
rlabel metal1 19182 37230 19182 37230 0 gpio_oeb[11]
rlabel metal1 15594 37162 15594 37162 0 gpio_oeb[12]
rlabel metal1 11408 37230 11408 37230 0 gpio_oeb[13]
rlabel metal1 8372 37230 8372 37230 0 gpio_oeb[14]
rlabel metal1 4232 36822 4232 36822 0 gpio_oeb[15]
rlabel metal1 56442 37162 56442 37162 0 gpio_oeb[1]
rlabel metal1 52532 37230 52532 37230 0 gpio_oeb[2]
rlabel metal1 48806 37162 48806 37162 0 gpio_oeb[3]
rlabel metal1 44942 36686 44942 36686 0 gpio_oeb[4]
rlabel metal1 41492 37230 41492 37230 0 gpio_oeb[5]
rlabel metal1 37398 37230 37398 37230 0 gpio_oeb[6]
rlabel metal1 33810 37298 33810 37298 0 gpio_oeb[7]
rlabel metal1 30406 36754 30406 36754 0 gpio_oeb[8]
rlabel metal2 26174 38192 26174 38192 0 gpio_oeb[9]
rlabel metal1 58604 37162 58604 37162 0 gpio_out[0]
rlabel metal1 20792 37230 20792 37230 0 gpio_out[10]
rlabel metal1 17480 36822 17480 36822 0 gpio_out[11]
rlabel metal1 13432 37298 13432 37298 0 gpio_out[12]
rlabel metal1 9752 36822 9752 36822 0 gpio_out[13]
rlabel metal2 5934 38226 5934 38226 0 gpio_out[14]
rlabel metal1 2392 37298 2392 37298 0 gpio_out[15]
rlabel metal1 54280 37162 54280 37162 0 gpio_out[1]
rlabel metal1 50370 36686 50370 36686 0 gpio_out[2]
rlabel metal1 46920 37162 46920 37162 0 gpio_out[3]
rlabel metal1 43516 37162 43516 37162 0 gpio_out[4]
rlabel metal1 39330 37298 39330 37298 0 gpio_out[5]
rlabel metal2 35374 37954 35374 37954 0 gpio_out[6]
rlabel metal1 31740 37230 31740 37230 0 gpio_out[7]
rlabel metal1 28152 37230 28152 37230 0 gpio_out[8]
rlabel metal1 24472 36822 24472 36822 0 gpio_out[9]
rlabel metal1 15364 3502 15364 3502 0 last_HADDR\[0\]
rlabel metal2 35098 4539 35098 4539 0 last_HADDR\[10\]
rlabel metal2 36202 4454 36202 4454 0 last_HADDR\[11\]
rlabel metal1 40802 3162 40802 3162 0 last_HADDR\[12\]
rlabel metal1 40618 4250 40618 4250 0 last_HADDR\[13\]
rlabel metal1 45034 2414 45034 2414 0 last_HADDR\[14\]
rlabel metal1 44988 3502 44988 3502 0 last_HADDR\[15\]
rlabel metal2 9154 2210 9154 2210 0 last_HADDR\[1\]
rlabel metal1 17756 7310 17756 7310 0 last_HADDR\[2\]
rlabel metal1 21206 4182 21206 4182 0 last_HADDR\[3\]
rlabel metal1 26772 10030 26772 10030 0 last_HADDR\[4\]
rlabel metal1 27232 3162 27232 3162 0 last_HADDR\[5\]
rlabel metal2 19366 5967 19366 5967 0 last_HADDR\[6\]
rlabel metal1 17250 4726 17250 4726 0 last_HADDR\[7\]
rlabel metal1 31694 4522 31694 4522 0 last_HADDR\[8\]
rlabel metal1 33396 3162 33396 3162 0 last_HADDR\[9\]
rlabel metal1 11914 2958 11914 2958 0 last_HSEL
rlabel metal1 12167 5678 12167 5678 0 last_HTRANS\[1\]
rlabel metal1 13294 3570 13294 3570 0 last_HWRITE
rlabel metal2 7958 4284 7958 4284 0 net1
rlabel metal1 16008 6222 16008 6222 0 net10
rlabel metal2 17618 4590 17618 4590 0 net100
rlabel metal1 39790 4624 39790 4624 0 net101
rlabel metal2 16330 2315 16330 2315 0 net102
rlabel metal1 19228 9690 19228 9690 0 net103
rlabel metal1 24012 9350 24012 9350 0 net104
rlabel metal2 34316 7718 34316 7718 0 net105
rlabel metal2 28750 4454 28750 4454 0 net106
rlabel metal1 19274 36720 19274 36720 0 net107
rlabel metal1 44390 36652 44390 36652 0 net108
rlabel metal1 23651 7786 23651 7786 0 net109
rlabel metal2 13202 5185 13202 5185 0 net11
rlabel metal1 25859 4182 25859 4182 0 net110
rlabel metal2 28106 10064 28106 10064 0 net111
rlabel metal2 13018 8398 13018 8398 0 net112
rlabel metal2 10166 6035 10166 6035 0 net113
rlabel metal2 10074 3570 10074 3570 0 net114
rlabel metal1 44850 2482 44850 2482 0 net115
rlabel metal2 49634 1656 49634 1656 0 net116
rlabel metal2 55430 1588 55430 1588 0 net117
rlabel metal2 59294 1792 59294 1792 0 net118
rlabel metal2 63158 1588 63158 1588 0 net119
rlabel metal2 11914 3876 11914 3876 0 net12
rlabel metal2 72818 1622 72818 1622 0 net120
rlabel metal2 10350 2183 10350 2183 0 net121
rlabel metal1 13478 4794 13478 4794 0 net122
rlabel metal2 26174 6732 26174 6732 0 net123
rlabel metal2 13018 2210 13018 2210 0 net124
rlabel metal2 32430 9452 32430 9452 0 net125
rlabel metal2 33534 3791 33534 3791 0 net126
rlabel metal2 32430 4199 32430 4199 0 net127
rlabel metal1 10120 2890 10120 2890 0 net128
rlabel metal2 19182 4182 19182 4182 0 net129
rlabel metal2 12190 5151 12190 5151 0 net13
rlabel metal1 11454 3638 11454 3638 0 net130
rlabel metal1 36110 9554 36110 9554 0 net131
rlabel metal1 36156 3366 36156 3366 0 net132
rlabel metal2 35650 5406 35650 5406 0 net133
rlabel metal2 47426 2176 47426 2176 0 net134
rlabel metal1 41147 2958 41147 2958 0 net135
rlabel metal2 41722 4794 41722 4794 0 net136
rlabel metal2 22034 9758 22034 9758 0 net137
rlabel metal1 23552 4454 23552 4454 0 net138
rlabel metal2 21482 3264 21482 3264 0 net139
rlabel metal2 24426 6324 24426 6324 0 net14
rlabel metal1 21068 12682 21068 12682 0 net140
rlabel metal2 28382 7004 28382 7004 0 net141
rlabel metal1 27002 3400 27002 3400 0 net142
rlabel via2 5842 2499 5842 2499 0 net143
rlabel metal1 19412 4046 19412 4046 0 net144
rlabel metal2 11454 3162 11454 3162 0 net145
rlabel metal1 26588 2278 26588 2278 0 net146
rlabel metal2 36110 4318 36110 4318 0 net147
rlabel metal2 37674 5712 37674 5712 0 net148
rlabel metal2 37214 9333 37214 9333 0 net149
rlabel metal1 24518 6188 24518 6188 0 net15
rlabel metal1 21666 5576 21666 5576 0 net150
rlabel metal2 30038 6494 30038 6494 0 net151
rlabel metal1 45540 5134 45540 5134 0 net152
rlabel metal2 45862 2516 45862 2516 0 net153
rlabel metal1 41952 2958 41952 2958 0 net154
rlabel metal2 8970 5508 8970 5508 0 net155
rlabel metal2 8326 2414 8326 2414 0 net156
rlabel metal1 17618 3570 17618 3570 0 net157
rlabel metal2 46966 5372 46966 5372 0 net158
rlabel metal1 44988 3570 44988 3570 0 net159
rlabel metal2 20378 1938 20378 1938 0 net16
rlabel metal1 43240 3570 43240 3570 0 net160
rlabel metal1 13984 2414 13984 2414 0 net161
rlabel metal2 31878 4828 31878 4828 0 net162
rlabel metal2 31234 3298 31234 3298 0 net163
rlabel metal2 41446 7854 41446 7854 0 net164
rlabel metal2 41262 2550 41262 2550 0 net165
rlabel metal1 38686 2958 38686 2958 0 net166
rlabel metal2 7590 4386 7590 4386 0 net167
rlabel metal1 10396 3706 10396 3706 0 net168
rlabel metal1 8694 3162 8694 3162 0 net169
rlabel metal1 5290 2618 5290 2618 0 net17
rlabel metal2 4370 4930 4370 4930 0 net170
rlabel metal2 15502 5134 15502 5134 0 net171
rlabel metal2 11638 6596 11638 6596 0 net172
rlabel metal2 11178 6902 11178 6902 0 net173
rlabel metal1 14444 5746 14444 5746 0 net174
rlabel metal1 12098 3944 12098 3944 0 net175
rlabel metal2 25990 9996 25990 9996 0 net176
rlabel metal1 19366 5882 19366 5882 0 net177
rlabel metal1 24334 6970 24334 6970 0 net178
rlabel metal1 15732 4046 15732 4046 0 net179
rlabel metal1 5336 3026 5336 3026 0 net18
rlabel metal1 23368 6834 23368 6834 0 net180
rlabel metal1 26818 6698 26818 6698 0 net181
rlabel metal1 19734 8058 19734 8058 0 net182
rlabel metal1 10810 4148 10810 4148 0 net183
rlabel metal1 23782 4012 23782 4012 0 net184
rlabel metal1 34960 2482 34960 2482 0 net185
rlabel metal1 36064 5134 36064 5134 0 net186
rlabel metal1 38032 4794 38032 4794 0 net187
rlabel metal1 22862 2618 22862 2618 0 net188
rlabel metal2 31878 6562 31878 6562 0 net189
rlabel metal2 5750 2788 5750 2788 0 net19
rlabel metal2 33902 8007 33902 8007 0 net190
rlabel metal3 35903 7956 35903 7956 0 net191
rlabel metal1 31878 6290 31878 6290 0 net192
rlabel metal2 35098 8670 35098 8670 0 net193
rlabel metal2 28658 9265 28658 9265 0 net194
rlabel metal1 29164 8398 29164 8398 0 net195
rlabel metal1 30130 8058 30130 8058 0 net196
rlabel metal1 9476 4658 9476 4658 0 net197
rlabel metal1 11960 4794 11960 4794 0 net198
rlabel metal1 24702 6834 24702 6834 0 net199
rlabel metal1 25622 2516 25622 2516 0 net2
rlabel metal1 13708 5678 13708 5678 0 net20
rlabel metal2 4002 5406 4002 5406 0 net200
rlabel metal2 18722 5882 18722 5882 0 net201
rlabel metal1 18906 5270 18906 5270 0 net202
rlabel metal1 5658 2414 5658 2414 0 net203
rlabel metal2 21758 8670 21758 8670 0 net204
rlabel metal2 22402 8024 22402 8024 0 net205
rlabel metal2 48070 3876 48070 3876 0 net206
rlabel metal1 34546 5202 34546 5202 0 net207
rlabel metal1 37214 5882 37214 5882 0 net208
rlabel metal2 32890 9826 32890 9826 0 net209
rlabel metal1 15134 7276 15134 7276 0 net21
rlabel metal1 32062 9010 32062 9010 0 net210
rlabel metal2 27278 4284 27278 4284 0 net211
rlabel metal1 29992 5270 29992 5270 0 net212
rlabel metal1 47748 4658 47748 4658 0 net213
rlabel metal2 38962 3774 38962 3774 0 net214
rlabel metal1 29486 5202 29486 5202 0 net215
rlabel metal1 33304 6358 33304 6358 0 net216
rlabel metal2 19274 5525 19274 5525 0 net217
rlabel metal2 27002 5712 27002 5712 0 net218
rlabel metal1 29716 7514 29716 7514 0 net219
rlabel metal2 20654 2176 20654 2176 0 net22
rlabel metal1 29762 7310 29762 7310 0 net220
rlabel metal2 8234 5984 8234 5984 0 net221
rlabel metal2 4554 4760 4554 4760 0 net222
rlabel metal2 14582 6732 14582 6732 0 net223
rlabel metal1 21436 6426 21436 6426 0 net224
rlabel metal2 50094 3604 50094 3604 0 net225
rlabel metal1 43424 4658 43424 4658 0 net226
rlabel metal1 36110 6324 36110 6324 0 net227
rlabel metal1 37490 6698 37490 6698 0 net228
rlabel metal1 11730 5338 11730 5338 0 net229
rlabel metal1 39146 4012 39146 4012 0 net23
rlabel metal2 14858 5916 14858 5916 0 net230
rlabel metal1 14674 4012 14674 4012 0 net231
rlabel metal1 38962 5780 38962 5780 0 net232
rlabel metal2 33994 4794 33994 4794 0 net233
rlabel metal1 36156 6970 36156 6970 0 net234
rlabel metal1 37680 8058 37680 8058 0 net235
rlabel metal1 14720 6426 14720 6426 0 net236
rlabel metal2 11178 4284 11178 4284 0 net237
rlabel metal1 18722 7242 18722 7242 0 net238
rlabel metal2 30314 4080 30314 4080 0 net239
rlabel metal1 38456 3162 38456 3162 0 net24
rlabel metal1 45540 2958 45540 2958 0 net240
rlabel metal1 19734 5542 19734 5542 0 net241
rlabel metal1 44344 2958 44344 2958 0 net242
rlabel metal1 31855 10098 31855 10098 0 net243
rlabel metal1 32476 4046 32476 4046 0 net244
rlabel metal2 28198 5814 28198 5814 0 net245
rlabel metal1 22494 2482 22494 2482 0 net246
rlabel metal1 30314 2414 30314 2414 0 net247
rlabel metal2 28290 6460 28290 6460 0 net248
rlabel metal1 19320 4658 19320 4658 0 net249
rlabel metal2 45402 3672 45402 3672 0 net25
rlabel metal2 29118 3774 29118 3774 0 net250
rlabel metal1 36892 4658 36892 4658 0 net251
rlabel metal2 32798 3740 32798 3740 0 net252
rlabel metal2 38686 3842 38686 3842 0 net253
rlabel metal1 35512 5678 35512 5678 0 net254
rlabel metal2 37950 7293 37950 7293 0 net255
rlabel metal2 36846 3842 36846 3842 0 net256
rlabel metal1 23000 5746 23000 5746 0 net257
rlabel metal1 18584 5882 18584 5882 0 net258
rlabel metal1 25162 2482 25162 2482 0 net259
rlabel metal1 46414 2550 46414 2550 0 net26
rlabel metal1 29946 6290 29946 6290 0 net260
rlabel metal2 25530 5916 25530 5916 0 net261
rlabel metal2 35282 3196 35282 3196 0 net262
rlabel metal2 16330 4794 16330 4794 0 net263
rlabel metal2 13478 6953 13478 6953 0 net264
rlabel metal2 22862 3842 22862 3842 0 net265
rlabel metal2 40526 5372 40526 5372 0 net266
rlabel metal1 41814 2448 41814 2448 0 net267
rlabel metal1 43194 2414 43194 2414 0 net268
rlabel metal2 22954 3757 22954 3757 0 net269
rlabel metal1 46828 2890 46828 2890 0 net27
rlabel metal2 13294 4726 13294 4726 0 net270
rlabel metal3 18653 2516 18653 2516 0 net271
rlabel metal1 41952 5338 41952 5338 0 net272
rlabel metal1 38548 3502 38548 3502 0 net273
rlabel metal1 37950 2380 37950 2380 0 net274
rlabel metal1 20148 7310 20148 7310 0 net275
rlabel metal1 16054 2448 16054 2448 0 net276
rlabel metal1 20378 2380 20378 2380 0 net277
rlabel metal2 39974 4828 39974 4828 0 net278
rlabel metal2 46138 3468 46138 3468 0 net279
rlabel metal1 19826 9452 19826 9452 0 net28
rlabel metal2 46506 3230 46506 3230 0 net280
rlabel metal1 16284 6290 16284 6290 0 net281
rlabel metal2 17802 7922 17802 7922 0 net282
rlabel metal2 18262 3774 18262 3774 0 net283
rlabel metal1 17756 4726 17756 4726 0 net284
rlabel metal1 43470 3026 43470 3026 0 net285
rlabel metal1 42642 2618 42642 2618 0 net287
rlabel metal2 77050 3808 77050 3808 0 net289
rlabel metal1 12328 5202 12328 5202 0 net29
rlabel metal2 28014 4709 28014 4709 0 net290
rlabel metal1 22310 9010 22310 9010 0 net291
rlabel metal2 15962 7242 15962 7242 0 net292
rlabel metal1 77326 2924 77326 2924 0 net295
rlabel metal1 76590 2482 76590 2482 0 net296
rlabel metal2 6026 3910 6026 3910 0 net297
rlabel metal2 8050 4250 8050 4250 0 net298
rlabel metal1 9982 5168 9982 5168 0 net299
rlabel metal1 38180 9010 38180 9010 0 net3
rlabel metal1 16790 5202 16790 5202 0 net30
rlabel metal1 27232 4046 27232 4046 0 net300
rlabel metal2 17250 5372 17250 5372 0 net302
rlabel via2 52670 4165 52670 4165 0 net305
rlabel metal2 58098 3332 58098 3332 0 net306
rlabel metal1 58512 2482 58512 2482 0 net307
rlabel metal1 5290 3400 5290 3400 0 net31
rlabel metal1 57178 3060 57178 3060 0 net312
rlabel metal2 65458 3604 65458 3604 0 net313
rlabel metal2 65550 2754 65550 2754 0 net314
rlabel metal2 18446 7616 18446 7616 0 net318
rlabel metal1 27278 9010 27278 9010 0 net32
rlabel metal1 52256 3162 52256 3162 0 net320
rlabel metal2 52118 2754 52118 2754 0 net321
rlabel metal2 56074 3196 56074 3196 0 net327
rlabel metal2 54050 2754 54050 2754 0 net328
rlabel metal2 19458 4709 19458 4709 0 net33
rlabel metal2 67942 3876 67942 3876 0 net334
rlabel metal2 67666 2754 67666 2754 0 net335
rlabel metal2 14122 4301 14122 4301 0 net34
rlabel metal1 61916 3162 61916 3162 0 net341
rlabel metal2 61778 2754 61778 2754 0 net342
rlabel metal2 71530 3196 71530 3196 0 net348
rlabel metal2 69506 2754 69506 2754 0 net349
rlabel metal3 32476 8568 32476 8568 0 net35
rlabel metal2 72450 3740 72450 3740 0 net355
rlabel metal2 72634 2754 72634 2754 0 net356
rlabel metal1 7912 3638 7912 3638 0 net357
rlabel metal2 6762 3230 6762 3230 0 net358
rlabel metal1 27002 3570 27002 3570 0 net359
rlabel metal1 24380 2550 24380 2550 0 net36
rlabel metal1 10672 3094 10672 3094 0 net360
rlabel metal2 40894 6018 40894 6018 0 net366
rlabel metal1 49956 3910 49956 3910 0 net367
rlabel metal1 49634 2482 49634 2482 0 net368
rlabel metal1 10350 6630 10350 6630 0 net37
rlabel metal2 76958 4964 76958 4964 0 net373
rlabel metal2 75486 2958 75486 2958 0 net374
rlabel metal1 29026 7922 29026 7922 0 net376
rlabel metal2 32706 7004 32706 7004 0 net377
rlabel metal1 33396 9894 33396 9894 0 net378
rlabel metal2 35742 6698 35742 6698 0 net379
rlabel metal1 16974 7514 16974 7514 0 net38
rlabel metal1 32614 6120 32614 6120 0 net380
rlabel metal2 28566 10710 28566 10710 0 net381
rlabel via2 11730 4029 11730 4029 0 net383
rlabel metal1 18262 2414 18262 2414 0 net384
rlabel metal1 24932 3502 24932 3502 0 net385
rlabel metal1 14996 5882 14996 5882 0 net386
rlabel metal1 27940 4046 27940 4046 0 net387
rlabel metal2 35282 5032 35282 5032 0 net39
rlabel metal2 74566 3196 74566 3196 0 net390
rlabel metal2 76222 2618 76222 2618 0 net391
rlabel metal2 76682 2822 76682 2822 0 net392
rlabel metal1 11500 6290 11500 6290 0 net393
rlabel metal2 7866 4454 7866 4454 0 net394
rlabel metal1 11454 3468 11454 3468 0 net395
rlabel metal1 12788 2482 12788 2482 0 net396
rlabel metal1 28934 5134 28934 5134 0 net397
rlabel metal1 23736 5814 23736 5814 0 net398
rlabel metal1 21758 5746 21758 5746 0 net399
rlabel metal2 35834 2210 35834 2210 0 net4
rlabel metal1 33994 4692 33994 4692 0 net40
rlabel metal1 23644 2278 23644 2278 0 net400
rlabel metal1 38410 7310 38410 7310 0 net401
rlabel metal1 36248 4794 36248 4794 0 net402
rlabel metal1 31280 4046 31280 4046 0 net403
rlabel metal1 29762 6834 29762 6834 0 net404
rlabel metal1 28888 6426 28888 6426 0 net405
rlabel metal1 21666 4624 21666 4624 0 net406
rlabel metal2 18538 4505 18538 4505 0 net407
rlabel metal1 22448 5746 22448 5746 0 net408
rlabel metal1 26818 8058 26818 8058 0 net409
rlabel metal2 40158 6494 40158 6494 0 net41
rlabel metal1 17802 5678 17802 5678 0 net410
rlabel metal1 25208 4590 25208 4590 0 net411
rlabel metal1 36524 7310 36524 7310 0 net412
rlabel metal1 32614 2890 32614 2890 0 net413
rlabel metal2 31878 5423 31878 5423 0 net414
rlabel metal1 36524 3502 36524 3502 0 net415
rlabel metal1 15824 4590 15824 4590 0 net416
rlabel metal4 13708 5780 13708 5780 0 net417
rlabel metal2 24150 9860 24150 9860 0 net418
rlabel metal1 21206 3502 21206 3502 0 net419
rlabel metal1 41538 4692 41538 4692 0 net42
rlabel metal1 34316 7514 34316 7514 0 net420
rlabel via2 32338 7701 32338 7701 0 net421
rlabel metal1 27554 5338 27554 5338 0 net422
rlabel metal1 32614 4046 32614 4046 0 net423
rlabel metal1 40940 6222 40940 6222 0 net424
rlabel metal1 41860 5202 41860 5202 0 net425
rlabel metal1 40020 2482 40020 2482 0 net426
rlabel metal1 39284 5202 39284 5202 0 net427
rlabel metal1 41584 5882 41584 5882 0 net428
rlabel metal2 34914 4862 34914 4862 0 net429
rlabel metal1 36662 2856 36662 2856 0 net43
rlabel metal1 21114 7412 21114 7412 0 net430
rlabel metal2 22310 9078 22310 9078 0 net431
rlabel metal1 9752 3026 9752 3026 0 net432
rlabel metal1 40020 5678 40020 5678 0 net434
rlabel metal1 40986 4726 40986 4726 0 net435
rlabel metal1 44206 4114 44206 4114 0 net436
rlabel metal2 23414 7956 23414 7956 0 net437
rlabel metal2 16698 8500 16698 8500 0 net438
rlabel metal1 11592 4046 11592 4046 0 net439
rlabel metal1 42504 4046 42504 4046 0 net44
rlabel metal1 13616 4658 13616 4658 0 net441
rlabel metal3 11799 3876 11799 3876 0 net442
rlabel metal1 13570 4114 13570 4114 0 net443
rlabel metal2 34822 10268 34822 10268 0 net444
rlabel metal2 20194 2108 20194 2108 0 net445
rlabel metal1 21390 4590 21390 4590 0 net446
rlabel metal2 9062 6443 9062 6443 0 net447
rlabel via2 15226 5355 15226 5355 0 net448
rlabel metal1 16054 6426 16054 6426 0 net449
rlabel metal1 48484 3978 48484 3978 0 net45
rlabel via2 15318 5627 15318 5627 0 net450
rlabel metal2 22586 10370 22586 10370 0 net451
rlabel metal1 14996 5270 14996 5270 0 net452
rlabel metal2 21574 2057 21574 2057 0 net453
rlabel metal1 28750 8942 28750 8942 0 net454
rlabel metal1 21390 6290 21390 6290 0 net455
rlabel metal1 35006 9146 35006 9146 0 net456
rlabel metal3 34339 8500 34339 8500 0 net457
rlabel metal3 35397 7684 35397 7684 0 net458
rlabel metal1 47518 2482 47518 2482 0 net459
rlabel metal2 51290 3332 51290 3332 0 net46
rlabel metal1 40480 2414 40480 2414 0 net460
rlabel metal1 43102 5746 43102 5746 0 net461
rlabel metal1 26772 9622 26772 9622 0 net462
rlabel via2 17066 4811 17066 4811 0 net463
rlabel metal3 20263 12444 20263 12444 0 net464
rlabel metal3 36225 8364 36225 8364 0 net465
rlabel metal1 28428 5542 28428 5542 0 net466
rlabel via2 37398 8891 37398 8891 0 net467
rlabel metal1 44574 5202 44574 5202 0 net468
rlabel metal2 45862 4012 45862 4012 0 net469
rlabel metal2 53682 3332 53682 3332 0 net47
rlabel metal2 49818 4556 49818 4556 0 net470
rlabel metal1 17342 8058 17342 8058 0 net471
rlabel metal2 6394 3400 6394 3400 0 net472
rlabel metal2 10810 6426 10810 6426 0 net473
rlabel metal1 40112 8398 40112 8398 0 net474
rlabel metal1 38180 1938 38180 1938 0 net475
rlabel metal2 32798 2108 32798 2108 0 net476
rlabel metal1 8418 4692 8418 4692 0 net477
rlabel metal2 3634 4148 3634 4148 0 net478
rlabel metal2 7038 4726 7038 4726 0 net479
rlabel via3 10925 4012 10925 4012 0 net48
rlabel metal2 31878 10081 31878 10081 0 net480
rlabel metal1 17618 3094 17618 3094 0 net481
rlabel metal1 25484 6426 25484 6426 0 net482
rlabel metal1 9844 5338 9844 5338 0 net483
rlabel metal2 4922 3570 4922 3570 0 net484
rlabel metal1 8004 2278 8004 2278 0 net485
rlabel metal1 48852 3706 48852 3706 0 net486
rlabel metal1 46138 3502 46138 3502 0 net487
rlabel metal1 47886 4046 47886 4046 0 net488
rlabel metal1 27508 10234 27508 10234 0 net489
rlabel metal2 57362 3332 57362 3332 0 net49
rlabel metal1 54372 3502 54372 3502 0 net493
rlabel metal2 55338 2618 55338 2618 0 net494
rlabel metal2 27462 4301 27462 4301 0 net495
rlabel metal2 57454 3196 57454 3196 0 net499
rlabel metal1 41492 2550 41492 2550 0 net5
rlabel metal2 60950 3332 60950 3332 0 net50
rlabel metal2 58650 2890 58650 2890 0 net500
rlabel metal1 10258 2482 10258 2482 0 net501
rlabel metal2 51474 3196 51474 3196 0 net505
rlabel metal2 53038 2890 53038 2890 0 net506
rlabel metal2 43838 3570 43838 3570 0 net507
rlabel metal2 64722 3332 64722 3332 0 net51
rlabel metal2 64906 3196 64906 3196 0 net511
rlabel metal2 66286 3162 66286 3162 0 net512
rlabel metal2 19274 9622 19274 9622 0 net515
rlabel metal2 61134 3196 61134 3196 0 net516
rlabel metal2 62790 2890 62790 2890 0 net517
rlabel metal1 30222 4658 30222 4658 0 net518
rlabel metal1 26082 7922 26082 7922 0 net519
rlabel metal1 67160 3162 67160 3162 0 net52
rlabel metal1 69828 3502 69828 3502 0 net521
rlabel metal2 70518 2618 70518 2618 0 net522
rlabel metal1 68172 3502 68172 3502 0 net526
rlabel metal2 68310 3162 68310 3162 0 net527
rlabel metal2 69138 3332 69138 3332 0 net53
rlabel metal2 71714 3876 71714 3876 0 net531
rlabel metal2 73094 2890 73094 2890 0 net532
rlabel metal1 9844 4114 9844 4114 0 net533
rlabel metal1 18676 8058 18676 8058 0 net534
rlabel metal1 14306 5882 14306 5882 0 net535
rlabel metal1 15272 2482 15272 2482 0 net536
rlabel metal2 8970 2006 8970 2006 0 net539
rlabel metal1 71576 2618 71576 2618 0 net54
rlabel metal1 23276 10642 23276 10642 0 net540
rlabel metal1 10350 4046 10350 4046 0 net541
rlabel metal1 22862 5100 22862 5100 0 net542
rlabel metal1 25116 9894 25116 9894 0 net543
rlabel metal3 4991 3604 4991 3604 0 net544
rlabel metal1 15732 4794 15732 4794 0 net545
rlabel metal1 22862 6222 22862 6222 0 net546
rlabel metal1 18124 5746 18124 5746 0 net547
rlabel metal1 17802 10438 17802 10438 0 net548
rlabel metal1 22908 6834 22908 6834 0 net549
rlabel metal2 22678 10268 22678 10268 0 net55
rlabel metal2 27278 7378 27278 7378 0 net550
rlabel metal1 44620 4658 44620 4658 0 net551
rlabel metal1 34316 2618 34316 2618 0 net552
rlabel metal1 39928 7310 39928 7310 0 net553
rlabel metal1 36800 5202 36800 5202 0 net554
rlabel metal1 16008 2618 16008 2618 0 net555
rlabel metal1 28336 9690 28336 9690 0 net556
rlabel via2 20010 4437 20010 4437 0 net557
rlabel metal1 25990 6698 25990 6698 0 net558
rlabel metal1 11040 3978 11040 3978 0 net559
rlabel metal2 74474 3332 74474 3332 0 net56
rlabel metal1 10396 4794 10396 4794 0 net560
rlabel metal1 11500 4658 11500 4658 0 net561
rlabel metal2 21574 8126 21574 8126 0 net562
rlabel metal1 20746 2516 20746 2516 0 net563
rlabel metal1 25760 2346 25760 2346 0 net564
rlabel metal1 28244 4726 28244 4726 0 net565
rlabel metal1 32706 6970 32706 6970 0 net566
rlabel metal2 38778 9724 38778 9724 0 net567
rlabel metal1 20470 2380 20470 2380 0 net568
rlabel metal1 28842 4794 28842 4794 0 net569
rlabel metal1 75302 4080 75302 4080 0 net57
rlabel metal1 34960 6970 34960 6970 0 net570
rlabel metal1 9016 2618 9016 2618 0 net571
rlabel via2 5658 2363 5658 2363 0 net572
rlabel metal1 20516 9486 20516 9486 0 net573
rlabel metal1 21022 7854 21022 7854 0 net574
rlabel metal2 47518 3468 47518 3468 0 net575
rlabel metal1 45632 3026 45632 3026 0 net576
rlabel metal1 45586 4012 45586 4012 0 net577
rlabel metal1 12742 3162 12742 3162 0 net58
rlabel metal2 50554 4284 50554 4284 0 net581
rlabel metal2 32246 9061 32246 9061 0 net582
rlabel metal2 32890 4352 32890 4352 0 net583
rlabel metal2 18722 4845 18722 4845 0 net584
rlabel metal1 12558 2482 12558 2482 0 net585
rlabel metal1 48990 4522 48990 4522 0 net586
rlabel metal1 48576 4454 48576 4454 0 net587
rlabel metal2 34270 5899 34270 5899 0 net588
rlabel via2 28842 2363 28842 2363 0 net589
rlabel metal1 24012 2822 24012 2822 0 net59
rlabel metal2 50646 3196 50646 3196 0 net590
rlabel metal1 48806 3026 48806 3026 0 net591
rlabel metal2 6854 4012 6854 4012 0 net592
rlabel metal2 4738 3978 4738 3978 0 net593
rlabel metal2 13846 5338 13846 5338 0 net595
rlabel metal2 77602 4148 77602 4148 0 net598
rlabel metal2 76682 4250 76682 4250 0 net599
rlabel metal1 45816 3162 45816 3162 0 net6
rlabel metal1 25898 9010 25898 9010 0 net60
rlabel metal2 74658 3366 74658 3366 0 net600
rlabel metal1 34224 6834 34224 6834 0 net601
rlabel metal1 33442 5202 33442 5202 0 net602
rlabel metal2 30498 6494 30498 6494 0 net603
rlabel metal2 33258 4556 33258 4556 0 net604
rlabel metal1 14214 6222 14214 6222 0 net605
rlabel metal1 18400 8398 18400 8398 0 net606
rlabel metal1 39790 6290 39790 6290 0 net607
rlabel metal1 41630 6290 41630 6290 0 net608
rlabel metal1 41262 5746 41262 5746 0 net609
rlabel metal1 29348 9010 29348 9010 0 net61
rlabel metal1 38318 5100 38318 5100 0 net610
rlabel metal1 40756 5134 40756 5134 0 net611
rlabel metal2 39146 6188 39146 6188 0 net612
rlabel metal2 39054 5338 39054 5338 0 net613
rlabel metal2 28842 9180 28842 9180 0 net62
rlabel metal1 32016 3638 32016 3638 0 net63
rlabel metal2 25714 5491 25714 5491 0 net64
rlabel metal1 59018 36618 59018 36618 0 net65
rlabel metal1 21022 9044 21022 9044 0 net652
rlabel metal1 14582 6086 14582 6086 0 net653
rlabel metal2 22494 37060 22494 37060 0 net66
rlabel metal1 18906 36890 18906 36890 0 net67
rlabel metal2 37490 7548 37490 7548 0 net674
rlabel metal2 37306 6698 37306 6698 0 net675
rlabel metal2 15134 37060 15134 37060 0 net68
rlabel metal2 11914 37060 11914 37060 0 net69
rlabel metal1 47380 3366 47380 3366 0 net7
rlabel metal2 7774 37060 7774 37060 0 net70
rlabel metal1 19182 6358 19182 6358 0 net704
rlabel metal1 18584 7378 18584 7378 0 net705
rlabel metal2 11822 36686 11822 36686 0 net71
rlabel metal2 55614 37060 55614 37060 0 net72
rlabel metal2 51934 37060 51934 37060 0 net73
rlabel metal2 48254 37060 48254 37060 0 net74
rlabel metal1 44574 36686 44574 36686 0 net75
rlabel metal1 19320 6766 19320 6766 0 net758
rlabel metal1 14766 5338 14766 5338 0 net759
rlabel metal2 40894 37060 40894 37060 0 net76
rlabel metal2 37030 37060 37030 37060 0 net77
rlabel metal2 33810 37060 33810 37060 0 net78
rlabel metal2 18262 6426 18262 6426 0 net786
rlabel metal1 10672 5202 10672 5202 0 net787
rlabel metal1 14214 6290 14214 6290 0 net788
rlabel metal1 29854 36686 29854 36686 0 net79
rlabel metal2 3818 4386 3818 4386 0 net8
rlabel metal1 26128 36890 26128 36890 0 net80
rlabel metal2 58834 25840 58834 25840 0 net81
rlabel metal1 18584 6290 18584 6290 0 net816
rlabel metal1 14168 5678 14168 5678 0 net817
rlabel metal1 20194 7378 20194 7378 0 net818
rlabel metal2 21942 27625 21942 27625 0 net82
rlabel metal2 18998 33167 18998 33167 0 net83
rlabel metal2 14582 25857 14582 25857 0 net84
rlabel metal2 10902 31807 10902 31807 0 net85
rlabel via3 7061 36516 7061 36516 0 net86
rlabel metal2 3542 30685 3542 30685 0 net87
rlabel metal1 39790 26894 39790 26894 0 net88
rlabel metal1 38134 29614 38134 29614 0 net89
rlabel metal2 10258 6460 10258 6460 0 net9
rlabel metal1 36018 24106 36018 24106 0 net90
rlabel metal2 43378 34816 43378 34816 0 net91
rlabel metal2 39146 25857 39146 25857 0 net92
rlabel metal1 33580 17850 33580 17850 0 net93
rlabel via3 32821 36516 32821 36516 0 net94
rlabel metal1 30222 17850 30222 17850 0 net95
rlabel metal2 25806 34918 25806 34918 0 net96
rlabel metal2 23138 10166 23138 10166 0 net97
rlabel metal1 33718 10642 33718 10642 0 net98
rlabel metal1 26680 11118 26680 11118 0 net99
<< properties >>
string FIXED_BBOX 0 0 80000 40000
<< end >>
