VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2720.000 BY 2300.000 ;
  PIN HADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 258.110 -2.000 258.390 4.000 ;
    END
  END HADDR[0]
  PIN HADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 336.310 -2.000 336.590 4.000 ;
    END
  END HADDR[10]
  PIN HADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 344.130 -2.000 344.410 4.000 ;
    END
  END HADDR[11]
  PIN HADDR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 351.950 -2.000 352.230 4.000 ;
    END
  END HADDR[12]
  PIN HADDR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 359.770 -2.000 360.050 4.000 ;
    END
  END HADDR[13]
  PIN HADDR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 367.590 -2.000 367.870 4.000 ;
    END
  END HADDR[14]
  PIN HADDR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 375.410 -2.000 375.690 4.000 ;
    END
  END HADDR[15]
  PIN HADDR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.230 -2.000 383.510 4.000 ;
    END
  END HADDR[16]
  PIN HADDR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.050 -2.000 391.330 4.000 ;
    END
  END HADDR[17]
  PIN HADDR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.870 -2.000 399.150 4.000 ;
    END
  END HADDR[18]
  PIN HADDR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.690 -2.000 406.970 4.000 ;
    END
  END HADDR[19]
  PIN HADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 265.930 -2.000 266.210 4.000 ;
    END
  END HADDR[1]
  PIN HADDR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.510 -2.000 414.790 4.000 ;
    END
  END HADDR[20]
  PIN HADDR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.330 -2.000 422.610 4.000 ;
    END
  END HADDR[21]
  PIN HADDR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.150 -2.000 430.430 4.000 ;
    END
  END HADDR[22]
  PIN HADDR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.970 -2.000 438.250 4.000 ;
    END
  END HADDR[23]
  PIN HADDR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.790 -2.000 446.070 4.000 ;
    END
  END HADDR[24]
  PIN HADDR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.610 -2.000 453.890 4.000 ;
    END
  END HADDR[25]
  PIN HADDR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.430 -2.000 461.710 4.000 ;
    END
  END HADDR[26]
  PIN HADDR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.250 -2.000 469.530 4.000 ;
    END
  END HADDR[27]
  PIN HADDR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.070 -2.000 477.350 4.000 ;
    END
  END HADDR[28]
  PIN HADDR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.890 -2.000 485.170 4.000 ;
    END
  END HADDR[29]
  PIN HADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 273.750 -2.000 274.030 4.000 ;
    END
  END HADDR[2]
  PIN HADDR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.710 -2.000 492.990 4.000 ;
    END
  END HADDR[30]
  PIN HADDR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.530 -2.000 500.810 4.000 ;
    END
  END HADDR[31]
  PIN HADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 281.570 -2.000 281.850 4.000 ;
    END
  END HADDR[3]
  PIN HADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 289.390 -2.000 289.670 4.000 ;
    END
  END HADDR[4]
  PIN HADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 297.210 -2.000 297.490 4.000 ;
    END
  END HADDR[5]
  PIN HADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 305.030 -2.000 305.310 4.000 ;
    END
  END HADDR[6]
  PIN HADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 312.850 -2.000 313.130 4.000 ;
    END
  END HADDR[7]
  PIN HADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 320.670 -2.000 320.950 4.000 ;
    END
  END HADDR[8]
  PIN HADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 328.490 -2.000 328.770 4.000 ;
    END
  END HADDR[9]
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 234.650 -2.000 234.930 4.000 ;
    END
  END HCLK
  PIN HRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 813.330 -2.000 813.610 4.000 ;
    END
  END HRDATA[0]
  PIN HRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 891.530 -2.000 891.810 4.000 ;
    END
  END HRDATA[10]
  PIN HRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 899.350 -2.000 899.630 4.000 ;
    END
  END HRDATA[11]
  PIN HRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 907.170 -2.000 907.450 4.000 ;
    END
  END HRDATA[12]
  PIN HRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 914.990 -2.000 915.270 4.000 ;
    END
  END HRDATA[13]
  PIN HRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 922.810 -2.000 923.090 4.000 ;
    END
  END HRDATA[14]
  PIN HRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 930.630 -2.000 930.910 4.000 ;
    END
  END HRDATA[15]
  PIN HRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 938.450 -2.000 938.730 4.000 ;
    END
  END HRDATA[16]
  PIN HRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.270 -2.000 946.550 4.000 ;
    END
  END HRDATA[17]
  PIN HRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 954.090 -2.000 954.370 4.000 ;
    END
  END HRDATA[18]
  PIN HRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 961.910 -2.000 962.190 4.000 ;
    END
  END HRDATA[19]
  PIN HRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 821.150 -2.000 821.430 4.000 ;
    END
  END HRDATA[1]
  PIN HRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.730 -2.000 970.010 4.000 ;
    END
  END HRDATA[20]
  PIN HRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 977.550 -2.000 977.830 4.000 ;
    END
  END HRDATA[21]
  PIN HRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.370 -2.000 985.650 4.000 ;
    END
  END HRDATA[22]
  PIN HRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 993.190 -2.000 993.470 4.000 ;
    END
  END HRDATA[23]
  PIN HRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.010 -2.000 1001.290 4.000 ;
    END
  END HRDATA[24]
  PIN HRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1008.830 -2.000 1009.110 4.000 ;
    END
  END HRDATA[25]
  PIN HRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1016.650 -2.000 1016.930 4.000 ;
    END
  END HRDATA[26]
  PIN HRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1024.470 -2.000 1024.750 4.000 ;
    END
  END HRDATA[27]
  PIN HRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1032.290 -2.000 1032.570 4.000 ;
    END
  END HRDATA[28]
  PIN HRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.110 -2.000 1040.390 4.000 ;
    END
  END HRDATA[29]
  PIN HRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 828.970 -2.000 829.250 4.000 ;
    END
  END HRDATA[2]
  PIN HRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1047.930 -2.000 1048.210 4.000 ;
    END
  END HRDATA[30]
  PIN HRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1055.750 -2.000 1056.030 4.000 ;
    END
  END HRDATA[31]
  PIN HRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 836.790 -2.000 837.070 4.000 ;
    END
  END HRDATA[3]
  PIN HRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 844.610 -2.000 844.890 4.000 ;
    END
  END HRDATA[4]
  PIN HRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 852.430 -2.000 852.710 4.000 ;
    END
  END HRDATA[5]
  PIN HRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 860.250 -2.000 860.530 4.000 ;
    END
  END HRDATA[6]
  PIN HRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 868.070 -2.000 868.350 4.000 ;
    END
  END HRDATA[7]
  PIN HRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 875.890 -2.000 876.170 4.000 ;
    END
  END HRDATA[8]
  PIN HRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 883.710 -2.000 883.990 4.000 ;
    END
  END HRDATA[9]
  PIN HREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 758.590 -2.000 758.870 4.000 ;
    END
  END HREADY
  PIN HREADYOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.570 -2.000 1063.850 4.000 ;
    END
  END HREADYOUT
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 242.470 -2.000 242.750 4.000 ;
    END
  END HRESETn
  PIN HSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 250.290 -2.000 250.570 4.000 ;
    END
  END HSEL
  PIN HSIZE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.870 -2.000 790.150 4.000 ;
    END
  END HSIZE[0]
  PIN HSIZE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.690 -2.000 797.970 4.000 ;
    END
  END HSIZE[1]
  PIN HSIZE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.510 -2.000 805.790 4.000 ;
    END
  END HSIZE[2]
  PIN HTRANS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.230 -2.000 774.510 4.000 ;
    END
  END HTRANS[0]
  PIN HTRANS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 782.050 -2.000 782.330 4.000 ;
    END
  END HTRANS[1]
  PIN HWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 508.350 -2.000 508.630 4.000 ;
    END
  END HWDATA[0]
  PIN HWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 586.550 -2.000 586.830 4.000 ;
    END
  END HWDATA[10]
  PIN HWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 594.370 -2.000 594.650 4.000 ;
    END
  END HWDATA[11]
  PIN HWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 602.190 -2.000 602.470 4.000 ;
    END
  END HWDATA[12]
  PIN HWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 610.010 -2.000 610.290 4.000 ;
    END
  END HWDATA[13]
  PIN HWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 617.830 -2.000 618.110 4.000 ;
    END
  END HWDATA[14]
  PIN HWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 625.650 -2.000 625.930 4.000 ;
    END
  END HWDATA[15]
  PIN HWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.470 -2.000 633.750 4.000 ;
    END
  END HWDATA[16]
  PIN HWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.290 -2.000 641.570 4.000 ;
    END
  END HWDATA[17]
  PIN HWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.110 -2.000 649.390 4.000 ;
    END
  END HWDATA[18]
  PIN HWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.930 -2.000 657.210 4.000 ;
    END
  END HWDATA[19]
  PIN HWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 516.170 -2.000 516.450 4.000 ;
    END
  END HWDATA[1]
  PIN HWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.750 -2.000 665.030 4.000 ;
    END
  END HWDATA[20]
  PIN HWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.570 -2.000 672.850 4.000 ;
    END
  END HWDATA[21]
  PIN HWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.390 -2.000 680.670 4.000 ;
    END
  END HWDATA[22]
  PIN HWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.210 -2.000 688.490 4.000 ;
    END
  END HWDATA[23]
  PIN HWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.030 -2.000 696.310 4.000 ;
    END
  END HWDATA[24]
  PIN HWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.850 -2.000 704.130 4.000 ;
    END
  END HWDATA[25]
  PIN HWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.670 -2.000 711.950 4.000 ;
    END
  END HWDATA[26]
  PIN HWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.490 -2.000 719.770 4.000 ;
    END
  END HWDATA[27]
  PIN HWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.310 -2.000 727.590 4.000 ;
    END
  END HWDATA[28]
  PIN HWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.130 -2.000 735.410 4.000 ;
    END
  END HWDATA[29]
  PIN HWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 523.990 -2.000 524.270 4.000 ;
    END
  END HWDATA[2]
  PIN HWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.950 -2.000 743.230 4.000 ;
    END
  END HWDATA[30]
  PIN HWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.770 -2.000 751.050 4.000 ;
    END
  END HWDATA[31]
  PIN HWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 531.810 -2.000 532.090 4.000 ;
    END
  END HWDATA[3]
  PIN HWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 539.630 -2.000 539.910 4.000 ;
    END
  END HWDATA[4]
  PIN HWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 547.450 -2.000 547.730 4.000 ;
    END
  END HWDATA[5]
  PIN HWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 555.270 -2.000 555.550 4.000 ;
    END
  END HWDATA[6]
  PIN HWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 563.090 -2.000 563.370 4.000 ;
    END
  END HWDATA[7]
  PIN HWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 570.910 -2.000 571.190 4.000 ;
    END
  END HWDATA[8]
  PIN HWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 578.730 -2.000 579.010 4.000 ;
    END
  END HWDATA[9]
  PIN HWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 766.410 -2.000 766.690 4.000 ;
    END
  END HWRITE
  PIN adc0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1698.125 2298.500 1698.765 2300.000 ;
    END
  END adc0
  PIN adc1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1700.685 2298.500 1701.325 2300.000 ;
    END
  END adc1
  PIN comp_n
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1703.245 2298.500 1703.885 2300.000 ;
    END
  END comp_n
  PIN comp_p
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1705.805 2298.500 1706.445 2300.000 ;
    END
  END comp_p
  PIN dac0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1682.765 2298.500 1683.405 2300.000 ;
    END
  END dac0
  PIN dac1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1685.325 2298.500 1685.965 2300.000 ;
    END
  END dac1
  PIN gpio0_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 97.090 2722.000 97.690 ;
    END
  END gpio0_in[0]
  PIN gpio0_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 166.450 2722.000 167.050 ;
    END
  END gpio0_in[1]
  PIN gpio0_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 235.810 2722.000 236.410 ;
    END
  END gpio0_in[2]
  PIN gpio0_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 305.170 2722.000 305.770 ;
    END
  END gpio0_in[3]
  PIN gpio0_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 374.530 2722.000 375.130 ;
    END
  END gpio0_in[4]
  PIN gpio0_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 443.890 2722.000 444.490 ;
    END
  END gpio0_in[5]
  PIN gpio0_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 513.250 2722.000 513.850 ;
    END
  END gpio0_in[6]
  PIN gpio0_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 582.610 2722.000 583.210 ;
    END
  END gpio0_in[7]
  PIN gpio0_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 143.330 2722.000 143.930 ;
    END
  END gpio0_oeb[0]
  PIN gpio0_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 212.690 2722.000 213.290 ;
    END
  END gpio0_oeb[1]
  PIN gpio0_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 282.050 2722.000 282.650 ;
    END
  END gpio0_oeb[2]
  PIN gpio0_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 351.410 2722.000 352.010 ;
    END
  END gpio0_oeb[3]
  PIN gpio0_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 420.770 2722.000 421.370 ;
    END
  END gpio0_oeb[4]
  PIN gpio0_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 490.130 2722.000 490.730 ;
    END
  END gpio0_oeb[5]
  PIN gpio0_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 559.490 2722.000 560.090 ;
    END
  END gpio0_oeb[6]
  PIN gpio0_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 628.850 2722.000 629.450 ;
    END
  END gpio0_oeb[7]
  PIN gpio0_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 120.210 2722.000 120.810 ;
    END
  END gpio0_out[0]
  PIN gpio0_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 189.570 2722.000 190.170 ;
    END
  END gpio0_out[1]
  PIN gpio0_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 258.930 2722.000 259.530 ;
    END
  END gpio0_out[2]
  PIN gpio0_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 328.290 2722.000 328.890 ;
    END
  END gpio0_out[3]
  PIN gpio0_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 397.650 2722.000 398.250 ;
    END
  END gpio0_out[4]
  PIN gpio0_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 467.010 2722.000 467.610 ;
    END
  END gpio0_out[5]
  PIN gpio0_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 536.370 2722.000 536.970 ;
    END
  END gpio0_out[6]
  PIN gpio0_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 605.730 2722.000 606.330 ;
    END
  END gpio0_out[7]
  PIN gpio1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 894.920 2722.000 895.520 ;
    END
  END gpio1_in[0]
  PIN gpio1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 964.280 2722.000 964.880 ;
    END
  END gpio1_in[1]
  PIN gpio1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1033.640 2722.000 1034.240 ;
    END
  END gpio1_in[2]
  PIN gpio1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1103.000 2722.000 1103.600 ;
    END
  END gpio1_in[3]
  PIN gpio1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1172.360 2722.000 1172.960 ;
    END
  END gpio1_in[4]
  PIN gpio1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1241.720 2722.000 1242.320 ;
    END
  END gpio1_in[5]
  PIN gpio1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1311.080 2722.000 1311.680 ;
    END
  END gpio1_in[6]
  PIN gpio1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1380.440 2722.000 1381.040 ;
    END
  END gpio1_in[7]
  PIN gpio1_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 941.160 2722.000 941.760 ;
    END
  END gpio1_oeb[0]
  PIN gpio1_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1010.520 2722.000 1011.120 ;
    END
  END gpio1_oeb[1]
  PIN gpio1_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1079.880 2722.000 1080.480 ;
    END
  END gpio1_oeb[2]
  PIN gpio1_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1149.240 2722.000 1149.840 ;
    END
  END gpio1_oeb[3]
  PIN gpio1_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1218.600 2722.000 1219.200 ;
    END
  END gpio1_oeb[4]
  PIN gpio1_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1287.960 2722.000 1288.560 ;
    END
  END gpio1_oeb[5]
  PIN gpio1_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1357.320 2722.000 1357.920 ;
    END
  END gpio1_oeb[6]
  PIN gpio1_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1426.680 2722.000 1427.280 ;
    END
  END gpio1_oeb[7]
  PIN gpio1_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 918.040 2722.000 918.640 ;
    END
  END gpio1_out[0]
  PIN gpio1_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 987.400 2722.000 988.000 ;
    END
  END gpio1_out[1]
  PIN gpio1_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1056.760 2722.000 1057.360 ;
    END
  END gpio1_out[2]
  PIN gpio1_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1126.120 2722.000 1126.720 ;
    END
  END gpio1_out[3]
  PIN gpio1_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1195.480 2722.000 1196.080 ;
    END
  END gpio1_out[4]
  PIN gpio1_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1264.840 2722.000 1265.440 ;
    END
  END gpio1_out[5]
  PIN gpio1_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1334.200 2722.000 1334.800 ;
    END
  END gpio1_out[6]
  PIN gpio1_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1403.560 2722.000 1404.160 ;
    END
  END gpio1_out[7]
  PIN gpio2_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1449.800 2722.000 1450.400 ;
    END
  END gpio2_in[0]
  PIN gpio2_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1519.160 2722.000 1519.760 ;
    END
  END gpio2_in[1]
  PIN gpio2_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1588.520 2722.000 1589.120 ;
    END
  END gpio2_in[2]
  PIN gpio2_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1657.880 2722.000 1658.480 ;
    END
  END gpio2_in[3]
  PIN gpio2_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2027.800 2722.000 2028.400 ;
    END
  END gpio2_in[4]
  PIN gpio2_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2097.160 2722.000 2097.760 ;
    END
  END gpio2_in[5]
  PIN gpio2_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2166.520 2722.000 2167.120 ;
    END
  END gpio2_in[6]
  PIN gpio2_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2235.880 2722.000 2236.480 ;
    END
  END gpio2_in[7]
  PIN gpio2_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1496.040 2722.000 1496.640 ;
    END
  END gpio2_oeb[0]
  PIN gpio2_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1565.400 2722.000 1566.000 ;
    END
  END gpio2_oeb[1]
  PIN gpio2_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1634.760 2722.000 1635.360 ;
    END
  END gpio2_oeb[2]
  PIN gpio2_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1704.120 2722.000 1704.720 ;
    END
  END gpio2_oeb[3]
  PIN gpio2_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2074.040 2722.000 2074.640 ;
    END
  END gpio2_oeb[4]
  PIN gpio2_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2143.400 2722.000 2144.000 ;
    END
  END gpio2_oeb[5]
  PIN gpio2_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2212.760 2722.000 2213.360 ;
    END
  END gpio2_oeb[6]
  PIN gpio2_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2282.120 2722.000 2282.720 ;
    END
  END gpio2_oeb[7]
  PIN gpio2_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1472.920 2722.000 1473.520 ;
    END
  END gpio2_out[0]
  PIN gpio2_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1542.280 2722.000 1542.880 ;
    END
  END gpio2_out[1]
  PIN gpio2_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1611.640 2722.000 1612.240 ;
    END
  END gpio2_out[2]
  PIN gpio2_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 1681.000 2722.000 1681.600 ;
    END
  END gpio2_out[3]
  PIN gpio2_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2050.920 2722.000 2051.520 ;
    END
  END gpio2_out[4]
  PIN gpio2_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2120.280 2722.000 2120.880 ;
    END
  END gpio2_out[5]
  PIN gpio2_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2189.640 2722.000 2190.240 ;
    END
  END gpio2_out[6]
  PIN gpio2_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2716.000 2259.000 2722.000 2259.600 ;
    END
  END gpio2_out[7]
  PIN gpio3_0_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1751.885 2298.500 1752.525 2300.000 ;
    END
  END gpio3_0_analog
  PIN gpio3_1_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1749.325 2298.500 1749.965 2300.000 ;
    END
  END gpio3_1_analog
  PIN gpio3_2_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1746.765 2298.500 1747.405 2300.000 ;
    END
  END gpio3_2_analog
  PIN gpio3_3_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1744.205 2298.500 1744.845 2300.000 ;
    END
  END gpio3_3_analog
  PIN gpio3_4_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1741.645 2298.500 1742.285 2300.000 ;
    END
  END gpio3_4_analog
  PIN gpio3_5_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1739.085 2298.500 1739.725 2300.000 ;
    END
  END gpio3_5_analog
  PIN gpio3_6_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1736.525 2298.500 1737.165 2300.000 ;
    END
  END gpio3_6_analog
  PIN gpio3_7_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1733.965 2298.500 1734.605 2300.000 ;
    END
  END gpio3_7_analog
  PIN gpio3_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2657.050 2296.000 2657.330 2302.000 ;
    END
  END gpio3_in[0]
  PIN gpio3_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2629.450 2296.000 2629.730 2302.000 ;
    END
  END gpio3_in[1]
  PIN gpio3_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2601.850 2296.000 2602.130 2302.000 ;
    END
  END gpio3_in[2]
  PIN gpio3_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2574.250 2296.000 2574.530 2302.000 ;
    END
  END gpio3_in[3]
  PIN gpio3_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2546.650 2296.000 2546.930 2302.000 ;
    END
  END gpio3_in[4]
  PIN gpio3_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2519.050 2296.000 2519.330 2302.000 ;
    END
  END gpio3_in[5]
  PIN gpio3_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2491.450 2296.000 2491.730 2302.000 ;
    END
  END gpio3_in[6]
  PIN gpio3_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2463.850 2296.000 2464.130 2302.000 ;
    END
  END gpio3_in[7]
  PIN gpio3_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.650 2296.000 2638.930 2302.000 ;
    END
  END gpio3_oeb[0]
  PIN gpio3_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2611.050 2296.000 2611.330 2302.000 ;
    END
  END gpio3_oeb[1]
  PIN gpio3_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2583.450 2296.000 2583.730 2302.000 ;
    END
  END gpio3_oeb[2]
  PIN gpio3_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2555.850 2296.000 2556.130 2302.000 ;
    END
  END gpio3_oeb[3]
  PIN gpio3_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2528.250 2296.000 2528.530 2302.000 ;
    END
  END gpio3_oeb[4]
  PIN gpio3_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.650 2296.000 2500.930 2302.000 ;
    END
  END gpio3_oeb[5]
  PIN gpio3_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.050 2296.000 2473.330 2302.000 ;
    END
  END gpio3_oeb[6]
  PIN gpio3_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2445.450 2296.000 2445.730 2302.000 ;
    END
  END gpio3_oeb[7]
  PIN gpio3_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2647.850 2296.000 2648.130 2302.000 ;
    END
  END gpio3_out[0]
  PIN gpio3_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2620.250 2296.000 2620.530 2302.000 ;
    END
  END gpio3_out[1]
  PIN gpio3_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2592.650 2296.000 2592.930 2302.000 ;
    END
  END gpio3_out[2]
  PIN gpio3_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2565.050 2296.000 2565.330 2302.000 ;
    END
  END gpio3_out[3]
  PIN gpio3_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2537.450 2296.000 2537.730 2302.000 ;
    END
  END gpio3_out[4]
  PIN gpio3_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2509.850 2296.000 2510.130 2302.000 ;
    END
  END gpio3_out[5]
  PIN gpio3_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2482.250 2296.000 2482.530 2302.000 ;
    END
  END gpio3_out[6]
  PIN gpio3_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2454.650 2296.000 2454.930 2302.000 ;
    END
  END gpio3_out[7]
  PIN gpio4_0_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1731.405 2298.500 1732.045 2300.000 ;
    END
  END gpio4_0_analog
  PIN gpio4_1_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1728.845 2298.500 1729.485 2300.000 ;
    END
  END gpio4_1_analog
  PIN gpio4_2_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1726.285 2298.500 1726.925 2300.000 ;
    END
  END gpio4_2_analog
  PIN gpio4_3_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1723.725 2298.500 1724.365 2300.000 ;
    END
  END gpio4_3_analog
  PIN gpio4_4_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1721.165 2298.500 1721.805 2300.000 ;
    END
  END gpio4_4_analog
  PIN gpio4_5_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1718.605 2298.500 1719.245 2300.000 ;
    END
  END gpio4_5_analog
  PIN gpio4_6_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1716.045 2298.500 1716.685 2300.000 ;
    END
  END gpio4_6_analog
  PIN gpio4_7_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1713.485 2298.500 1714.125 2300.000 ;
    END
  END gpio4_7_analog
  PIN gpio4_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 2296.000 274.530 2302.000 ;
    END
  END gpio4_in[0]
  PIN gpio4_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 2296.000 246.930 2302.000 ;
    END
  END gpio4_in[1]
  PIN gpio4_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 2296.000 219.330 2302.000 ;
    END
  END gpio4_in[2]
  PIN gpio4_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 2296.000 191.730 2302.000 ;
    END
  END gpio4_in[3]
  PIN gpio4_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 2296.000 164.130 2302.000 ;
    END
  END gpio4_in[4]
  PIN gpio4_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 2296.000 136.530 2302.000 ;
    END
  END gpio4_in[5]
  PIN gpio4_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 2296.000 108.930 2302.000 ;
    END
  END gpio4_in[6]
  PIN gpio4_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 2296.000 81.330 2302.000 ;
    END
  END gpio4_in[7]
  PIN gpio4_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 2296.000 256.130 2302.000 ;
    END
  END gpio4_oeb[0]
  PIN gpio4_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 2296.000 228.530 2302.000 ;
    END
  END gpio4_oeb[1]
  PIN gpio4_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 2296.000 200.930 2302.000 ;
    END
  END gpio4_oeb[2]
  PIN gpio4_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 2296.000 173.330 2302.000 ;
    END
  END gpio4_oeb[3]
  PIN gpio4_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 2296.000 145.730 2302.000 ;
    END
  END gpio4_oeb[4]
  PIN gpio4_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 2296.000 118.130 2302.000 ;
    END
  END gpio4_oeb[5]
  PIN gpio4_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 2296.000 90.530 2302.000 ;
    END
  END gpio4_oeb[6]
  PIN gpio4_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 2296.000 62.930 2302.000 ;
    END
  END gpio4_oeb[7]
  PIN gpio4_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 2296.000 265.330 2302.000 ;
    END
  END gpio4_out[0]
  PIN gpio4_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 2296.000 237.730 2302.000 ;
    END
  END gpio4_out[1]
  PIN gpio4_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 2296.000 210.130 2302.000 ;
    END
  END gpio4_out[2]
  PIN gpio4_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 2296.000 182.530 2302.000 ;
    END
  END gpio4_out[3]
  PIN gpio4_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 2296.000 154.930 2302.000 ;
    END
  END gpio4_out[4]
  PIN gpio4_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 2296.000 127.330 2302.000 ;
    END
  END gpio4_out[5]
  PIN gpio4_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 2296.000 99.730 2302.000 ;
    END
  END gpio4_out[6]
  PIN gpio4_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 2296.000 72.130 2302.000 ;
    END
  END gpio4_out[7]
  PIN gpio5_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2284.120 4.000 2284.720 ;
    END
  END gpio5_in[0]
  PIN gpio5_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2214.760 4.000 2215.360 ;
    END
  END gpio5_in[1]
  PIN gpio5_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2145.400 4.000 2146.000 ;
    END
  END gpio5_in[2]
  PIN gpio5_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2076.040 4.000 2076.640 ;
    END
  END gpio5_in[3]
  PIN gpio5_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1704.120 4.000 1704.720 ;
    END
  END gpio5_in[4]
  PIN gpio5_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1634.760 4.000 1635.360 ;
    END
  END gpio5_in[5]
  PIN gpio5_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1565.400 4.000 1566.000 ;
    END
  END gpio5_in[6]
  PIN gpio5_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1496.040 4.000 1496.640 ;
    END
  END gpio5_in[7]
  PIN gpio5_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2237.880 4.000 2238.480 ;
    END
  END gpio5_oeb[0]
  PIN gpio5_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2168.520 4.000 2169.120 ;
    END
  END gpio5_oeb[1]
  PIN gpio5_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2099.160 4.000 2099.760 ;
    END
  END gpio5_oeb[2]
  PIN gpio5_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2029.800 4.000 2030.400 ;
    END
  END gpio5_oeb[3]
  PIN gpio5_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1657.880 4.000 1658.480 ;
    END
  END gpio5_oeb[4]
  PIN gpio5_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1588.520 4.000 1589.120 ;
    END
  END gpio5_oeb[5]
  PIN gpio5_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1519.160 4.000 1519.760 ;
    END
  END gpio5_oeb[6]
  PIN gpio5_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1449.800 4.000 1450.400 ;
    END
  END gpio5_oeb[7]
  PIN gpio5_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2261.000 4.000 2261.600 ;
    END
  END gpio5_out[0]
  PIN gpio5_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2191.640 4.000 2192.240 ;
    END
  END gpio5_out[1]
  PIN gpio5_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2122.280 4.000 2122.880 ;
    END
  END gpio5_out[2]
  PIN gpio5_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 2052.920 4.000 2053.520 ;
    END
  END gpio5_out[3]
  PIN gpio5_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1681.000 4.000 1681.600 ;
    END
  END gpio5_out[4]
  PIN gpio5_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1611.640 4.000 1612.240 ;
    END
  END gpio5_out[5]
  PIN gpio5_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1542.280 4.000 1542.880 ;
    END
  END gpio5_out[6]
  PIN gpio5_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1472.920 4.000 1473.520 ;
    END
  END gpio5_out[7]
  PIN gpio6_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1426.680 4.000 1427.280 ;
    END
  END gpio6_in[0]
  PIN gpio6_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1357.320 4.000 1357.920 ;
    END
  END gpio6_in[1]
  PIN gpio6_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1287.960 4.000 1288.560 ;
    END
  END gpio6_in[2]
  PIN gpio6_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1218.600 4.000 1219.200 ;
    END
  END gpio6_in[3]
  PIN gpio6_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1149.240 4.000 1149.840 ;
    END
  END gpio6_in[4]
  PIN gpio6_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1079.880 4.000 1080.480 ;
    END
  END gpio6_in[5]
  PIN gpio6_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 1010.520 4.000 1011.120 ;
    END
  END gpio6_in[6]
  PIN gpio6_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 941.160 4.000 941.760 ;
    END
  END gpio6_in[7]
  PIN gpio6_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1380.440 4.000 1381.040 ;
    END
  END gpio6_oeb[0]
  PIN gpio6_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1311.080 4.000 1311.680 ;
    END
  END gpio6_oeb[1]
  PIN gpio6_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1241.720 4.000 1242.320 ;
    END
  END gpio6_oeb[2]
  PIN gpio6_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1172.360 4.000 1172.960 ;
    END
  END gpio6_oeb[3]
  PIN gpio6_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1103.000 4.000 1103.600 ;
    END
  END gpio6_oeb[4]
  PIN gpio6_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1033.640 4.000 1034.240 ;
    END
  END gpio6_oeb[5]
  PIN gpio6_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 964.280 4.000 964.880 ;
    END
  END gpio6_oeb[6]
  PIN gpio6_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 894.920 4.000 895.520 ;
    END
  END gpio6_oeb[7]
  PIN gpio6_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1403.560 4.000 1404.160 ;
    END
  END gpio6_out[0]
  PIN gpio6_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1334.200 4.000 1334.800 ;
    END
  END gpio6_out[1]
  PIN gpio6_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1264.840 4.000 1265.440 ;
    END
  END gpio6_out[2]
  PIN gpio6_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1195.480 4.000 1196.080 ;
    END
  END gpio6_out[3]
  PIN gpio6_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1126.120 4.000 1126.720 ;
    END
  END gpio6_out[4]
  PIN gpio6_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 1056.760 4.000 1057.360 ;
    END
  END gpio6_out[5]
  PIN gpio6_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 987.400 4.000 988.000 ;
    END
  END gpio6_out[6]
  PIN gpio6_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -2.000 918.040 4.000 918.640 ;
    END
  END gpio6_out[7]
  PIN gpio7_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 870.320 4.000 870.920 ;
    END
  END gpio7_in[0]
  PIN gpio7_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 800.960 4.000 801.560 ;
    END
  END gpio7_in[1]
  PIN gpio7_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 731.600 4.000 732.200 ;
    END
  END gpio7_in[2]
  PIN gpio7_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 571.240 4.000 571.840 ;
    END
  END gpio7_in[3]
  PIN gpio7_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 501.880 4.000 502.480 ;
    END
  END gpio7_in[4]
  PIN gpio7_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 432.520 4.000 433.120 ;
    END
  END gpio7_in[5]
  PIN gpio7_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 363.160 4.000 363.760 ;
    END
  END gpio7_in[6]
  PIN gpio7_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 293.800 4.000 294.400 ;
    END
  END gpio7_in[7]
  PIN gpio7_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 824.080 4.000 824.680 ;
    END
  END gpio7_oeb[0]
  PIN gpio7_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 754.720 4.000 755.320 ;
    END
  END gpio7_oeb[1]
  PIN gpio7_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 594.360 4.000 594.960 ;
    END
  END gpio7_oeb[2]
  PIN gpio7_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 525.000 4.000 525.600 ;
    END
  END gpio7_oeb[3]
  PIN gpio7_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 455.640 4.000 456.240 ;
    END
  END gpio7_oeb[4]
  PIN gpio7_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 386.280 4.000 386.880 ;
    END
  END gpio7_oeb[5]
  PIN gpio7_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 316.920 4.000 317.520 ;
    END
  END gpio7_oeb[6]
  PIN gpio7_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 247.560 4.000 248.160 ;
    END
  END gpio7_oeb[7]
  PIN gpio7_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 847.200 4.000 847.800 ;
    END
  END gpio7_out[0]
  PIN gpio7_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 777.840 4.000 778.440 ;
    END
  END gpio7_out[1]
  PIN gpio7_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 617.480 4.000 618.080 ;
    END
  END gpio7_out[2]
  PIN gpio7_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 548.120 4.000 548.720 ;
    END
  END gpio7_out[3]
  PIN gpio7_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 478.760 4.000 479.360 ;
    END
  END gpio7_out[4]
  PIN gpio7_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 409.400 4.000 410.000 ;
    END
  END gpio7_out[5]
  PIN gpio7_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 340.040 4.000 340.640 ;
    END
  END gpio7_out[6]
  PIN gpio7_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -2.000 270.680 4.000 271.280 ;
    END
  END gpio7_out[7]
  PIN ibias100
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1695.565 2298.500 1696.205 2300.000 ;
    END
  END ibias100
  PIN ibias50
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1693.005 2298.500 1693.645 2300.000 ;
    END
  END ibias50
  PIN left_vref
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1675.085 2298.500 1675.725 2300.000 ;
    END
  END left_vref
  PIN right_vref
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1677.645 2298.500 1678.285 2300.000 ;
    END
  END right_vref
  PIN sio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2445.970 -2.000 2446.250 4.000 ;
    END
  END sio_in[0]
  PIN sio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2469.430 -2.000 2469.710 4.000 ;
    END
  END sio_in[1]
  PIN sio_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.610 -2.000 2461.890 4.000 ;
    END
  END sio_oeb[0]
  PIN sio_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.070 -2.000 2485.350 4.000 ;
    END
  END sio_oeb[1]
  PIN sio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2453.790 -2.000 2454.070 4.000 ;
    END
  END sio_out[0]
  PIN sio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2477.250 -2.000 2477.530 4.000 ;
    END
  END sio_out[1]
  PIN tempsense
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1680.205 2298.500 1680.845 2300.000 ;
    END
  END tempsense
  PIN ulpcomp_n
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1708.365 2298.500 1709.005 2300.000 ;
    END
  END ulpcomp_n
  PIN ulpcomp_p
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1710.925 2298.500 1711.565 2300.000 ;
    END
  END ulpcomp_p
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.390 -2.000 1071.670 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.590 -2.000 1149.870 4.000 ;
    END
  END user_irq[10]
  PIN user_irq[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.410 -2.000 1157.690 4.000 ;
    END
  END user_irq[11]
  PIN user_irq[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.230 -2.000 1165.510 4.000 ;
    END
  END user_irq[12]
  PIN user_irq[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.050 -2.000 1173.330 4.000 ;
    END
  END user_irq[13]
  PIN user_irq[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.870 -2.000 1181.150 4.000 ;
    END
  END user_irq[14]
  PIN user_irq[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.690 -2.000 1188.970 4.000 ;
    END
  END user_irq[15]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.210 -2.000 1079.490 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.030 -2.000 1087.310 4.000 ;
    END
  END user_irq[2]
  PIN user_irq[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.850 -2.000 1095.130 4.000 ;
    END
  END user_irq[3]
  PIN user_irq[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.670 -2.000 1102.950 4.000 ;
    END
  END user_irq[4]
  PIN user_irq[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.490 -2.000 1110.770 4.000 ;
    END
  END user_irq[5]
  PIN user_irq[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.310 -2.000 1118.590 4.000 ;
    END
  END user_irq[6]
  PIN user_irq[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.130 -2.000 1126.410 4.000 ;
    END
  END user_irq[7]
  PIN user_irq[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.950 -2.000 1134.230 4.000 ;
    END
  END user_irq[8]
  PIN user_irq[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.770 -2.000 1142.050 4.000 ;
    END
  END user_irq[9]
  PIN vbgsc
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1690.445 2298.500 1691.085 2300.000 ;
    END
  END vbgsc
  PIN vbgtc
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1687.885 2298.500 1688.525 2300.000 ;
    END
  END vbgtc
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -7.980 -7.220 -4.880 2305.620 ;
    END
    PORT
      LAYER met5 ;
        RECT -7.980 -7.220 2727.960 -4.120 ;
    END
    PORT
      LAYER met5 ;
        RECT -7.980 2302.520 2727.960 2305.620 ;
    END
    PORT
      LAYER met4 ;
        RECT 2724.860 -7.220 2727.960 2305.620 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.570 4.400 26.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.570 4.400 116.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.570 4.400 206.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 293.570 -21.620 296.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.570 -21.620 386.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.570 -21.620 476.670 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.570 298.620 476.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 -21.620 566.670 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.570 293.145 566.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.570 -21.620 656.670 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.570 293.145 656.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 -21.620 746.670 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.570 293.145 746.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 833.570 -21.620 836.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.570 -21.620 926.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.570 -21.620 1016.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.570 -21.620 1106.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1193.570 -21.620 1196.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.570 -21.620 1286.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.570 -21.620 1376.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.570 -21.620 1466.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1553.570 -21.620 1556.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1643.570 -21.620 1646.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.570 -21.620 1736.670 2292.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1823.570 -21.620 1826.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.570 -21.620 1916.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2003.570 -21.620 2006.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2093.570 -21.620 2096.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2183.570 -21.620 2186.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2273.570 -21.620 2276.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2363.570 -21.620 2366.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2453.570 -21.620 2456.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2543.570 4.400 2546.670 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2633.570 4.400 2636.670 2320.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 24.330 2742.360 27.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 114.330 461.980 117.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 204.330 2742.360 207.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 294.330 2742.360 297.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 384.330 2742.360 387.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 474.330 2742.360 477.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 564.330 2742.360 567.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 654.330 2742.360 657.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 744.330 2742.360 747.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 834.330 2742.360 837.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 924.330 2742.360 927.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1014.330 2742.360 1017.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1104.330 2742.360 1107.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1194.330 2742.360 1197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1284.330 2742.360 1287.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1374.330 2742.360 1377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1464.330 2742.360 1467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1554.330 2742.360 1557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1644.330 2742.360 1647.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1734.330 2742.360 1737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1824.330 2742.360 1827.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1914.330 2742.360 1917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2004.330 2742.360 2007.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2094.330 2742.360 2097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2184.330 2742.360 2187.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2274.330 2742.360 2277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 832.700 114.330 2742.360 117.430 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -17.580 -16.820 -14.480 2315.220 ;
    END
    PORT
      LAYER met5 ;
        RECT -17.580 -16.820 2737.560 -13.720 ;
    END
    PORT
      LAYER met5 ;
        RECT -17.580 2312.120 2737.560 2315.220 ;
    END
    PORT
      LAYER met4 ;
        RECT 2734.460 -16.820 2737.560 2315.220 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.770 4.400 63.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 150.770 4.400 153.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 240.770 -21.620 243.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 330.770 -21.620 333.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 420.770 -21.620 423.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 510.770 -21.620 513.870 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 510.770 293.145 513.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 600.770 -21.620 603.870 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 600.770 293.145 603.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 690.770 -21.620 693.870 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 690.770 293.145 693.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 780.770 -21.620 783.870 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 780.770 298.620 783.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 870.770 -21.620 873.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 960.770 -21.620 963.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1050.770 -21.620 1053.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1140.770 -21.620 1143.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1230.770 -21.620 1233.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1320.770 -21.620 1323.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.770 -21.620 1413.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1500.770 -21.620 1503.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1590.770 -21.620 1593.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1680.770 -21.620 1683.870 2292.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1770.770 -21.620 1773.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1860.770 -21.620 1863.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1950.770 -21.620 1953.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2040.770 -21.620 2043.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2130.770 -21.620 2133.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2220.770 -21.620 2223.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2310.770 -21.620 2313.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2400.770 -21.620 2403.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2490.770 -21.620 2493.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2580.770 4.400 2583.870 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2670.770 4.400 2673.870 2320.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 61.530 2742.360 64.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 151.530 461.980 154.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 241.530 2742.360 244.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 331.530 2742.360 334.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 421.530 2742.360 424.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 511.530 2742.360 514.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 601.530 2742.360 604.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 691.530 2742.360 694.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 781.530 2742.360 784.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 871.530 2742.360 874.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 961.530 2742.360 964.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1051.530 2742.360 1054.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1141.530 2742.360 1144.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1231.530 2742.360 1234.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1321.530 2742.360 1324.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1411.530 2742.360 1414.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1501.530 2742.360 1504.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1591.530 2742.360 1594.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1681.530 2742.360 1684.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1771.530 2742.360 1774.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1861.530 2742.360 1864.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1951.530 2742.360 1954.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2041.530 2742.360 2044.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2131.530 2742.360 2134.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2221.530 2742.360 2224.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 832.700 151.530 2742.360 154.630 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 2716.780 1722.860 2720.000 1746.760 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 2716.780 1772.755 2720.000 1796.655 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2501.510 0.000 2525.410 3.190 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2551.405 0.000 2575.305 3.190 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 1786.540 3.220 1810.440 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 1736.645 3.220 1760.545 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 144.695 0.000 168.595 3.190 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 194.590 0.000 218.490 3.190 ;
    END
  END vdda2
  PIN vinref
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1672.525 2298.500 1673.165 2300.000 ;
    END
  END vinref
  PIN voutref
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1669.965 2298.500 1670.605 2300.000 ;
    END
  END voutref
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 2716.780 1892.750 2720.000 1916.650 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 2716.780 1842.855 2720.000 1866.755 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2671.405 0.000 2695.305 3.190 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2621.510 0.000 2645.410 3.190 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 1901.540 3.220 1925.440 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 1851.645 3.220 1875.545 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 74.590 0.000 98.490 3.190 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.695 0.000 48.595 3.190 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -12.780 -12.020 -9.680 2310.420 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.780 -12.020 2732.760 -8.920 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.780 2307.320 2732.760 2310.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 2729.660 -12.020 2732.760 2310.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 42.170 4.400 45.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.170 4.400 135.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 222.170 4.400 225.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 312.170 -21.620 315.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 402.170 -21.620 405.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 492.170 -21.620 495.270 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 492.170 293.145 495.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 582.170 -21.620 585.270 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 582.170 293.145 585.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 672.170 -21.620 675.270 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 672.170 293.145 675.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 762.170 -21.620 765.270 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 762.170 293.145 765.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 852.170 -21.620 855.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.170 -21.620 945.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.170 -21.620 1035.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1122.170 -21.620 1125.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1212.170 -21.620 1215.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1302.170 -21.620 1305.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1392.170 -21.620 1395.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1482.170 -21.620 1485.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1572.170 -21.620 1575.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.170 -21.620 1665.270 2292.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1752.170 -21.620 1755.270 2292.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1842.170 -21.620 1845.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.170 -21.620 1935.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2022.170 -21.620 2025.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2112.170 -21.620 2115.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2202.170 -21.620 2205.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2292.170 -21.620 2295.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2382.170 -21.620 2385.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2472.170 -21.620 2475.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2562.170 4.400 2565.270 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2652.170 4.400 2655.270 2320.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 42.930 2742.360 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 132.930 461.980 136.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 222.930 2742.360 226.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 312.930 2742.360 316.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 402.930 2742.360 406.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 492.930 2742.360 496.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 582.930 2742.360 586.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 672.930 2742.360 676.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 762.930 2742.360 766.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 852.930 2742.360 856.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 942.930 2742.360 946.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1032.930 2742.360 1036.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1122.930 2742.360 1126.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1212.930 2742.360 1216.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1302.930 2742.360 1306.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1392.930 2742.360 1396.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1482.930 2742.360 1486.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1572.930 2742.360 1576.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1662.930 2742.360 1666.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1752.930 2742.360 1756.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1842.930 2742.360 1846.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1932.930 2742.360 1936.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2022.930 2742.360 2026.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2112.930 2742.360 2116.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2202.930 2742.360 2206.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 832.700 132.930 2742.360 136.030 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -22.380 -21.620 -19.280 2320.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 -21.620 2742.360 -18.520 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2316.920 2742.360 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2739.260 -21.620 2742.360 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.370 4.400 82.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 169.370 4.400 172.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 259.370 -21.620 262.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 349.370 -21.620 352.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 439.370 -21.620 442.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 529.370 -21.620 532.470 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 529.370 293.145 532.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 619.370 -21.620 622.470 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 619.370 293.145 622.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 709.370 -21.620 712.470 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 709.370 293.145 712.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 799.370 -21.620 802.470 94.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 799.370 293.145 802.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 889.370 -21.620 892.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 979.370 -21.620 982.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1069.370 -21.620 1072.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1159.370 -21.620 1162.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.370 -21.620 1252.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1339.370 -21.620 1342.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1429.370 -21.620 1432.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1519.370 -21.620 1522.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1609.370 -21.620 1612.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1699.370 -21.620 1702.470 2292.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1789.370 -21.620 1792.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1879.370 -21.620 1882.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1969.370 -21.620 1972.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2059.370 -21.620 2062.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2149.370 -21.620 2152.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2239.370 -21.620 2242.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2329.370 -21.620 2332.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2419.370 -21.620 2422.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2509.370 4.400 2512.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2599.370 4.400 2602.470 2320.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2689.370 4.400 2692.470 2320.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 80.130 2742.360 83.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 170.130 2742.360 173.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 260.130 2742.360 263.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 350.130 2742.360 353.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 440.130 2742.360 443.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 530.130 2742.360 533.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 620.130 2742.360 623.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 710.130 2742.360 713.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 800.130 2742.360 803.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 890.130 2742.360 893.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 980.130 2742.360 983.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1070.130 2742.360 1073.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1160.130 2742.360 1163.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1250.130 2742.360 1253.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1340.130 2742.360 1343.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1430.130 2742.360 1433.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1520.130 2742.360 1523.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1610.130 2742.360 1613.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1700.130 2742.360 1703.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1790.130 2742.360 1793.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1880.130 2742.360 1883.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 1970.130 2742.360 1973.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2060.130 2742.360 2063.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2150.130 2742.360 2153.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -22.380 2240.130 2742.360 2243.230 ;
    END
  END vssd2
  OBS
      LAYER nwell ;
        RECT 459.930 110.795 839.810 287.870 ;
      LAYER li1 ;
        RECT 460.120 110.795 839.620 287.765 ;
      LAYER met1 ;
        RECT 460.120 0.040 1063.450 287.920 ;
      LAYER met2 ;
        RECT 0.550 4.280 2716.670 1427.165 ;
        RECT 0.550 0.010 234.370 4.280 ;
        RECT 235.210 0.010 242.190 4.280 ;
        RECT 243.030 0.010 250.010 4.280 ;
        RECT 250.850 0.010 257.830 4.280 ;
        RECT 258.670 0.010 265.650 4.280 ;
        RECT 266.490 0.010 273.470 4.280 ;
        RECT 274.310 0.010 281.290 4.280 ;
        RECT 282.130 0.010 289.110 4.280 ;
        RECT 289.950 0.010 296.930 4.280 ;
        RECT 297.770 0.010 304.750 4.280 ;
        RECT 305.590 0.010 312.570 4.280 ;
        RECT 313.410 0.010 320.390 4.280 ;
        RECT 321.230 0.010 328.210 4.280 ;
        RECT 329.050 0.010 336.030 4.280 ;
        RECT 336.870 0.010 343.850 4.280 ;
        RECT 344.690 0.010 351.670 4.280 ;
        RECT 352.510 0.010 359.490 4.280 ;
        RECT 360.330 0.010 367.310 4.280 ;
        RECT 368.150 0.010 375.130 4.280 ;
        RECT 375.970 0.010 382.950 4.280 ;
        RECT 383.790 0.010 390.770 4.280 ;
        RECT 391.610 0.010 398.590 4.280 ;
        RECT 399.430 0.010 406.410 4.280 ;
        RECT 407.250 0.010 414.230 4.280 ;
        RECT 415.070 0.010 422.050 4.280 ;
        RECT 422.890 0.010 429.870 4.280 ;
        RECT 430.710 0.010 437.690 4.280 ;
        RECT 438.530 0.010 445.510 4.280 ;
        RECT 446.350 0.010 453.330 4.280 ;
        RECT 454.170 0.010 461.150 4.280 ;
        RECT 461.990 0.010 468.970 4.280 ;
        RECT 469.810 0.010 476.790 4.280 ;
        RECT 477.630 0.010 484.610 4.280 ;
        RECT 485.450 0.010 492.430 4.280 ;
        RECT 493.270 0.010 500.250 4.280 ;
        RECT 501.090 0.010 508.070 4.280 ;
        RECT 508.910 0.010 515.890 4.280 ;
        RECT 516.730 0.010 523.710 4.280 ;
        RECT 524.550 0.010 531.530 4.280 ;
        RECT 532.370 0.010 539.350 4.280 ;
        RECT 540.190 0.010 547.170 4.280 ;
        RECT 548.010 0.010 554.990 4.280 ;
        RECT 555.830 0.010 562.810 4.280 ;
        RECT 563.650 0.010 570.630 4.280 ;
        RECT 571.470 0.010 578.450 4.280 ;
        RECT 579.290 0.010 586.270 4.280 ;
        RECT 587.110 0.010 594.090 4.280 ;
        RECT 594.930 0.010 601.910 4.280 ;
        RECT 602.750 0.010 609.730 4.280 ;
        RECT 610.570 0.010 617.550 4.280 ;
        RECT 618.390 0.010 625.370 4.280 ;
        RECT 626.210 0.010 633.190 4.280 ;
        RECT 634.030 0.010 641.010 4.280 ;
        RECT 641.850 0.010 648.830 4.280 ;
        RECT 649.670 0.010 656.650 4.280 ;
        RECT 657.490 0.010 664.470 4.280 ;
        RECT 665.310 0.010 672.290 4.280 ;
        RECT 673.130 0.010 680.110 4.280 ;
        RECT 680.950 0.010 687.930 4.280 ;
        RECT 688.770 0.010 695.750 4.280 ;
        RECT 696.590 0.010 703.570 4.280 ;
        RECT 704.410 0.010 711.390 4.280 ;
        RECT 712.230 0.010 719.210 4.280 ;
        RECT 720.050 0.010 727.030 4.280 ;
        RECT 727.870 0.010 734.850 4.280 ;
        RECT 735.690 0.010 742.670 4.280 ;
        RECT 743.510 0.010 750.490 4.280 ;
        RECT 751.330 0.010 758.310 4.280 ;
        RECT 759.150 0.010 766.130 4.280 ;
        RECT 766.970 0.010 773.950 4.280 ;
        RECT 774.790 0.010 781.770 4.280 ;
        RECT 782.610 0.010 789.590 4.280 ;
        RECT 790.430 0.010 797.410 4.280 ;
        RECT 798.250 0.010 805.230 4.280 ;
        RECT 806.070 0.010 813.050 4.280 ;
        RECT 813.890 0.010 820.870 4.280 ;
        RECT 821.710 0.010 828.690 4.280 ;
        RECT 829.530 0.010 836.510 4.280 ;
        RECT 837.350 0.010 844.330 4.280 ;
        RECT 845.170 0.010 852.150 4.280 ;
        RECT 852.990 0.010 859.970 4.280 ;
        RECT 860.810 0.010 867.790 4.280 ;
        RECT 868.630 0.010 875.610 4.280 ;
        RECT 876.450 0.010 883.430 4.280 ;
        RECT 884.270 0.010 891.250 4.280 ;
        RECT 892.090 0.010 899.070 4.280 ;
        RECT 899.910 0.010 906.890 4.280 ;
        RECT 907.730 0.010 914.710 4.280 ;
        RECT 915.550 0.010 922.530 4.280 ;
        RECT 923.370 0.010 930.350 4.280 ;
        RECT 931.190 0.010 938.170 4.280 ;
        RECT 939.010 0.010 945.990 4.280 ;
        RECT 946.830 0.010 953.810 4.280 ;
        RECT 954.650 0.010 961.630 4.280 ;
        RECT 962.470 0.010 969.450 4.280 ;
        RECT 970.290 0.010 977.270 4.280 ;
        RECT 978.110 0.010 985.090 4.280 ;
        RECT 985.930 0.010 992.910 4.280 ;
        RECT 993.750 0.010 1000.730 4.280 ;
        RECT 1001.570 0.010 1008.550 4.280 ;
        RECT 1009.390 0.010 1016.370 4.280 ;
        RECT 1017.210 0.010 1024.190 4.280 ;
        RECT 1025.030 0.010 1032.010 4.280 ;
        RECT 1032.850 0.010 1039.830 4.280 ;
        RECT 1040.670 0.010 1047.650 4.280 ;
        RECT 1048.490 0.010 1055.470 4.280 ;
        RECT 1056.310 0.010 1063.290 4.280 ;
        RECT 1064.130 0.010 1071.110 4.280 ;
        RECT 1071.950 0.010 1078.930 4.280 ;
        RECT 1079.770 0.010 1086.750 4.280 ;
        RECT 1087.590 0.010 1094.570 4.280 ;
        RECT 1095.410 0.010 1102.390 4.280 ;
        RECT 1103.230 0.010 1110.210 4.280 ;
        RECT 1111.050 0.010 1118.030 4.280 ;
        RECT 1118.870 0.010 1125.850 4.280 ;
        RECT 1126.690 0.010 1133.670 4.280 ;
        RECT 1134.510 0.010 1141.490 4.280 ;
        RECT 1142.330 0.010 1149.310 4.280 ;
        RECT 1150.150 0.010 1157.130 4.280 ;
        RECT 1157.970 0.010 1164.950 4.280 ;
        RECT 1165.790 0.010 1172.770 4.280 ;
        RECT 1173.610 0.010 1180.590 4.280 ;
        RECT 1181.430 0.010 1188.410 4.280 ;
        RECT 1189.250 0.010 2445.690 4.280 ;
        RECT 2446.530 0.010 2453.510 4.280 ;
        RECT 2454.350 0.010 2461.330 4.280 ;
        RECT 2462.170 0.010 2469.150 4.280 ;
        RECT 2469.990 0.010 2476.970 4.280 ;
        RECT 2477.810 0.010 2484.790 4.280 ;
        RECT 2485.630 0.010 2716.670 4.280 ;
      LAYER met3 ;
        RECT 4.400 1426.280 2715.600 1427.145 ;
        RECT 0.270 1404.560 2716.695 1426.280 ;
        RECT 4.400 1403.160 2715.600 1404.560 ;
        RECT 0.270 1381.440 2716.695 1403.160 ;
        RECT 4.400 1380.040 2715.600 1381.440 ;
        RECT 0.270 1358.320 2716.695 1380.040 ;
        RECT 4.400 1356.920 2715.600 1358.320 ;
        RECT 0.270 1335.200 2716.695 1356.920 ;
        RECT 4.400 1333.800 2715.600 1335.200 ;
        RECT 0.270 1312.080 2716.695 1333.800 ;
        RECT 4.400 1310.680 2715.600 1312.080 ;
        RECT 0.270 1288.960 2716.695 1310.680 ;
        RECT 4.400 1287.560 2715.600 1288.960 ;
        RECT 0.270 1265.840 2716.695 1287.560 ;
        RECT 4.400 1264.440 2715.600 1265.840 ;
        RECT 0.270 1242.720 2716.695 1264.440 ;
        RECT 4.400 1241.320 2715.600 1242.720 ;
        RECT 0.270 1219.600 2716.695 1241.320 ;
        RECT 4.400 1218.200 2715.600 1219.600 ;
        RECT 0.270 1196.480 2716.695 1218.200 ;
        RECT 4.400 1195.080 2715.600 1196.480 ;
        RECT 0.270 1173.360 2716.695 1195.080 ;
        RECT 4.400 1171.960 2715.600 1173.360 ;
        RECT 0.270 1150.240 2716.695 1171.960 ;
        RECT 4.400 1148.840 2715.600 1150.240 ;
        RECT 0.270 1127.120 2716.695 1148.840 ;
        RECT 4.400 1125.720 2715.600 1127.120 ;
        RECT 0.270 1104.000 2716.695 1125.720 ;
        RECT 4.400 1102.600 2715.600 1104.000 ;
        RECT 0.270 1080.880 2716.695 1102.600 ;
        RECT 4.400 1079.480 2715.600 1080.880 ;
        RECT 0.270 1057.760 2716.695 1079.480 ;
        RECT 4.400 1056.360 2715.600 1057.760 ;
        RECT 0.270 1034.640 2716.695 1056.360 ;
        RECT 4.400 1033.240 2715.600 1034.640 ;
        RECT 0.270 1011.520 2716.695 1033.240 ;
        RECT 4.400 1010.120 2715.600 1011.520 ;
        RECT 0.270 988.400 2716.695 1010.120 ;
        RECT 4.400 987.000 2715.600 988.400 ;
        RECT 0.270 965.280 2716.695 987.000 ;
        RECT 4.400 963.880 2715.600 965.280 ;
        RECT 0.270 942.160 2716.695 963.880 ;
        RECT 4.400 940.760 2715.600 942.160 ;
        RECT 0.270 919.040 2716.695 940.760 ;
        RECT 4.400 917.640 2715.600 919.040 ;
        RECT 0.270 895.920 2716.695 917.640 ;
        RECT 4.400 894.520 2715.600 895.920 ;
        RECT 0.270 871.320 2716.695 894.520 ;
        RECT 4.400 869.920 2716.695 871.320 ;
        RECT 0.270 848.200 2716.695 869.920 ;
        RECT 4.400 846.800 2716.695 848.200 ;
        RECT 0.270 825.080 2716.695 846.800 ;
        RECT 4.400 823.680 2716.695 825.080 ;
        RECT 0.270 801.960 2716.695 823.680 ;
        RECT 4.400 800.560 2716.695 801.960 ;
        RECT 0.270 778.840 2716.695 800.560 ;
        RECT 4.400 777.440 2716.695 778.840 ;
        RECT 0.270 755.720 2716.695 777.440 ;
        RECT 4.400 754.320 2716.695 755.720 ;
        RECT 0.270 732.600 2716.695 754.320 ;
        RECT 4.400 731.200 2716.695 732.600 ;
        RECT 0.270 629.850 2716.695 731.200 ;
        RECT 0.270 628.450 2715.600 629.850 ;
        RECT 0.270 618.480 2716.695 628.450 ;
        RECT 4.400 617.080 2716.695 618.480 ;
        RECT 0.270 606.730 2716.695 617.080 ;
        RECT 0.270 605.330 2715.600 606.730 ;
        RECT 0.270 595.360 2716.695 605.330 ;
        RECT 4.400 593.960 2716.695 595.360 ;
        RECT 0.270 583.610 2716.695 593.960 ;
        RECT 0.270 582.210 2715.600 583.610 ;
        RECT 0.270 572.240 2716.695 582.210 ;
        RECT 4.400 570.840 2716.695 572.240 ;
        RECT 0.270 560.490 2716.695 570.840 ;
        RECT 0.270 559.090 2715.600 560.490 ;
        RECT 0.270 549.120 2716.695 559.090 ;
        RECT 4.400 547.720 2716.695 549.120 ;
        RECT 0.270 537.370 2716.695 547.720 ;
        RECT 0.270 535.970 2715.600 537.370 ;
        RECT 0.270 526.000 2716.695 535.970 ;
        RECT 4.400 524.600 2716.695 526.000 ;
        RECT 0.270 514.250 2716.695 524.600 ;
        RECT 0.270 512.850 2715.600 514.250 ;
        RECT 0.270 502.880 2716.695 512.850 ;
        RECT 4.400 501.480 2716.695 502.880 ;
        RECT 0.270 491.130 2716.695 501.480 ;
        RECT 0.270 489.730 2715.600 491.130 ;
        RECT 0.270 479.760 2716.695 489.730 ;
        RECT 4.400 478.360 2716.695 479.760 ;
        RECT 0.270 468.010 2716.695 478.360 ;
        RECT 0.270 466.610 2715.600 468.010 ;
        RECT 0.270 456.640 2716.695 466.610 ;
        RECT 4.400 455.240 2716.695 456.640 ;
        RECT 0.270 444.890 2716.695 455.240 ;
        RECT 0.270 443.490 2715.600 444.890 ;
        RECT 0.270 433.520 2716.695 443.490 ;
        RECT 4.400 432.120 2716.695 433.520 ;
        RECT 0.270 421.770 2716.695 432.120 ;
        RECT 0.270 420.370 2715.600 421.770 ;
        RECT 0.270 410.400 2716.695 420.370 ;
        RECT 4.400 409.000 2716.695 410.400 ;
        RECT 0.270 398.650 2716.695 409.000 ;
        RECT 0.270 397.250 2715.600 398.650 ;
        RECT 0.270 387.280 2716.695 397.250 ;
        RECT 4.400 385.880 2716.695 387.280 ;
        RECT 0.270 375.530 2716.695 385.880 ;
        RECT 0.270 374.130 2715.600 375.530 ;
        RECT 0.270 364.160 2716.695 374.130 ;
        RECT 4.400 362.760 2716.695 364.160 ;
        RECT 0.270 352.410 2716.695 362.760 ;
        RECT 0.270 351.010 2715.600 352.410 ;
        RECT 0.270 341.040 2716.695 351.010 ;
        RECT 4.400 339.640 2716.695 341.040 ;
        RECT 0.270 329.290 2716.695 339.640 ;
        RECT 0.270 327.890 2715.600 329.290 ;
        RECT 0.270 317.920 2716.695 327.890 ;
        RECT 4.400 316.520 2716.695 317.920 ;
        RECT 0.270 306.170 2716.695 316.520 ;
        RECT 0.270 304.770 2715.600 306.170 ;
        RECT 0.270 294.800 2716.695 304.770 ;
        RECT 4.400 293.400 2716.695 294.800 ;
        RECT 0.270 283.050 2716.695 293.400 ;
        RECT 0.270 281.650 2715.600 283.050 ;
        RECT 0.270 271.680 2716.695 281.650 ;
        RECT 4.400 270.280 2716.695 271.680 ;
        RECT 0.270 259.930 2716.695 270.280 ;
        RECT 0.270 258.530 2715.600 259.930 ;
        RECT 0.270 248.560 2716.695 258.530 ;
        RECT 4.400 247.160 2716.695 248.560 ;
        RECT 0.270 236.810 2716.695 247.160 ;
        RECT 0.270 235.410 2715.600 236.810 ;
        RECT 0.270 213.690 2716.695 235.410 ;
        RECT 0.270 212.290 2715.600 213.690 ;
        RECT 0.270 190.570 2716.695 212.290 ;
        RECT 0.270 189.170 2715.600 190.570 ;
        RECT 0.270 167.450 2716.695 189.170 ;
        RECT 0.270 166.050 2715.600 167.450 ;
        RECT 0.270 144.330 2716.695 166.050 ;
        RECT 0.270 142.930 2715.600 144.330 ;
        RECT 0.270 121.210 2716.695 142.930 ;
        RECT 0.270 119.810 2715.600 121.210 ;
        RECT 0.270 98.090 2716.695 119.810 ;
        RECT 0.270 96.690 2715.600 98.090 ;
        RECT 0.270 0.175 2716.695 96.690 ;
      LAYER met4 ;
        RECT 0.295 4.000 23.170 1402.665 ;
        RECT 27.070 4.000 41.770 1402.665 ;
        RECT 45.670 4.000 60.370 1402.665 ;
        RECT 64.270 4.000 78.970 1402.665 ;
        RECT 82.870 4.000 113.170 1402.665 ;
        RECT 117.070 4.000 131.770 1402.665 ;
        RECT 135.670 4.000 150.370 1402.665 ;
        RECT 154.270 4.000 168.970 1402.665 ;
        RECT 172.870 4.000 203.170 1402.665 ;
        RECT 207.070 4.000 221.770 1402.665 ;
        RECT 225.670 4.000 240.370 1402.665 ;
        RECT 0.295 3.590 240.370 4.000 ;
        RECT 0.295 1.110 24.295 3.590 ;
        RECT 48.995 1.110 74.190 3.590 ;
        RECT 98.890 1.110 144.295 3.590 ;
        RECT 168.995 1.110 194.190 3.590 ;
        RECT 218.890 1.110 240.370 3.590 ;
        RECT 244.270 1.110 258.970 1402.665 ;
        RECT 262.870 1.110 293.170 1402.665 ;
        RECT 297.070 1.110 311.770 1402.665 ;
        RECT 315.670 1.110 330.370 1402.665 ;
        RECT 334.270 1.110 348.970 1402.665 ;
        RECT 352.870 1.110 383.170 1402.665 ;
        RECT 387.070 1.110 401.770 1402.665 ;
        RECT 405.670 1.110 420.370 1402.665 ;
        RECT 424.270 1.110 438.970 1402.665 ;
        RECT 442.870 298.220 473.170 1402.665 ;
        RECT 477.070 298.220 491.770 1402.665 ;
        RECT 442.870 292.745 491.770 298.220 ;
        RECT 495.670 292.745 510.370 1402.665 ;
        RECT 514.270 292.745 528.970 1402.665 ;
        RECT 532.870 292.745 563.170 1402.665 ;
        RECT 567.070 292.745 581.770 1402.665 ;
        RECT 585.670 292.745 600.370 1402.665 ;
        RECT 604.270 292.745 618.970 1402.665 ;
        RECT 622.870 292.745 653.170 1402.665 ;
        RECT 657.070 292.745 671.770 1402.665 ;
        RECT 675.670 292.745 690.370 1402.665 ;
        RECT 694.270 292.745 708.970 1402.665 ;
        RECT 712.870 292.745 743.170 1402.665 ;
        RECT 747.070 292.745 761.770 1402.665 ;
        RECT 765.670 298.220 780.370 1402.665 ;
        RECT 784.270 298.220 798.970 1402.665 ;
        RECT 765.670 292.745 798.970 298.220 ;
        RECT 802.870 292.745 820.890 1402.665 ;
        RECT 442.870 94.935 820.890 292.745 ;
        RECT 442.870 1.110 473.170 94.935 ;
        RECT 477.070 1.110 491.770 94.935 ;
        RECT 495.670 1.110 510.370 94.935 ;
        RECT 514.270 1.110 528.970 94.935 ;
        RECT 532.870 1.110 563.170 94.935 ;
        RECT 567.070 1.110 581.770 94.935 ;
        RECT 585.670 1.110 600.370 94.935 ;
        RECT 604.270 1.110 618.970 94.935 ;
        RECT 622.870 1.110 653.170 94.935 ;
        RECT 657.070 1.110 671.770 94.935 ;
        RECT 675.670 1.110 690.370 94.935 ;
        RECT 694.270 1.110 708.970 94.935 ;
        RECT 712.870 1.110 743.170 94.935 ;
        RECT 747.070 1.110 761.770 94.935 ;
        RECT 765.670 1.110 780.370 94.935 ;
        RECT 784.270 1.110 798.970 94.935 ;
        RECT 802.870 1.110 820.890 94.935 ;
      LAYER met5 ;
        RECT 0.580 299.030 821.100 301.700 ;
        RECT 0.580 264.830 821.100 292.730 ;
        RECT 0.580 246.230 821.100 258.530 ;
        RECT 0.580 227.630 821.100 239.930 ;
        RECT 0.580 209.030 821.100 221.330 ;
        RECT 0.580 174.830 821.100 202.730 ;
        RECT 0.580 156.230 821.100 168.530 ;
        RECT 463.580 149.930 821.100 156.230 ;
        RECT 0.580 137.630 821.100 149.930 ;
        RECT 463.580 131.330 821.100 137.630 ;
        RECT 0.580 119.030 821.100 131.330 ;
        RECT 463.580 112.730 821.100 119.030 ;
        RECT 0.580 84.830 821.100 112.730 ;
        RECT 0.580 66.230 821.100 78.530 ;
        RECT 0.580 47.630 821.100 59.930 ;
        RECT 0.580 29.030 821.100 41.330 ;
        RECT 0.580 0.900 821.100 22.730 ;
  END
END user_project_wrapper
END LIBRARY

