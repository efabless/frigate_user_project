magic
tech sky130A
magscale 1 2
timestamp 1740783570
<< viali >>
rect 2513 37281 2547 37315
rect 13553 37281 13587 37315
rect 34069 37281 34103 37315
rect 39589 37281 39623 37315
rect 3525 37213 3559 37247
rect 5917 37213 5951 37247
rect 7113 37213 7147 37247
rect 7849 37213 7883 37247
rect 8769 37213 8803 37247
rect 11345 37213 11379 37247
rect 12081 37213 12115 37247
rect 14565 37213 14599 37247
rect 15209 37213 15243 37247
rect 18705 37213 18739 37247
rect 19533 37213 19567 37247
rect 20913 37213 20947 37247
rect 21925 37213 21959 37247
rect 22753 37213 22787 37247
rect 26249 37213 26283 37247
rect 28273 37213 28307 37247
rect 29469 37213 29503 37247
rect 31769 37213 31803 37247
rect 32689 37213 32723 37247
rect 33793 37213 33827 37247
rect 36829 37213 36863 37247
rect 37565 37213 37599 37247
rect 39129 37213 39163 37247
rect 40969 37213 41003 37247
rect 41889 37213 41923 37247
rect 43361 37213 43395 37247
rect 46489 37213 46523 37247
rect 48513 37213 48547 37247
rect 52009 37213 52043 37247
rect 52929 37213 52963 37247
rect 53849 37213 53883 37247
rect 56241 37213 56275 37247
rect 58817 37213 58851 37247
rect 16129 37145 16163 37179
rect 23673 37145 23707 37179
rect 27169 37145 27203 37179
rect 44281 37145 44315 37179
rect 47409 37145 47443 37179
rect 49433 37145 49467 37179
rect 54769 37145 54803 37179
rect 57161 37145 57195 37179
rect 59737 37145 59771 37179
rect 7757 36873 7791 36907
rect 11897 36873 11931 36907
rect 15117 36873 15151 36907
rect 19073 36873 19107 36907
rect 22477 36873 22511 36907
rect 26157 36873 26191 36907
rect 33793 36873 33827 36907
rect 37013 36873 37047 36907
rect 40877 36873 40911 36907
rect 48237 36873 48271 36907
rect 51917 36873 51951 36907
rect 55597 36873 55631 36907
rect 4353 36805 4387 36839
rect 9873 36805 9907 36839
rect 17969 36805 18003 36839
rect 24593 36805 24627 36839
rect 5457 36737 5491 36771
rect 7573 36737 7607 36771
rect 10977 36737 11011 36771
rect 11805 36737 11839 36771
rect 12081 36737 12115 36771
rect 14933 36737 14967 36771
rect 18797 36737 18831 36771
rect 19257 36737 19291 36771
rect 22293 36737 22327 36771
rect 25789 36737 25823 36771
rect 25973 36737 26007 36771
rect 29653 36737 29687 36771
rect 29929 36737 29963 36771
rect 33517 36737 33551 36771
rect 33701 36737 33735 36771
rect 33977 36737 34011 36771
rect 35449 36737 35483 36771
rect 37197 36737 37231 36771
rect 40693 36737 40727 36771
rect 44373 36737 44407 36771
rect 44649 36737 44683 36771
rect 48053 36737 48087 36771
rect 50169 36737 50203 36771
rect 51733 36737 51767 36771
rect 55413 36737 55447 36771
rect 58449 36737 58483 36771
rect 59369 36737 59403 36771
rect 11621 36669 11655 36703
rect 30389 36669 30423 36703
rect 35909 36669 35943 36703
rect 45109 36669 45143 36703
rect 50629 36669 50663 36703
rect 59829 36669 59863 36703
rect 29837 36601 29871 36635
rect 44557 36601 44591 36635
rect 58633 36601 58667 36635
rect 22109 11849 22143 11883
rect 26233 11849 26267 11883
rect 28825 11849 28859 11883
rect 29101 11849 29135 11883
rect 23765 11781 23799 11815
rect 26433 11781 26467 11815
rect 30021 11781 30055 11815
rect 30573 11781 30607 11815
rect 33241 11781 33275 11815
rect 22477 11713 22511 11747
rect 23673 11713 23707 11747
rect 24777 11713 24811 11747
rect 25145 11713 25179 11747
rect 26985 11713 27019 11747
rect 27169 11713 27203 11747
rect 27261 11713 27295 11747
rect 28641 11713 28675 11747
rect 28901 11713 28935 11747
rect 29009 11713 29043 11747
rect 29561 11713 29595 11747
rect 30481 11713 30515 11747
rect 30757 11713 30791 11747
rect 33333 11713 33367 11747
rect 33425 11713 33459 11747
rect 23305 11645 23339 11679
rect 28457 11645 28491 11679
rect 29471 11645 29505 11679
rect 33057 11577 33091 11611
rect 22293 11509 22327 11543
rect 22753 11509 22787 11543
rect 23489 11509 23523 11543
rect 25237 11509 25271 11543
rect 26065 11509 26099 11543
rect 26249 11509 26283 11543
rect 26801 11509 26835 11543
rect 29285 11509 29319 11543
rect 30113 11509 30147 11543
rect 30941 11509 30975 11543
rect 33609 11509 33643 11543
rect 22937 11305 22971 11339
rect 25329 11305 25363 11339
rect 26065 11305 26099 11339
rect 28825 11305 28859 11339
rect 31677 11305 31711 11339
rect 33057 11237 33091 11271
rect 23949 11169 23983 11203
rect 24225 11169 24259 11203
rect 24409 11169 24443 11203
rect 25881 11169 25915 11203
rect 26249 11169 26283 11203
rect 26801 11169 26835 11203
rect 30113 11169 30147 11203
rect 32229 11169 32263 11203
rect 33793 11169 33827 11203
rect 34161 11169 34195 11203
rect 34437 11169 34471 11203
rect 21741 11101 21775 11135
rect 22569 11101 22603 11135
rect 24685 11101 24719 11135
rect 24869 11101 24903 11135
rect 24961 11101 24995 11135
rect 26985 11101 27019 11135
rect 27721 11101 27755 11135
rect 28457 11101 28491 11135
rect 29377 11101 29411 11135
rect 31401 11101 31435 11135
rect 33609 11101 33643 11135
rect 33977 11101 34011 11135
rect 34069 11101 34103 11135
rect 34253 11101 34287 11135
rect 34713 11101 34747 11135
rect 34805 11101 34839 11135
rect 21833 11033 21867 11067
rect 22385 11033 22419 11067
rect 23213 11033 23247 11067
rect 23397 11033 23431 11067
rect 24501 11033 24535 11067
rect 27905 11033 27939 11067
rect 29561 11033 29595 11067
rect 30757 11033 30791 11067
rect 34621 11033 34655 11067
rect 34989 11033 35023 11067
rect 22753 10965 22787 10999
rect 25053 10965 25087 10999
rect 27169 10965 27203 10999
rect 24501 10761 24535 10795
rect 27721 10761 27755 10795
rect 33333 10761 33367 10795
rect 20545 10625 20579 10659
rect 21005 10625 21039 10659
rect 21557 10625 21591 10659
rect 21741 10625 21775 10659
rect 22753 10625 22787 10659
rect 22937 10625 22971 10659
rect 23673 10625 23707 10659
rect 24409 10625 24443 10659
rect 25237 10625 25271 10659
rect 26065 10625 26099 10659
rect 26249 10625 26283 10659
rect 26617 10625 26651 10659
rect 28089 10625 28123 10659
rect 32045 10625 32079 10659
rect 34069 10625 34103 10659
rect 21281 10557 21315 10591
rect 22385 10557 22419 10591
rect 24133 10557 24167 10591
rect 26433 10557 26467 10591
rect 27077 10557 27111 10591
rect 28825 10557 28859 10591
rect 29745 10557 29779 10591
rect 30481 10557 30515 10591
rect 30941 10557 30975 10591
rect 32781 10557 32815 10591
rect 33149 10557 33183 10591
rect 34805 10557 34839 10591
rect 35541 10557 35575 10591
rect 21649 10489 21683 10523
rect 23857 10489 23891 10523
rect 30849 10489 30883 10523
rect 33517 10489 33551 10523
rect 34989 10489 35023 10523
rect 20637 10421 20671 10455
rect 20821 10421 20855 10455
rect 21189 10421 21223 10455
rect 21833 10421 21867 10455
rect 23121 10421 23155 10455
rect 24041 10421 24075 10455
rect 24685 10421 24719 10455
rect 25513 10421 25547 10455
rect 26801 10421 26835 10455
rect 27905 10421 27939 10455
rect 28273 10421 28307 10455
rect 29009 10421 29043 10455
rect 29193 10421 29227 10455
rect 29929 10421 29963 10455
rect 31493 10421 31527 10455
rect 32229 10421 32263 10455
rect 34253 10421 34287 10455
rect 26341 10217 26375 10251
rect 27169 10217 27203 10251
rect 20269 10149 20303 10183
rect 33609 10149 33643 10183
rect 21373 10081 21407 10115
rect 22385 10081 22419 10115
rect 22937 10081 22971 10115
rect 23673 10081 23707 10115
rect 26249 10081 26283 10115
rect 28917 10081 28951 10115
rect 29561 10081 29595 10115
rect 19625 10013 19659 10047
rect 19901 10013 19935 10047
rect 20453 10013 20487 10047
rect 20545 10013 20579 10047
rect 22109 10013 22143 10047
rect 23305 10013 23339 10047
rect 24501 10013 24535 10047
rect 26985 10013 27019 10047
rect 27997 10013 28031 10047
rect 28181 10013 28215 10047
rect 29745 10013 29779 10047
rect 31125 10013 31159 10047
rect 31309 10013 31343 10047
rect 31953 10013 31987 10047
rect 32597 10013 32631 10047
rect 33425 10013 33459 10047
rect 34253 10013 34287 10047
rect 34897 10013 34931 10047
rect 36461 10013 36495 10047
rect 36645 10013 36679 10047
rect 37289 10013 37323 10047
rect 23397 9945 23431 9979
rect 23581 9945 23615 9979
rect 19441 9877 19475 9911
rect 19717 9877 19751 9911
rect 20821 9877 20855 9911
rect 21557 9877 21591 9911
rect 23121 9877 23155 9911
rect 23305 9877 23339 9911
rect 24317 9877 24351 9911
rect 25053 9877 25087 9911
rect 25605 9877 25639 9911
rect 27445 9877 27479 9911
rect 28825 9877 28859 9911
rect 30297 9877 30331 9911
rect 30573 9877 30607 9911
rect 32045 9877 32079 9911
rect 32873 9877 32907 9911
rect 34345 9877 34379 9911
rect 35909 9877 35943 9911
rect 34805 9673 34839 9707
rect 20913 9605 20947 9639
rect 27353 9605 27387 9639
rect 19257 9537 19291 9571
rect 22201 9537 22235 9571
rect 22569 9537 22603 9571
rect 24225 9537 24259 9571
rect 25145 9537 25179 9571
rect 25329 9537 25363 9571
rect 26617 9537 26651 9571
rect 26801 9537 26835 9571
rect 27445 9537 27479 9571
rect 27997 9537 28031 9571
rect 28733 9537 28767 9571
rect 29561 9537 29595 9571
rect 33517 9537 33551 9571
rect 35817 9537 35851 9571
rect 37565 9537 37599 9571
rect 37657 9537 37691 9571
rect 37841 9537 37875 9571
rect 19901 9469 19935 9503
rect 20729 9469 20763 9503
rect 21557 9469 21591 9503
rect 22477 9469 22511 9503
rect 23489 9469 23523 9503
rect 25973 9469 26007 9503
rect 28641 9469 28675 9503
rect 30113 9469 30147 9503
rect 30389 9469 30423 9503
rect 31217 9469 31251 9503
rect 31861 9469 31895 9503
rect 34161 9469 34195 9503
rect 35081 9469 35115 9503
rect 35725 9469 35759 9503
rect 36369 9469 36403 9503
rect 37289 9469 37323 9503
rect 38853 9469 38887 9503
rect 20085 9401 20119 9435
rect 21649 9401 21683 9435
rect 27629 9401 27663 9435
rect 36553 9401 36587 9435
rect 37749 9401 37783 9435
rect 18613 9333 18647 9367
rect 19349 9333 19383 9367
rect 22937 9333 22971 9367
rect 23673 9333 23707 9367
rect 24501 9333 24535 9367
rect 25881 9333 25915 9367
rect 29377 9333 29411 9367
rect 30205 9333 30239 9367
rect 31033 9333 31067 9367
rect 31769 9333 31803 9367
rect 32505 9333 32539 9367
rect 34069 9333 34103 9367
rect 34897 9333 34931 9367
rect 36737 9333 36771 9367
rect 38025 9333 38059 9367
rect 38209 9333 38243 9367
rect 11713 9129 11747 9163
rect 19257 9129 19291 9163
rect 21281 9129 21315 9163
rect 22201 9129 22235 9163
rect 28641 9129 28675 9163
rect 29653 9129 29687 9163
rect 32229 9129 32263 9163
rect 17141 9061 17175 9095
rect 20361 9061 20395 9095
rect 25513 9061 25547 9095
rect 35449 9061 35483 9095
rect 17693 8993 17727 9027
rect 18521 8993 18555 9027
rect 21097 8993 21131 9027
rect 23581 8993 23615 9027
rect 25697 8993 25731 9027
rect 27077 8993 27111 9027
rect 27997 8993 28031 9027
rect 29469 8993 29503 9027
rect 32781 8993 32815 9027
rect 34621 8993 34655 9027
rect 36829 8993 36863 9027
rect 40049 8993 40083 9027
rect 11621 8925 11655 8959
rect 16497 8925 16531 8959
rect 18613 8925 18647 8959
rect 19349 8925 19383 8959
rect 20269 8925 20303 8959
rect 20453 8925 20487 8959
rect 21833 8925 21867 8959
rect 22017 8925 22051 8959
rect 22201 8925 22235 8959
rect 22569 8925 22603 8959
rect 22661 8925 22695 8959
rect 22753 8925 22787 8959
rect 22937 8925 22971 8959
rect 23765 8925 23799 8959
rect 24685 8925 24719 8959
rect 24777 8925 24811 8959
rect 25329 8925 25363 8959
rect 26433 8925 26467 8959
rect 27629 8925 27663 8959
rect 28917 8925 28951 8959
rect 30205 8925 30239 8959
rect 31309 8925 31343 8959
rect 31401 8925 31435 8959
rect 33977 8925 34011 8959
rect 34805 8925 34839 8959
rect 34897 8925 34931 8959
rect 35173 8925 35207 8959
rect 35265 8925 35299 8959
rect 35817 8925 35851 8959
rect 36001 8925 36035 8959
rect 36645 8925 36679 8959
rect 37381 8925 37415 8959
rect 38209 8925 38243 8959
rect 38853 8925 38887 8959
rect 39497 8925 39531 8959
rect 20545 8857 20579 8891
rect 23029 8857 23063 8891
rect 24501 8857 24535 8891
rect 30941 8857 30975 8891
rect 31677 8857 31711 8891
rect 31769 8857 31803 8891
rect 35081 8857 35115 8891
rect 15945 8789 15979 8823
rect 17877 8789 17911 8823
rect 19993 8789 20027 8823
rect 22293 8789 22327 8823
rect 24409 8789 24443 8823
rect 25145 8789 25179 8823
rect 26249 8789 26283 8823
rect 26985 8789 27019 8823
rect 31125 8789 31159 8823
rect 33333 8789 33367 8823
rect 34069 8789 34103 8823
rect 35633 8789 35667 8823
rect 36093 8789 36127 8823
rect 37565 8789 37599 8823
rect 39405 8789 39439 8823
rect 18889 8585 18923 8619
rect 21833 8585 21867 8619
rect 32663 8585 32697 8619
rect 18153 8517 18187 8551
rect 24225 8517 24259 8551
rect 25973 8517 26007 8551
rect 27997 8517 28031 8551
rect 31677 8517 31711 8551
rect 32873 8517 32907 8551
rect 38209 8517 38243 8551
rect 17785 8449 17819 8483
rect 19625 8449 19659 8483
rect 21005 8449 21039 8483
rect 22017 8449 22051 8483
rect 22569 8449 22603 8483
rect 22845 8449 22879 8483
rect 23765 8449 23799 8483
rect 26801 8449 26835 8483
rect 26985 8449 27019 8483
rect 27077 8449 27111 8483
rect 27905 8449 27939 8483
rect 28089 8449 28123 8483
rect 28733 8449 28767 8483
rect 29469 8449 29503 8483
rect 33609 8449 33643 8483
rect 34897 8449 34931 8483
rect 39773 8449 39807 8483
rect 16037 8381 16071 8415
rect 16681 8381 16715 8415
rect 17325 8381 17359 8415
rect 18337 8381 18371 8415
rect 20269 8381 20303 8415
rect 21189 8381 21223 8415
rect 23213 8381 23247 8415
rect 23949 8381 23983 8415
rect 26617 8381 26651 8415
rect 27721 8381 27755 8415
rect 29653 8381 29687 8415
rect 29929 8381 29963 8415
rect 32321 8381 32355 8415
rect 33057 8381 33091 8415
rect 34069 8381 34103 8415
rect 34621 8381 34655 8415
rect 35173 8381 35207 8415
rect 36921 8381 36955 8415
rect 37565 8381 37599 8415
rect 38853 8381 38887 8415
rect 38945 8381 38979 8415
rect 39957 8381 39991 8415
rect 16773 8313 16807 8347
rect 20453 8313 20487 8347
rect 26801 8313 26835 8347
rect 28181 8313 28215 8347
rect 37013 8313 37047 8347
rect 39221 8313 39255 8347
rect 40601 8313 40635 8347
rect 18981 8245 19015 8279
rect 19717 8245 19751 8279
rect 22937 8245 22971 8279
rect 26065 8245 26099 8279
rect 28917 8245 28951 8279
rect 31769 8245 31803 8279
rect 32505 8245 32539 8279
rect 32689 8245 32723 8279
rect 19993 8041 20027 8075
rect 20177 8041 20211 8075
rect 20545 8041 20579 8075
rect 21281 8041 21315 8075
rect 24501 8041 24535 8075
rect 25329 8041 25363 8075
rect 27353 8041 27387 8075
rect 29561 8041 29595 8075
rect 35449 8041 35483 8075
rect 15669 7973 15703 8007
rect 17049 7973 17083 8007
rect 28181 7973 28215 8007
rect 34253 7973 34287 8007
rect 16405 7905 16439 7939
rect 17877 7905 17911 7939
rect 18705 7905 18739 7939
rect 21373 7905 21407 7939
rect 22017 7905 22051 7939
rect 22109 7905 22143 7939
rect 24133 7905 24167 7939
rect 25145 7905 25179 7939
rect 26801 7905 26835 7939
rect 28825 7905 28859 7939
rect 30297 7905 30331 7939
rect 32137 7905 32171 7939
rect 34805 7905 34839 7939
rect 36001 7905 36035 7939
rect 38025 7905 38059 7939
rect 38117 7905 38151 7939
rect 39589 7905 39623 7939
rect 41429 7905 41463 7939
rect 14105 7837 14139 7871
rect 15025 7837 15059 7871
rect 15209 7837 15243 7871
rect 15301 7837 15335 7871
rect 16221 7837 16255 7871
rect 17141 7837 17175 7871
rect 19257 7837 19291 7871
rect 19441 7837 19475 7871
rect 20177 7837 20211 7871
rect 20269 7837 20303 7871
rect 20729 7837 20763 7871
rect 24225 7837 24259 7871
rect 24409 7837 24443 7871
rect 25513 7837 25547 7871
rect 25605 7837 25639 7871
rect 25789 7837 25823 7871
rect 25881 7837 25915 7871
rect 25973 7837 26007 7871
rect 27445 7837 27479 7871
rect 28917 7837 28951 7871
rect 30481 7837 30515 7871
rect 30665 7837 30699 7871
rect 30849 7837 30883 7871
rect 31493 7837 31527 7871
rect 34437 7837 34471 7871
rect 34713 7837 34747 7871
rect 35633 7837 35667 7871
rect 35817 7837 35851 7871
rect 38853 7837 38887 7871
rect 40233 7837 40267 7871
rect 17785 7769 17819 7803
rect 22385 7769 22419 7803
rect 28089 7769 28123 7803
rect 32413 7769 32447 7803
rect 34161 7769 34195 7803
rect 35725 7769 35759 7803
rect 36277 7769 36311 7803
rect 41613 7769 41647 7803
rect 14749 7701 14783 7735
rect 15117 7701 15151 7735
rect 15485 7701 15519 7735
rect 18521 7701 18555 7735
rect 24317 7701 24351 7735
rect 26617 7701 26651 7735
rect 29653 7701 29687 7735
rect 30941 7701 30975 7735
rect 34621 7701 34655 7735
rect 38761 7701 38795 7735
rect 39497 7701 39531 7735
rect 40785 7701 40819 7735
rect 41889 7701 41923 7735
rect 11897 7497 11931 7531
rect 15945 7497 15979 7531
rect 17601 7497 17635 7531
rect 18889 7497 18923 7531
rect 21097 7497 21131 7531
rect 21189 7497 21223 7531
rect 22569 7497 22603 7531
rect 24961 7497 24995 7531
rect 27721 7497 27755 7531
rect 32229 7497 32263 7531
rect 33977 7497 34011 7531
rect 34897 7497 34931 7531
rect 35909 7497 35943 7531
rect 42073 7497 42107 7531
rect 25329 7429 25363 7463
rect 27077 7429 27111 7463
rect 27445 7429 27479 7463
rect 28825 7429 28859 7463
rect 30021 7429 30055 7463
rect 31769 7429 31803 7463
rect 35081 7429 35115 7463
rect 35449 7429 35483 7463
rect 13737 7361 13771 7395
rect 13829 7361 13863 7395
rect 14105 7361 14139 7395
rect 14381 7361 14415 7395
rect 14473 7361 14507 7395
rect 14565 7361 14599 7395
rect 16589 7361 16623 7395
rect 17417 7361 17451 7395
rect 17785 7361 17819 7395
rect 17877 7361 17911 7395
rect 18153 7361 18187 7395
rect 20453 7361 20487 7395
rect 20601 7361 20635 7395
rect 20729 7361 20763 7395
rect 20821 7361 20855 7395
rect 20959 7361 20993 7395
rect 21833 7361 21867 7395
rect 22017 7361 22051 7395
rect 25053 7361 25087 7395
rect 27169 7361 27203 7395
rect 27353 7361 27387 7395
rect 27537 7361 27571 7395
rect 29745 7361 29779 7395
rect 31861 7361 31895 7395
rect 31953 7361 31987 7395
rect 32137 7361 32171 7395
rect 32505 7361 32539 7395
rect 33057 7361 33091 7395
rect 33241 7361 33275 7395
rect 34621 7361 34655 7395
rect 34805 7361 34839 7395
rect 35173 7361 35207 7395
rect 35265 7361 35299 7395
rect 35541 7361 35575 7395
rect 35633 7361 35667 7395
rect 36553 7361 36587 7395
rect 37289 7361 37323 7395
rect 38301 7361 38335 7395
rect 40233 7361 40267 7395
rect 41153 7361 41187 7395
rect 42625 7361 42659 7395
rect 11253 7293 11287 7327
rect 13369 7293 13403 7327
rect 15301 7293 15335 7327
rect 16037 7293 16071 7327
rect 18337 7293 18371 7327
rect 18981 7293 19015 7327
rect 19717 7293 19751 7327
rect 23213 7293 23247 7327
rect 23765 7293 23799 7327
rect 24317 7293 24351 7327
rect 28273 7293 28307 7327
rect 28917 7293 28951 7327
rect 29561 7293 29595 7327
rect 32413 7293 32447 7327
rect 32781 7293 32815 7327
rect 32873 7293 32907 7327
rect 33425 7293 33459 7327
rect 34069 7293 34103 7327
rect 37381 7293 37415 7327
rect 38853 7293 38887 7327
rect 39497 7293 39531 7327
rect 41429 7293 41463 7327
rect 16773 7225 16807 7259
rect 32137 7225 32171 7259
rect 39681 7225 39715 7259
rect 12817 7157 12851 7191
rect 13553 7157 13587 7191
rect 15209 7157 15243 7191
rect 18061 7157 18095 7191
rect 19625 7157 19659 7191
rect 20361 7157 20395 7191
rect 33149 7157 33183 7191
rect 35081 7157 35115 7191
rect 35817 7157 35851 7191
rect 36645 7157 36679 7191
rect 38025 7157 38059 7191
rect 38945 7157 38979 7191
rect 40601 7157 40635 7191
rect 41981 7157 42015 7191
rect 16681 6953 16715 6987
rect 18981 6953 19015 6987
rect 21937 6953 21971 6987
rect 22477 6953 22511 6987
rect 25881 6953 25915 6987
rect 26966 6953 27000 6987
rect 37736 6953 37770 6987
rect 25329 6885 25363 6919
rect 30297 6885 30331 6919
rect 11989 6817 12023 6851
rect 13369 6817 13403 6851
rect 14841 6817 14875 6851
rect 17417 6817 17451 6851
rect 22201 6817 22235 6851
rect 23673 6817 23707 6851
rect 24593 6817 24627 6851
rect 26525 6817 26559 6851
rect 26709 6817 26743 6851
rect 28733 6817 28767 6851
rect 28917 6817 28951 6851
rect 29561 6817 29595 6851
rect 29745 6817 29779 6851
rect 31401 6817 31435 6851
rect 31953 6817 31987 6851
rect 33241 6817 33275 6851
rect 33977 6817 34011 6851
rect 36553 6817 36587 6851
rect 37289 6817 37323 6851
rect 37473 6817 37507 6851
rect 42257 6817 42291 6851
rect 11161 6749 11195 6783
rect 12725 6749 12759 6783
rect 14105 6749 14139 6783
rect 15025 6749 15059 6783
rect 15209 6749 15243 6783
rect 15853 6749 15887 6783
rect 16129 6749 16163 6783
rect 16865 6749 16899 6783
rect 17509 6749 17543 6783
rect 18245 6749 18279 6783
rect 18797 6749 18831 6783
rect 19533 6749 19567 6783
rect 23489 6749 23523 6783
rect 25513 6749 25547 6783
rect 25697 6749 25731 6783
rect 25973 6749 26007 6783
rect 31309 6749 31343 6783
rect 32597 6749 32631 6783
rect 33333 6749 33367 6783
rect 34621 6749 34655 6783
rect 35357 6749 35391 6783
rect 35817 6749 35851 6783
rect 36737 6749 36771 6783
rect 40141 6749 40175 6783
rect 40785 6749 40819 6783
rect 42073 6749 42107 6783
rect 20177 6681 20211 6715
rect 22461 6681 22495 6715
rect 22661 6681 22695 6715
rect 24225 6681 24259 6715
rect 25145 6681 25179 6715
rect 34069 6681 34103 6715
rect 35909 6681 35943 6715
rect 39497 6681 39531 6715
rect 10057 6613 10091 6647
rect 11805 6613 11839 6647
rect 12633 6613 12667 6647
rect 13461 6613 13495 6647
rect 14197 6613 14231 6647
rect 15117 6613 15151 6647
rect 15301 6613 15335 6647
rect 18153 6613 18187 6647
rect 22293 6613 22327 6647
rect 22845 6613 22879 6647
rect 25605 6613 25639 6647
rect 30665 6613 30699 6647
rect 34805 6613 34839 6647
rect 35725 6613 35759 6647
rect 39589 6613 39623 6647
rect 41429 6613 41463 6647
rect 41521 6613 41555 6647
rect 42901 6613 42935 6647
rect 10885 6409 10919 6443
rect 13737 6409 13771 6443
rect 17417 6409 17451 6443
rect 23213 6409 23247 6443
rect 23397 6409 23431 6443
rect 24409 6409 24443 6443
rect 26893 6409 26927 6443
rect 27261 6409 27295 6443
rect 35633 6409 35667 6443
rect 10793 6341 10827 6375
rect 12265 6341 12299 6375
rect 21281 6341 21315 6375
rect 22201 6341 22235 6375
rect 22401 6341 22435 6375
rect 23029 6341 23063 6375
rect 26617 6341 26651 6375
rect 27353 6341 27387 6375
rect 35081 6341 35115 6375
rect 38025 6341 38059 6375
rect 38485 6341 38519 6375
rect 40233 6341 40267 6375
rect 9781 6273 9815 6307
rect 11529 6273 11563 6307
rect 12449 6273 12483 6307
rect 12817 6273 12851 6307
rect 13185 6273 13219 6307
rect 14657 6273 14691 6307
rect 15945 6273 15979 6307
rect 16681 6273 16715 6307
rect 16865 6273 16899 6307
rect 19809 6273 19843 6307
rect 21741 6273 21775 6307
rect 23305 6273 23339 6307
rect 23857 6273 23891 6307
rect 26065 6273 26099 6307
rect 27905 6273 27939 6307
rect 29837 6273 29871 6307
rect 30021 6273 30055 6307
rect 30113 6273 30147 6307
rect 30941 6273 30975 6307
rect 31861 6273 31895 6307
rect 32597 6273 32631 6307
rect 35173 6273 35207 6307
rect 35265 6273 35299 6307
rect 35449 6273 35483 6307
rect 36277 6273 36311 6307
rect 37381 6273 37415 6307
rect 41797 6273 41831 6307
rect 42717 6273 42751 6307
rect 42809 6273 42843 6307
rect 42993 6273 43027 6307
rect 44097 6273 44131 6307
rect 9597 6205 9631 6239
rect 10241 6205 10275 6239
rect 11621 6205 11655 6239
rect 13829 6205 13863 6239
rect 14381 6205 14415 6239
rect 15209 6205 15243 6239
rect 17693 6205 17727 6239
rect 18245 6205 18279 6239
rect 19073 6205 19107 6239
rect 19901 6205 19935 6239
rect 20637 6205 20671 6239
rect 21833 6205 21867 6239
rect 21925 6205 21959 6239
rect 24501 6205 24535 6239
rect 25329 6205 25363 6239
rect 27445 6205 27479 6239
rect 29653 6205 29687 6239
rect 29929 6205 29963 6239
rect 30297 6205 30331 6239
rect 31125 6205 31159 6239
rect 31769 6205 31803 6239
rect 32689 6205 32723 6239
rect 33057 6205 33091 6239
rect 33333 6205 33367 6239
rect 37289 6205 37323 6239
rect 38209 6205 38243 6239
rect 40601 6205 40635 6239
rect 41245 6205 41279 6239
rect 42625 6205 42659 6239
rect 43177 6205 43211 6239
rect 43361 6205 43395 6239
rect 9965 6137 9999 6171
rect 19165 6137 19199 6171
rect 20545 6137 20579 6171
rect 22569 6137 22603 6171
rect 23581 6137 23615 6171
rect 32505 6137 32539 6171
rect 35725 6137 35759 6171
rect 44005 6137 44039 6171
rect 9045 6069 9079 6103
rect 15301 6069 15335 6103
rect 16037 6069 16071 6103
rect 18429 6069 18463 6103
rect 21373 6069 21407 6103
rect 22345 6069 22379 6103
rect 25145 6069 25179 6103
rect 25881 6069 25915 6103
rect 30389 6069 30423 6103
rect 36645 6069 36679 6103
rect 41153 6069 41187 6103
rect 41981 6069 42015 6103
rect 44741 6069 44775 6103
rect 8585 5865 8619 5899
rect 12725 5865 12759 5899
rect 14841 5865 14875 5899
rect 18521 5865 18555 5899
rect 20177 5865 20211 5899
rect 20361 5865 20395 5899
rect 21465 5865 21499 5899
rect 24409 5865 24443 5899
rect 26617 5865 26651 5899
rect 30481 5865 30515 5899
rect 31309 5865 31343 5899
rect 32505 5865 32539 5899
rect 33885 5865 33919 5899
rect 42993 5865 43027 5899
rect 15577 5797 15611 5831
rect 16313 5797 16347 5831
rect 20729 5797 20763 5831
rect 30297 5797 30331 5831
rect 34437 5797 34471 5831
rect 34805 5797 34839 5831
rect 10609 5729 10643 5763
rect 11253 5729 11287 5763
rect 11897 5729 11931 5763
rect 15669 5729 15703 5763
rect 16957 5729 16991 5763
rect 19165 5729 19199 5763
rect 19441 5729 19475 5763
rect 22937 5729 22971 5763
rect 23673 5729 23707 5763
rect 24501 5729 24535 5763
rect 25329 5729 25363 5763
rect 25513 5729 25547 5763
rect 25789 5729 25823 5763
rect 25973 5729 26007 5763
rect 27353 5729 27387 5763
rect 28825 5729 28859 5763
rect 29561 5729 29595 5763
rect 29653 5729 29687 5763
rect 30941 5729 30975 5763
rect 31125 5729 31159 5763
rect 31953 5729 31987 5763
rect 36921 5729 36955 5763
rect 39313 5729 39347 5763
rect 42073 5729 42107 5763
rect 44465 5729 44499 5763
rect 45937 5729 45971 5763
rect 8033 5661 8067 5695
rect 9045 5661 9079 5695
rect 10149 5661 10183 5695
rect 10333 5661 10367 5695
rect 10425 5661 10459 5695
rect 11989 5661 12023 5695
rect 13277 5661 13311 5695
rect 14105 5661 14139 5695
rect 14289 5661 14323 5695
rect 15117 5661 15151 5695
rect 15209 5661 15243 5695
rect 15393 5661 15427 5695
rect 17693 5661 17727 5695
rect 17877 5661 17911 5695
rect 20913 5661 20947 5695
rect 22201 5661 22235 5695
rect 22385 5661 22419 5695
rect 23857 5661 23891 5695
rect 25605 5661 25639 5695
rect 25697 5661 25731 5695
rect 28089 5661 28123 5695
rect 30849 5661 30883 5695
rect 31493 5661 31527 5695
rect 31769 5661 31803 5695
rect 32597 5661 32631 5695
rect 34437 5661 34471 5695
rect 34529 5661 34563 5695
rect 35081 5661 35115 5695
rect 35173 5661 35207 5695
rect 35265 5661 35299 5695
rect 35449 5661 35483 5695
rect 35725 5661 35759 5695
rect 38945 5661 38979 5695
rect 39865 5661 39899 5695
rect 40509 5661 40543 5695
rect 41429 5661 41463 5695
rect 41521 5661 41555 5695
rect 42901 5661 42935 5695
rect 43637 5661 43671 5695
rect 44373 5661 44407 5695
rect 45109 5661 45143 5695
rect 9689 5593 9723 5627
rect 11161 5593 11195 5627
rect 13461 5593 13495 5627
rect 23029 5593 23063 5627
rect 28181 5593 28215 5627
rect 31677 5593 31711 5627
rect 34713 5593 34747 5627
rect 36369 5593 36403 5627
rect 37105 5593 37139 5627
rect 42257 5593 42291 5627
rect 9965 5525 9999 5559
rect 12633 5525 12667 5559
rect 16405 5525 16439 5559
rect 17141 5525 17175 5559
rect 18613 5525 18647 5559
rect 19993 5525 20027 5559
rect 20361 5525 20395 5559
rect 21557 5525 21591 5559
rect 25145 5525 25179 5559
rect 26709 5525 26743 5559
rect 27445 5525 27479 5559
rect 28917 5525 28951 5559
rect 36277 5525 36311 5559
rect 38393 5525 38427 5559
rect 39037 5525 39071 5559
rect 39957 5525 39991 5559
rect 40785 5525 40819 5559
rect 43729 5525 43763 5559
rect 46581 5525 46615 5559
rect 8401 5321 8435 5355
rect 9137 5321 9171 5355
rect 11529 5321 11563 5355
rect 12265 5321 12299 5355
rect 12633 5321 12667 5355
rect 15209 5321 15243 5355
rect 16129 5321 16163 5355
rect 20821 5321 20855 5355
rect 21281 5321 21315 5355
rect 21833 5321 21867 5355
rect 22569 5321 22603 5355
rect 24041 5321 24075 5355
rect 25513 5321 25547 5355
rect 29561 5321 29595 5355
rect 30297 5321 30331 5355
rect 32781 5321 32815 5355
rect 33609 5321 33643 5355
rect 35173 5321 35207 5355
rect 36553 5321 36587 5355
rect 41521 5321 41555 5355
rect 9965 5253 9999 5287
rect 13553 5253 13587 5287
rect 16681 5253 16715 5287
rect 19257 5253 19291 5287
rect 22753 5253 22787 5287
rect 30849 5253 30883 5287
rect 33241 5253 33275 5287
rect 36645 5253 36679 5287
rect 7481 5185 7515 5219
rect 8585 5185 8619 5219
rect 9781 5185 9815 5219
rect 11713 5185 11747 5219
rect 12449 5185 12483 5219
rect 13737 5185 13771 5219
rect 16405 5185 16439 5219
rect 17693 5185 17727 5219
rect 21189 5185 21223 5219
rect 21649 5185 21683 5219
rect 21925 5185 21959 5219
rect 24777 5185 24811 5219
rect 24961 5185 24995 5219
rect 26433 5185 26467 5219
rect 27905 5185 27939 5219
rect 32597 5185 32631 5219
rect 32873 5185 32907 5219
rect 33057 5185 33091 5219
rect 33333 5185 33367 5219
rect 33425 5185 33459 5219
rect 35081 5185 35115 5219
rect 35817 5185 35851 5219
rect 35909 5185 35943 5219
rect 36093 5185 36127 5219
rect 36185 5185 36219 5219
rect 36277 5185 36311 5219
rect 38209 5185 38243 5219
rect 38393 5185 38427 5219
rect 39497 5185 39531 5219
rect 40877 5185 40911 5219
rect 42349 5185 42383 5219
rect 44005 5185 44039 5219
rect 45477 5185 45511 5219
rect 47041 5185 47075 5219
rect 7849 5117 7883 5151
rect 10517 5117 10551 5151
rect 10885 5117 10919 5151
rect 13001 5117 13035 5151
rect 14473 5117 14507 5151
rect 14657 5117 14691 5151
rect 15945 5117 15979 5151
rect 16589 5117 16623 5151
rect 16773 5117 16807 5151
rect 17785 5117 17819 5151
rect 17877 5117 17911 5151
rect 17969 5117 18003 5151
rect 18337 5117 18371 5151
rect 18981 5117 19015 5151
rect 20729 5117 20763 5151
rect 21373 5117 21407 5151
rect 25697 5117 25731 5151
rect 27169 5117 27203 5151
rect 28273 5117 28307 5151
rect 28917 5117 28951 5151
rect 29745 5117 29779 5151
rect 30573 5117 30607 5151
rect 33701 5117 33735 5151
rect 37289 5117 37323 5151
rect 37933 5117 37967 5151
rect 38669 5117 38703 5151
rect 39313 5117 39347 5151
rect 40049 5117 40083 5151
rect 40693 5117 40727 5151
rect 41613 5117 41647 5151
rect 42901 5117 42935 5151
rect 44097 5117 44131 5151
rect 45569 5117 45603 5151
rect 46949 5117 46983 5151
rect 77493 5117 77527 5151
rect 9229 5049 9263 5083
rect 15301 5049 15335 5083
rect 26249 5049 26283 5083
rect 34437 5049 34471 5083
rect 38577 5049 38611 5083
rect 40141 5049 40175 5083
rect 44833 5049 44867 5083
rect 46213 5049 46247 5083
rect 7665 4981 7699 5015
rect 10701 4981 10735 5015
rect 14289 4981 14323 5015
rect 16221 4981 16255 5015
rect 16589 4981 16623 5015
rect 17417 4981 17451 5015
rect 18153 4981 18187 5015
rect 18889 4981 18923 5015
rect 24593 4981 24627 5015
rect 26985 4981 27019 5015
rect 27721 4981 27755 5015
rect 28089 4981 28123 5015
rect 28825 4981 28859 5015
rect 34345 4981 34379 5015
rect 37381 4981 37415 5015
rect 42257 4981 42291 5015
rect 43361 4981 43395 5015
rect 44741 4981 44775 5015
rect 46305 4981 46339 5015
rect 47685 4981 47719 5015
rect 76941 4981 76975 5015
rect 8953 4777 8987 4811
rect 10241 4777 10275 4811
rect 11897 4777 11931 4811
rect 16497 4777 16531 4811
rect 19073 4777 19107 4811
rect 23397 4777 23431 4811
rect 24317 4777 24351 4811
rect 27905 4777 27939 4811
rect 29653 4777 29687 4811
rect 31401 4777 31435 4811
rect 32689 4777 32723 4811
rect 32873 4777 32907 4811
rect 33333 4777 33367 4811
rect 37105 4777 37139 4811
rect 41429 4777 41463 4811
rect 42809 4777 42843 4811
rect 43545 4777 43579 4811
rect 45017 4777 45051 4811
rect 46673 4777 46707 4811
rect 76941 4777 76975 4811
rect 9689 4709 9723 4743
rect 12633 4709 12667 4743
rect 14105 4709 14139 4743
rect 17233 4709 17267 4743
rect 21833 4709 21867 4743
rect 26249 4709 26283 4743
rect 37013 4709 37047 4743
rect 44281 4709 44315 4743
rect 8309 4641 8343 4675
rect 13369 4641 13403 4675
rect 13553 4641 13587 4675
rect 15853 4641 15887 4675
rect 16589 4641 16623 4675
rect 19717 4641 19751 4675
rect 20545 4641 20579 4675
rect 21097 4641 21131 4675
rect 22569 4641 22603 4675
rect 23949 4641 23983 4675
rect 24777 4641 24811 4675
rect 24961 4641 24995 4675
rect 26433 4641 26467 4675
rect 28365 4641 28399 4675
rect 28457 4641 28491 4675
rect 28917 4641 28951 4675
rect 30757 4641 30791 4675
rect 31861 4641 31895 4675
rect 31953 4641 31987 4675
rect 32597 4641 32631 4675
rect 35633 4641 35667 4675
rect 36461 4641 36495 4675
rect 37749 4641 37783 4675
rect 38209 4641 38243 4675
rect 40877 4641 40911 4675
rect 44833 4641 44867 4675
rect 45937 4641 45971 4675
rect 47225 4641 47259 4675
rect 48881 4641 48915 4675
rect 6745 4573 6779 4607
rect 7481 4573 7515 4607
rect 7665 4573 7699 4607
rect 9137 4573 9171 4607
rect 10609 4573 10643 4607
rect 11161 4573 11195 4607
rect 11345 4573 11379 4607
rect 11989 4573 12023 4607
rect 12817 4573 12851 4607
rect 14197 4573 14231 4607
rect 15117 4573 15151 4607
rect 17417 4573 17451 4607
rect 21281 4573 21315 4607
rect 21925 4573 21959 4607
rect 22661 4573 22695 4607
rect 23765 4573 23799 4607
rect 23857 4573 23891 4607
rect 24685 4573 24719 4607
rect 25697 4573 25731 4607
rect 27721 4573 27755 4607
rect 30297 4573 30331 4607
rect 32689 4573 32723 4607
rect 33977 4573 34011 4607
rect 34161 4573 34195 4607
rect 34897 4573 34931 4607
rect 37933 4573 37967 4607
rect 40233 4573 40267 4607
rect 40325 4573 40359 4607
rect 40601 4573 40635 4607
rect 42257 4573 42291 4607
rect 43453 4573 43487 4607
rect 44189 4573 44223 4607
rect 45569 4573 45603 4607
rect 47409 4573 47443 4607
rect 48789 4573 48823 4607
rect 77585 4573 77619 4607
rect 10333 4505 10367 4539
rect 15761 4505 15795 4539
rect 18061 4505 18095 4539
rect 19441 4505 19475 4539
rect 19533 4505 19567 4539
rect 26985 4505 27019 4539
rect 31309 4505 31343 4539
rect 31769 4505 31803 4539
rect 32229 4505 32263 4539
rect 32965 4505 32999 4539
rect 33149 4505 33183 4539
rect 34713 4505 34747 4539
rect 35449 4505 35483 4539
rect 39957 4505 39991 4539
rect 40417 4505 40451 4539
rect 48053 4505 48087 4539
rect 6101 4437 6135 4471
rect 6837 4437 6871 4471
rect 8217 4437 8251 4471
rect 14841 4437 14875 4471
rect 17969 4437 18003 4471
rect 23305 4437 23339 4471
rect 27077 4437 27111 4471
rect 28273 4437 28307 4471
rect 29561 4437 29595 4471
rect 36277 4437 36311 4471
rect 37473 4437 37507 4471
rect 37565 4437 37599 4471
rect 40049 4437 40083 4471
rect 41705 4437 41739 4471
rect 46581 4437 46615 4471
rect 48145 4437 48179 4471
rect 49525 4437 49559 4471
rect 7113 4233 7147 4267
rect 20085 4233 20119 4267
rect 20821 4233 20855 4267
rect 22911 4233 22945 4267
rect 23949 4233 23983 4267
rect 36737 4233 36771 4267
rect 43729 4233 43763 4267
rect 47133 4233 47167 4267
rect 48329 4233 48363 4267
rect 49157 4233 49191 4267
rect 12541 4165 12575 4199
rect 13369 4165 13403 4199
rect 17417 4165 17451 4199
rect 19809 4165 19843 4199
rect 23121 4165 23155 4199
rect 27905 4165 27939 4199
rect 6377 4097 6411 4131
rect 6469 4097 6503 4131
rect 7573 4097 7607 4131
rect 7757 4097 7791 4131
rect 7849 4097 7883 4131
rect 8033 4097 8067 4131
rect 10149 4097 10183 4131
rect 10793 4097 10827 4131
rect 10977 4097 11011 4131
rect 11529 4097 11563 4131
rect 12265 4097 12299 4131
rect 12633 4097 12667 4131
rect 12725 4097 12759 4131
rect 14657 4097 14691 4131
rect 17601 4097 17635 4131
rect 17785 4097 17819 4131
rect 19901 4097 19935 4131
rect 21281 4097 21315 4131
rect 23397 4097 23431 4131
rect 23489 4097 23523 4131
rect 23765 4097 23799 4131
rect 23949 4097 23983 4131
rect 24225 4097 24259 4131
rect 26341 4097 26375 4131
rect 28089 4097 28123 4131
rect 28181 4097 28215 4131
rect 28641 4097 28675 4131
rect 30297 4097 30331 4131
rect 30849 4097 30883 4131
rect 31493 4097 31527 4131
rect 33057 4097 33091 4131
rect 33241 4097 33275 4131
rect 33977 4097 34011 4131
rect 34069 4097 34103 4131
rect 36277 4097 36311 4131
rect 36829 4097 36863 4131
rect 38025 4097 38059 4131
rect 38485 4097 38519 4131
rect 38577 4097 38611 4131
rect 40417 4097 40451 4131
rect 40509 4097 40543 4131
rect 41061 4097 41095 4131
rect 42533 4097 42567 4131
rect 42993 4097 43027 4131
rect 46397 4097 46431 4131
rect 46949 4097 46983 4131
rect 48053 4097 48087 4131
rect 48145 4097 48179 4131
rect 48513 4097 48547 4131
rect 74733 4097 74767 4131
rect 76205 4097 76239 4131
rect 5733 4029 5767 4063
rect 8769 4029 8803 4063
rect 9321 4029 9355 4063
rect 9505 4029 9539 4063
rect 10057 4029 10091 4063
rect 11621 4029 11655 4063
rect 14381 4029 14415 4063
rect 15117 4029 15151 4063
rect 15945 4029 15979 4063
rect 16865 4029 16899 4063
rect 20269 4029 20303 4063
rect 21373 4029 21407 4063
rect 21557 4029 21591 4063
rect 22017 4029 22051 4063
rect 22569 4029 22603 4063
rect 24501 4029 24535 4063
rect 26249 4029 26283 4063
rect 26893 4029 26927 4063
rect 29101 4029 29135 4063
rect 30389 4029 30423 4063
rect 30481 4029 30515 4063
rect 31953 4029 31987 4063
rect 33425 4029 33459 4063
rect 35265 4029 35299 4063
rect 35725 4029 35759 4063
rect 36921 4029 36955 4063
rect 37749 4029 37783 4063
rect 39037 4029 39071 4063
rect 40601 4029 40635 4063
rect 41153 4029 41187 4063
rect 41797 4029 41831 4063
rect 42901 4029 42935 4063
rect 43453 4029 43487 4063
rect 43637 4029 43671 4063
rect 44189 4029 44223 4063
rect 44741 4029 44775 4063
rect 45569 4029 45603 4063
rect 45661 4029 45695 4063
rect 46305 4029 46339 4063
rect 47777 4029 47811 4063
rect 49249 4029 49283 4063
rect 52193 4029 52227 4063
rect 53849 4029 53883 4063
rect 65533 4029 65567 4063
rect 67649 4029 67683 4063
rect 69305 4029 69339 4063
rect 71513 4029 71547 4063
rect 75929 4029 75963 4063
rect 77033 4029 77067 4063
rect 17969 3961 18003 3995
rect 18521 3961 18555 3995
rect 22753 3961 22787 3995
rect 28365 3961 28399 3995
rect 33241 3961 33275 3995
rect 44097 3961 44131 3995
rect 47869 3961 47903 3995
rect 7389 3893 7423 3927
rect 8585 3893 8619 3927
rect 15761 3893 15795 3927
rect 16497 3893 16531 3927
rect 17601 3893 17635 3927
rect 20913 3893 20947 3927
rect 21833 3893 21867 3927
rect 22937 3893 22971 3927
rect 27905 3893 27939 3927
rect 29929 3893 29963 3927
rect 31401 3893 31435 3927
rect 36369 3893 36403 3927
rect 38301 3893 38335 3927
rect 40049 3893 40083 3927
rect 40877 3893 40911 3927
rect 41889 3893 41923 3927
rect 42717 3893 42751 3927
rect 44925 3893 44959 3927
rect 49893 3893 49927 3927
rect 52745 3893 52779 3927
rect 54401 3893 54435 3927
rect 66177 3893 66211 3927
rect 68201 3893 68235 3927
rect 69857 3893 69891 3927
rect 72065 3893 72099 3927
rect 5825 3689 5859 3723
rect 13737 3689 13771 3723
rect 14841 3689 14875 3723
rect 19993 3689 20027 3723
rect 22017 3689 22051 3723
rect 25605 3689 25639 3723
rect 34069 3689 34103 3723
rect 34713 3689 34747 3723
rect 41245 3689 41279 3723
rect 41981 3689 42015 3723
rect 43563 3689 43597 3723
rect 45569 3689 45603 3723
rect 47409 3689 47443 3723
rect 49617 3689 49651 3723
rect 53205 3689 53239 3723
rect 68661 3689 68695 3723
rect 71697 3689 71731 3723
rect 77585 3689 77619 3723
rect 7297 3621 7331 3655
rect 16129 3621 16163 3655
rect 26525 3621 26559 3655
rect 28457 3621 28491 3655
rect 32045 3621 32079 3655
rect 34621 3621 34655 3655
rect 42073 3621 42107 3655
rect 46673 3621 46707 3655
rect 6561 3553 6595 3587
rect 8217 3553 8251 3587
rect 9689 3553 9723 3587
rect 10241 3553 10275 3587
rect 10885 3553 10919 3587
rect 12265 3553 12299 3587
rect 14381 3553 14415 3587
rect 15301 3553 15335 3587
rect 16681 3553 16715 3587
rect 18153 3553 18187 3587
rect 18705 3553 18739 3587
rect 20821 3553 20855 3587
rect 23949 3553 23983 3587
rect 26341 3553 26375 3587
rect 29377 3553 29411 3587
rect 32321 3553 32355 3587
rect 35265 3553 35299 3587
rect 38577 3553 38611 3587
rect 45937 3553 45971 3587
rect 47225 3553 47259 3587
rect 48697 3553 48731 3587
rect 48881 3553 48915 3587
rect 52377 3553 52411 3587
rect 53849 3553 53883 3587
rect 54033 3553 54067 3587
rect 67833 3553 67867 3587
rect 69213 3553 69247 3587
rect 69489 3553 69523 3587
rect 73721 3553 73755 3587
rect 77033 3553 77067 3587
rect 5273 3485 5307 3519
rect 6745 3485 6779 3519
rect 7389 3485 7423 3519
rect 8033 3485 8067 3519
rect 9045 3485 9079 3519
rect 11989 3485 12023 3519
rect 14197 3485 14231 3519
rect 14289 3485 14323 3519
rect 14657 3485 14691 3519
rect 15577 3485 15611 3519
rect 16313 3485 16347 3519
rect 16405 3485 16439 3519
rect 18245 3485 18279 3519
rect 19809 3485 19843 3519
rect 20361 3485 20395 3519
rect 22293 3485 22327 3519
rect 25145 3485 25179 3519
rect 25329 3485 25363 3519
rect 26709 3485 26743 3519
rect 28733 3485 28767 3519
rect 29101 3485 29135 3519
rect 31677 3485 31711 3519
rect 32229 3485 32263 3519
rect 34161 3485 34195 3519
rect 34437 3485 34471 3519
rect 35633 3485 35667 3519
rect 35725 3485 35759 3519
rect 35909 3485 35943 3519
rect 36093 3485 36127 3519
rect 36369 3485 36403 3519
rect 37289 3485 37323 3519
rect 39129 3485 39163 3519
rect 40601 3485 40635 3519
rect 40969 3485 41003 3519
rect 41061 3485 41095 3519
rect 41245 3485 41279 3519
rect 41337 3485 41371 3519
rect 43821 3485 43855 3519
rect 43913 3485 43947 3519
rect 45385 3485 45419 3519
rect 46581 3485 46615 3519
rect 47961 3485 47995 3519
rect 50261 3485 50295 3519
rect 51825 3485 51859 3519
rect 52469 3485 52503 3519
rect 53021 3485 53055 3519
rect 54585 3485 54619 3519
rect 54677 3485 54711 3519
rect 58081 3485 58115 3519
rect 58173 3485 58207 3519
rect 58725 3485 58759 3519
rect 59461 3485 59495 3519
rect 62037 3485 62071 3519
rect 62129 3485 62163 3519
rect 62681 3485 62715 3519
rect 63417 3485 63451 3519
rect 64521 3485 64555 3519
rect 65073 3485 65107 3519
rect 65717 3485 65751 3519
rect 67281 3485 67315 3519
rect 67925 3485 67959 3519
rect 68477 3485 68511 3519
rect 70041 3485 70075 3519
rect 70133 3485 70167 3519
rect 72341 3485 72375 3519
rect 72433 3485 72467 3519
rect 72985 3485 73019 3519
rect 75101 3485 75135 3519
rect 76665 3485 76699 3519
rect 5917 3417 5951 3451
rect 20269 3417 20303 3451
rect 21985 3417 22019 3451
rect 22201 3417 22235 3451
rect 23213 3417 23247 3451
rect 25605 3417 25639 3451
rect 26065 3417 26099 3451
rect 26157 3417 26191 3451
rect 26985 3417 27019 3451
rect 30665 3417 30699 3451
rect 32597 3417 32631 3451
rect 34253 3417 34287 3451
rect 39405 3417 39439 3451
rect 45109 3417 45143 3451
rect 49525 3417 49559 3451
rect 75469 3417 75503 3451
rect 8769 3349 8803 3383
rect 8953 3349 8987 3383
rect 10793 3349 10827 3383
rect 11529 3349 11563 3383
rect 13829 3349 13863 3383
rect 15485 3349 15519 3383
rect 15945 3349 15979 3383
rect 21833 3349 21867 3383
rect 25421 3349 25455 3383
rect 25697 3349 25731 3383
rect 28641 3349 28675 3383
rect 35081 3349 35115 3383
rect 35173 3349 35207 3383
rect 40785 3349 40819 3383
rect 48145 3349 48179 3383
rect 55321 3349 55355 3383
rect 57437 3349 57471 3383
rect 58909 3349 58943 3383
rect 61393 3349 61427 3383
rect 62865 3349 62899 3383
rect 65165 3349 65199 3383
rect 70777 3349 70811 3383
rect 73169 3349 73203 3383
rect 74549 3349 74583 3383
rect 3801 3145 3835 3179
rect 7297 3145 7331 3179
rect 8217 3145 8251 3179
rect 8953 3145 8987 3179
rect 9689 3145 9723 3179
rect 12265 3145 12299 3179
rect 12909 3145 12943 3179
rect 17417 3145 17451 3179
rect 17601 3145 17635 3179
rect 21649 3145 21683 3179
rect 22569 3145 22603 3179
rect 23029 3145 23063 3179
rect 25053 3145 25087 3179
rect 26985 3145 27019 3179
rect 27445 3145 27479 3179
rect 27537 3145 27571 3179
rect 28549 3145 28583 3179
rect 33517 3145 33551 3179
rect 34069 3145 34103 3179
rect 42073 3145 42107 3179
rect 42717 3145 42751 3179
rect 43177 3145 43211 3179
rect 45109 3145 45143 3179
rect 48145 3145 48179 3179
rect 50813 3145 50847 3179
rect 51733 3145 51767 3179
rect 53849 3145 53883 3179
rect 57345 3145 57379 3179
rect 58081 3145 58115 3179
rect 60933 3145 60967 3179
rect 61669 3145 61703 3179
rect 64521 3145 64555 3179
rect 65441 3145 65475 3179
rect 67189 3145 67223 3179
rect 69305 3145 69339 3179
rect 74457 3145 74491 3179
rect 10793 3077 10827 3111
rect 12633 3077 12667 3111
rect 18337 3077 18371 3111
rect 24501 3077 24535 3111
rect 25421 3077 25455 3111
rect 30021 3077 30055 3111
rect 30481 3077 30515 3111
rect 32413 3077 32447 3111
rect 33425 3077 33459 3111
rect 35633 3077 35667 3111
rect 38669 3077 38703 3111
rect 43637 3077 43671 3111
rect 50077 3077 50111 3111
rect 3249 3009 3283 3043
rect 4905 3009 4939 3043
rect 7481 3009 7515 3043
rect 7573 3009 7607 3043
rect 9781 3009 9815 3043
rect 10425 3009 10459 3043
rect 10517 3009 10551 3043
rect 13093 3009 13127 3043
rect 14933 3009 14967 3043
rect 16865 3009 16899 3043
rect 18061 3009 18095 3043
rect 19901 3009 19935 3043
rect 21925 3009 21959 3043
rect 22753 3009 22787 3043
rect 24777 3009 24811 3043
rect 24869 3009 24903 3043
rect 25145 3009 25179 3043
rect 25237 3009 25271 3043
rect 26893 3009 26927 3043
rect 27353 3009 27387 3043
rect 27997 3009 28031 3043
rect 28181 3009 28215 3043
rect 30389 3009 30423 3043
rect 30665 3009 30699 3043
rect 30849 3009 30883 3043
rect 32689 3009 32723 3043
rect 33885 3009 33919 3043
rect 34069 3009 34103 3043
rect 35909 3009 35943 3043
rect 36185 3009 36219 3043
rect 38393 3009 38427 3043
rect 41981 3009 42015 3043
rect 42257 3009 42291 3043
rect 42809 3009 42843 3043
rect 43361 3009 43395 3043
rect 45201 3009 45235 3043
rect 46765 3009 46799 3043
rect 48329 3009 48363 3043
rect 49801 3009 49835 3043
rect 51365 3009 51399 3043
rect 51549 3009 51583 3043
rect 52101 3009 52135 3043
rect 53665 3009 53699 3043
rect 54033 3009 54067 3043
rect 56057 3009 56091 3043
rect 57161 3009 57195 3043
rect 57437 3009 57471 3043
rect 60749 3009 60783 3043
rect 61117 3009 61151 3043
rect 61761 3009 61795 3043
rect 64705 3009 64739 3043
rect 64889 3009 64923 3043
rect 65533 3009 65567 3043
rect 67005 3009 67039 3043
rect 67649 3009 67683 3043
rect 69121 3009 69155 3043
rect 69489 3009 69523 3043
rect 71513 3009 71547 3043
rect 72985 3009 73019 3043
rect 74273 3009 74307 3043
rect 74549 3009 74583 3043
rect 76665 3009 76699 3043
rect 4353 2941 4387 2975
rect 5089 2941 5123 2975
rect 5641 2941 5675 2975
rect 5733 2941 5767 2975
rect 7113 2941 7147 2975
rect 8309 2941 8343 2975
rect 9137 2941 9171 2975
rect 13369 2941 13403 2975
rect 15209 2941 15243 2975
rect 16681 2941 16715 2975
rect 20177 2941 20211 2975
rect 26433 2941 26467 2975
rect 28089 2941 28123 2975
rect 28273 2941 28307 2975
rect 30308 2941 30342 2975
rect 33609 2941 33643 2975
rect 36461 2941 36495 2975
rect 40233 2941 40267 2975
rect 41705 2941 41739 2975
rect 42533 2941 42567 2975
rect 45661 2941 45695 2975
rect 47133 2941 47167 2975
rect 48789 2941 48823 2975
rect 50629 2941 50663 2975
rect 52561 2941 52595 2975
rect 54493 2941 54527 2975
rect 62221 2941 62255 2975
rect 65993 2941 66027 2975
rect 68017 2941 68051 2975
rect 69949 2941 69983 2975
rect 71973 2941 72007 2975
rect 75469 2941 75503 2975
rect 77309 2941 77343 2975
rect 6377 2873 6411 2907
rect 27169 2873 27203 2907
rect 28457 2873 28491 2907
rect 34161 2873 34195 2907
rect 37933 2873 37967 2907
rect 40141 2873 40175 2907
rect 75193 2873 75227 2907
rect 6469 2805 6503 2839
rect 14841 2805 14875 2839
rect 19809 2805 19843 2839
rect 21833 2805 21867 2839
rect 22937 2805 22971 2839
rect 25421 2805 25455 2839
rect 27721 2805 27755 2839
rect 30941 2805 30975 2839
rect 33057 2805 33091 2839
rect 55505 2805 55539 2839
rect 59369 2805 59403 2839
rect 70961 2805 70995 2839
rect 76757 2805 76791 2839
rect 3801 2601 3835 2635
rect 6377 2601 6411 2635
rect 8585 2601 8619 2635
rect 11161 2601 11195 2635
rect 12449 2601 12483 2635
rect 16865 2601 16899 2635
rect 20821 2601 20855 2635
rect 23305 2601 23339 2635
rect 27077 2601 27111 2635
rect 27353 2601 27387 2635
rect 30481 2601 30515 2635
rect 31401 2601 31435 2635
rect 35725 2601 35759 2635
rect 41613 2601 41647 2635
rect 47409 2601 47443 2635
rect 49985 2601 50019 2635
rect 70869 2601 70903 2635
rect 74089 2601 74123 2635
rect 76849 2601 76883 2635
rect 3065 2533 3099 2567
rect 8217 2533 8251 2567
rect 22753 2533 22787 2567
rect 38209 2533 38243 2567
rect 39129 2533 39163 2567
rect 50721 2533 50755 2567
rect 3249 2465 3283 2499
rect 3985 2465 4019 2499
rect 4537 2465 4571 2499
rect 4997 2465 5031 2499
rect 6561 2465 6595 2499
rect 7113 2465 7147 2499
rect 7665 2465 7699 2499
rect 10057 2465 10091 2499
rect 11805 2465 11839 2499
rect 13093 2465 13127 2499
rect 16497 2465 16531 2499
rect 18245 2465 18279 2499
rect 19533 2465 19567 2499
rect 20177 2465 20211 2499
rect 22109 2465 22143 2499
rect 25329 2465 25363 2499
rect 29837 2465 29871 2499
rect 30849 2465 30883 2499
rect 32229 2465 32263 2499
rect 37105 2465 37139 2499
rect 38577 2465 38611 2499
rect 39957 2465 39991 2499
rect 40969 2465 41003 2499
rect 44833 2465 44867 2499
rect 45385 2465 45419 2499
rect 46765 2465 46799 2499
rect 49433 2465 49467 2499
rect 50537 2465 50571 2499
rect 52101 2465 52135 2499
rect 54033 2465 54067 2499
rect 58173 2465 58207 2499
rect 59277 2465 59311 2499
rect 61761 2465 61795 2499
rect 65533 2465 65567 2499
rect 67649 2465 67683 2499
rect 69489 2465 69523 2499
rect 72617 2465 72651 2499
rect 73169 2465 73203 2499
rect 73537 2465 73571 2499
rect 75745 2465 75779 2499
rect 77401 2465 77435 2499
rect 2513 2397 2547 2431
rect 4721 2397 4755 2431
rect 5641 2397 5675 2431
rect 5733 2397 5767 2431
rect 7481 2397 7515 2431
rect 9137 2397 9171 2431
rect 10609 2397 10643 2431
rect 11713 2397 11747 2431
rect 12081 2397 12115 2431
rect 12817 2397 12851 2431
rect 14657 2397 14691 2431
rect 15301 2397 15335 2431
rect 18061 2397 18095 2431
rect 19809 2397 19843 2431
rect 20913 2397 20947 2431
rect 22477 2397 22511 2431
rect 22937 2397 22971 2431
rect 23397 2397 23431 2431
rect 27537 2397 27571 2431
rect 28089 2397 28123 2431
rect 28273 2397 28307 2431
rect 30297 2397 30331 2431
rect 30665 2397 30699 2431
rect 31493 2397 31527 2431
rect 33057 2397 33091 2431
rect 33425 2397 33459 2431
rect 35265 2397 35299 2431
rect 35633 2397 35667 2431
rect 35817 2397 35851 2431
rect 36001 2397 36035 2431
rect 36829 2397 36863 2431
rect 38393 2397 38427 2431
rect 39405 2397 39439 2431
rect 41245 2397 41279 2431
rect 41981 2397 42015 2431
rect 42993 2397 43027 2431
rect 43361 2397 43395 2431
rect 45753 2397 45787 2431
rect 45937 2397 45971 2431
rect 47961 2397 47995 2431
rect 48329 2397 48363 2431
rect 49709 2397 49743 2431
rect 52837 2397 52871 2431
rect 55045 2397 55079 2431
rect 55505 2397 55539 2431
rect 58633 2397 58667 2431
rect 58817 2397 58851 2431
rect 62773 2397 62807 2431
rect 63233 2397 63267 2431
rect 66269 2397 66303 2431
rect 68293 2397 68327 2431
rect 70501 2397 70535 2431
rect 70685 2397 70719 2431
rect 73077 2397 73111 2431
rect 76205 2397 76239 2431
rect 10333 2329 10367 2363
rect 12909 2329 12943 2363
rect 13645 2329 13679 2363
rect 16957 2329 16991 2363
rect 17325 2329 17359 2363
rect 17969 2329 18003 2363
rect 23121 2329 23155 2363
rect 25605 2329 25639 2363
rect 27721 2329 27755 2363
rect 28825 2329 28859 2363
rect 34253 2329 34287 2363
rect 44281 2329 44315 2363
rect 4905 2261 4939 2295
rect 7297 2261 7331 2295
rect 11253 2261 11287 2295
rect 11621 2261 11655 2295
rect 12265 2261 12299 2295
rect 17601 2261 17635 2295
rect 21097 2261 21131 2295
rect 23029 2261 23063 2295
rect 24685 2261 24719 2295
rect 33241 2261 33275 2295
rect 33977 2261 34011 2295
rect 36553 2261 36587 2295
rect 41153 2261 41187 2295
rect 45569 2261 45603 2295
rect 48145 2261 48179 2295
<< metal1 >>
rect 2024 37562 77924 37584
rect 2024 37510 5134 37562
rect 5186 37510 5198 37562
rect 5250 37510 5262 37562
rect 5314 37510 5326 37562
rect 5378 37510 5390 37562
rect 5442 37510 35854 37562
rect 35906 37510 35918 37562
rect 35970 37510 35982 37562
rect 36034 37510 36046 37562
rect 36098 37510 36110 37562
rect 36162 37510 66574 37562
rect 66626 37510 66638 37562
rect 66690 37510 66702 37562
rect 66754 37510 66766 37562
rect 66818 37510 66830 37562
rect 66882 37510 77924 37562
rect 2024 37488 77924 37510
rect 2222 37272 2228 37324
rect 2280 37312 2286 37324
rect 2501 37315 2559 37321
rect 2501 37312 2513 37315
rect 2280 37284 2513 37312
rect 2280 37272 2286 37284
rect 2501 37281 2513 37284
rect 2547 37281 2559 37315
rect 2501 37275 2559 37281
rect 13262 37272 13268 37324
rect 13320 37312 13326 37324
rect 13541 37315 13599 37321
rect 13541 37312 13553 37315
rect 13320 37284 13553 37312
rect 13320 37272 13326 37284
rect 13541 37281 13553 37284
rect 13587 37281 13599 37315
rect 13541 37275 13599 37281
rect 33502 37272 33508 37324
rect 33560 37312 33566 37324
rect 34057 37315 34115 37321
rect 34057 37312 34069 37315
rect 33560 37284 34069 37312
rect 33560 37272 33566 37284
rect 34057 37281 34069 37284
rect 34103 37281 34115 37315
rect 34057 37275 34115 37281
rect 39022 37272 39028 37324
rect 39080 37312 39086 37324
rect 39577 37315 39635 37321
rect 39577 37312 39589 37315
rect 39080 37284 39589 37312
rect 39080 37272 39086 37284
rect 39577 37281 39589 37284
rect 39623 37281 39635 37315
rect 39577 37275 39635 37281
rect 3510 37204 3516 37256
rect 3568 37204 3574 37256
rect 5902 37204 5908 37256
rect 5960 37204 5966 37256
rect 7098 37204 7104 37256
rect 7156 37204 7162 37256
rect 7742 37204 7748 37256
rect 7800 37244 7806 37256
rect 7837 37247 7895 37253
rect 7837 37244 7849 37247
rect 7800 37216 7849 37244
rect 7800 37204 7806 37216
rect 7837 37213 7849 37216
rect 7883 37213 7895 37247
rect 7837 37207 7895 37213
rect 7926 37204 7932 37256
rect 7984 37244 7990 37256
rect 8757 37247 8815 37253
rect 8757 37244 8769 37247
rect 7984 37216 8769 37244
rect 7984 37204 7990 37216
rect 8757 37213 8769 37216
rect 8803 37213 8815 37247
rect 8757 37207 8815 37213
rect 11333 37247 11391 37253
rect 11333 37213 11345 37247
rect 11379 37244 11391 37247
rect 11422 37244 11428 37256
rect 11379 37216 11428 37244
rect 11379 37213 11391 37216
rect 11333 37207 11391 37213
rect 11422 37204 11428 37216
rect 11480 37204 11486 37256
rect 11882 37204 11888 37256
rect 11940 37244 11946 37256
rect 12069 37247 12127 37253
rect 12069 37244 12081 37247
rect 11940 37216 12081 37244
rect 11940 37204 11946 37216
rect 12069 37213 12081 37216
rect 12115 37213 12127 37247
rect 12069 37207 12127 37213
rect 14550 37204 14556 37256
rect 14608 37204 14614 37256
rect 15102 37204 15108 37256
rect 15160 37244 15166 37256
rect 15197 37247 15255 37253
rect 15197 37244 15209 37247
rect 15160 37216 15209 37244
rect 15160 37204 15166 37216
rect 15197 37213 15209 37216
rect 15243 37213 15255 37247
rect 15197 37207 15255 37213
rect 18690 37204 18696 37256
rect 18748 37204 18754 37256
rect 18782 37204 18788 37256
rect 18840 37244 18846 37256
rect 19521 37247 19579 37253
rect 19521 37244 19533 37247
rect 18840 37216 19533 37244
rect 18840 37204 18846 37216
rect 19521 37213 19533 37216
rect 19567 37213 19579 37247
rect 19521 37207 19579 37213
rect 20622 37204 20628 37256
rect 20680 37244 20686 37256
rect 20901 37247 20959 37253
rect 20901 37244 20913 37247
rect 20680 37216 20913 37244
rect 20680 37204 20686 37216
rect 20901 37213 20913 37216
rect 20947 37213 20959 37247
rect 20901 37207 20959 37213
rect 21910 37204 21916 37256
rect 21968 37204 21974 37256
rect 22462 37204 22468 37256
rect 22520 37244 22526 37256
rect 22741 37247 22799 37253
rect 22741 37244 22753 37247
rect 22520 37216 22753 37244
rect 22520 37204 22526 37216
rect 22741 37213 22753 37216
rect 22787 37213 22799 37247
rect 22741 37207 22799 37213
rect 26050 37204 26056 37256
rect 26108 37244 26114 37256
rect 26237 37247 26295 37253
rect 26237 37244 26249 37247
rect 26108 37216 26249 37244
rect 26108 37204 26114 37216
rect 26237 37213 26249 37216
rect 26283 37213 26295 37247
rect 26237 37207 26295 37213
rect 27982 37204 27988 37256
rect 28040 37244 28046 37256
rect 28261 37247 28319 37253
rect 28261 37244 28273 37247
rect 28040 37216 28273 37244
rect 28040 37204 28046 37216
rect 28261 37213 28273 37216
rect 28307 37213 28319 37247
rect 28261 37207 28319 37213
rect 29457 37247 29515 37253
rect 29457 37213 29469 37247
rect 29503 37213 29515 37247
rect 29457 37207 29515 37213
rect 15010 37136 15016 37188
rect 15068 37176 15074 37188
rect 16117 37179 16175 37185
rect 16117 37176 16129 37179
rect 15068 37148 16129 37176
rect 15068 37136 15074 37148
rect 16117 37145 16129 37148
rect 16163 37145 16175 37179
rect 16117 37139 16175 37145
rect 22554 37136 22560 37188
rect 22612 37176 22618 37188
rect 23661 37179 23719 37185
rect 23661 37176 23673 37179
rect 22612 37148 23673 37176
rect 22612 37136 22618 37148
rect 23661 37145 23673 37148
rect 23707 37145 23719 37179
rect 23661 37139 23719 37145
rect 26142 37136 26148 37188
rect 26200 37176 26206 37188
rect 27157 37179 27215 37185
rect 27157 37176 27169 37179
rect 26200 37148 27169 37176
rect 26200 37136 26206 37148
rect 27157 37145 27169 37148
rect 27203 37145 27215 37179
rect 29472 37176 29500 37207
rect 31662 37204 31668 37256
rect 31720 37244 31726 37256
rect 31757 37247 31815 37253
rect 31757 37244 31769 37247
rect 31720 37216 31769 37244
rect 31720 37204 31726 37216
rect 31757 37213 31769 37216
rect 31803 37213 31815 37247
rect 31757 37207 31815 37213
rect 32674 37204 32680 37256
rect 32732 37204 32738 37256
rect 33778 37204 33784 37256
rect 33836 37204 33842 37256
rect 36817 37247 36875 37253
rect 36817 37213 36829 37247
rect 36863 37244 36875 37247
rect 36998 37244 37004 37256
rect 36863 37216 37004 37244
rect 36863 37213 36875 37216
rect 36817 37207 36875 37213
rect 36998 37204 37004 37216
rect 37056 37204 37062 37256
rect 37182 37204 37188 37256
rect 37240 37244 37246 37256
rect 37553 37247 37611 37253
rect 37553 37244 37565 37247
rect 37240 37216 37565 37244
rect 37240 37204 37246 37216
rect 37553 37213 37565 37216
rect 37599 37213 37611 37247
rect 37553 37207 37611 37213
rect 39114 37204 39120 37256
rect 39172 37204 39178 37256
rect 40862 37204 40868 37256
rect 40920 37244 40926 37256
rect 40957 37247 41015 37253
rect 40957 37244 40969 37247
rect 40920 37216 40969 37244
rect 40920 37204 40926 37216
rect 40957 37213 40969 37216
rect 41003 37213 41015 37247
rect 40957 37207 41015 37213
rect 41046 37204 41052 37256
rect 41104 37244 41110 37256
rect 41877 37247 41935 37253
rect 41877 37244 41889 37247
rect 41104 37216 41889 37244
rect 41104 37204 41110 37216
rect 41877 37213 41889 37216
rect 41923 37213 41935 37247
rect 41877 37207 41935 37213
rect 43346 37204 43352 37256
rect 43404 37204 43410 37256
rect 46474 37204 46480 37256
rect 46532 37204 46538 37256
rect 48222 37204 48228 37256
rect 48280 37244 48286 37256
rect 48501 37247 48559 37253
rect 48501 37244 48513 37247
rect 48280 37216 48513 37244
rect 48280 37204 48286 37216
rect 48501 37213 48513 37216
rect 48547 37213 48559 37247
rect 48501 37207 48559 37213
rect 51902 37204 51908 37256
rect 51960 37244 51966 37256
rect 51997 37247 52055 37253
rect 51997 37244 52009 37247
rect 51960 37216 52009 37244
rect 51960 37204 51966 37216
rect 51997 37213 52009 37216
rect 52043 37213 52055 37247
rect 51997 37207 52055 37213
rect 52086 37204 52092 37256
rect 52144 37244 52150 37256
rect 52917 37247 52975 37253
rect 52917 37244 52929 37247
rect 52144 37216 52929 37244
rect 52144 37204 52150 37216
rect 52917 37213 52929 37216
rect 52963 37213 52975 37247
rect 52917 37207 52975 37213
rect 53834 37204 53840 37256
rect 53892 37204 53898 37256
rect 55582 37204 55588 37256
rect 55640 37244 55646 37256
rect 56229 37247 56287 37253
rect 56229 37244 56241 37247
rect 55640 37216 56241 37244
rect 55640 37204 55646 37216
rect 56229 37213 56241 37216
rect 56275 37213 56287 37247
rect 56229 37207 56287 37213
rect 58802 37204 58808 37256
rect 58860 37204 58866 37256
rect 33042 37176 33048 37188
rect 29472 37148 33048 37176
rect 27157 37139 27215 37145
rect 33042 37136 33048 37148
rect 33100 37136 33106 37188
rect 42702 37136 42708 37188
rect 42760 37176 42766 37188
rect 44269 37179 44327 37185
rect 44269 37176 44281 37179
rect 42760 37148 44281 37176
rect 42760 37136 42766 37148
rect 44269 37145 44281 37148
rect 44315 37145 44327 37179
rect 44269 37139 44327 37145
rect 46382 37136 46388 37188
rect 46440 37176 46446 37188
rect 47397 37179 47455 37185
rect 47397 37176 47409 37179
rect 46440 37148 47409 37176
rect 46440 37136 46446 37148
rect 47397 37145 47409 37148
rect 47443 37145 47455 37179
rect 47397 37139 47455 37145
rect 48130 37136 48136 37188
rect 48188 37176 48194 37188
rect 49421 37179 49479 37185
rect 49421 37176 49433 37179
rect 48188 37148 49433 37176
rect 48188 37136 48194 37148
rect 49421 37145 49433 37148
rect 49467 37145 49479 37179
rect 49421 37139 49479 37145
rect 53742 37136 53748 37188
rect 53800 37176 53806 37188
rect 54757 37179 54815 37185
rect 54757 37176 54769 37179
rect 53800 37148 54769 37176
rect 53800 37136 53806 37148
rect 54757 37145 54769 37148
rect 54803 37145 54815 37179
rect 54757 37139 54815 37145
rect 55674 37136 55680 37188
rect 55732 37176 55738 37188
rect 57149 37179 57207 37185
rect 57149 37176 57161 37179
rect 55732 37148 57161 37176
rect 55732 37136 55738 37148
rect 57149 37145 57161 37148
rect 57195 37145 57207 37179
rect 57149 37139 57207 37145
rect 57422 37136 57428 37188
rect 57480 37176 57486 37188
rect 59725 37179 59783 37185
rect 59725 37176 59737 37179
rect 57480 37148 59737 37176
rect 57480 37136 57486 37148
rect 59725 37145 59737 37148
rect 59771 37145 59783 37179
rect 59725 37139 59783 37145
rect 2024 37018 77924 37040
rect 2024 36966 5794 37018
rect 5846 36966 5858 37018
rect 5910 36966 5922 37018
rect 5974 36966 5986 37018
rect 6038 36966 6050 37018
rect 6102 36966 36514 37018
rect 36566 36966 36578 37018
rect 36630 36966 36642 37018
rect 36694 36966 36706 37018
rect 36758 36966 36770 37018
rect 36822 36966 67234 37018
rect 67286 36966 67298 37018
rect 67350 36966 67362 37018
rect 67414 36966 67426 37018
rect 67478 36966 67490 37018
rect 67542 36966 77924 37018
rect 2024 36944 77924 36966
rect 7742 36864 7748 36916
rect 7800 36864 7806 36916
rect 11882 36864 11888 36916
rect 11940 36864 11946 36916
rect 15102 36864 15108 36916
rect 15160 36864 15166 36916
rect 18690 36864 18696 36916
rect 18748 36904 18754 36916
rect 19061 36907 19119 36913
rect 19061 36904 19073 36907
rect 18748 36876 19073 36904
rect 18748 36864 18754 36876
rect 19061 36873 19073 36876
rect 19107 36873 19119 36907
rect 19061 36867 19119 36873
rect 22462 36864 22468 36916
rect 22520 36864 22526 36916
rect 26050 36864 26056 36916
rect 26108 36904 26114 36916
rect 26145 36907 26203 36913
rect 26145 36904 26157 36907
rect 26108 36876 26157 36904
rect 26108 36864 26114 36876
rect 26145 36873 26157 36876
rect 26191 36873 26203 36907
rect 26145 36867 26203 36873
rect 29656 36876 30604 36904
rect 4062 36796 4068 36848
rect 4120 36836 4126 36848
rect 4341 36839 4399 36845
rect 4341 36836 4353 36839
rect 4120 36808 4353 36836
rect 4120 36796 4126 36808
rect 4341 36805 4353 36808
rect 4387 36805 4399 36839
rect 4341 36799 4399 36805
rect 9582 36796 9588 36848
rect 9640 36836 9646 36848
rect 9861 36839 9919 36845
rect 9861 36836 9873 36839
rect 9640 36808 9873 36836
rect 9640 36796 9646 36808
rect 9861 36805 9873 36808
rect 9907 36805 9919 36839
rect 9861 36799 9919 36805
rect 16942 36796 16948 36848
rect 17000 36836 17006 36848
rect 17957 36839 18015 36845
rect 17957 36836 17969 36839
rect 17000 36808 17969 36836
rect 17000 36796 17006 36808
rect 17957 36805 17969 36808
rect 18003 36805 18015 36839
rect 17957 36799 18015 36805
rect 24302 36796 24308 36848
rect 24360 36836 24366 36848
rect 24581 36839 24639 36845
rect 24581 36836 24593 36839
rect 24360 36808 24593 36836
rect 24360 36796 24366 36808
rect 24581 36805 24593 36808
rect 24627 36805 24639 36839
rect 24581 36799 24639 36805
rect 5445 36771 5503 36777
rect 5445 36737 5457 36771
rect 5491 36768 5503 36771
rect 7561 36771 7619 36777
rect 7561 36768 7573 36771
rect 5491 36740 7573 36768
rect 5491 36737 5503 36740
rect 5445 36731 5503 36737
rect 7561 36737 7573 36740
rect 7607 36737 7619 36771
rect 7561 36731 7619 36737
rect 7576 36700 7604 36731
rect 10962 36728 10968 36780
rect 11020 36728 11026 36780
rect 11790 36728 11796 36780
rect 11848 36728 11854 36780
rect 12069 36771 12127 36777
rect 12069 36737 12081 36771
rect 12115 36768 12127 36771
rect 14921 36771 14979 36777
rect 14921 36768 14933 36771
rect 12115 36740 14933 36768
rect 12115 36737 12127 36740
rect 12069 36731 12127 36737
rect 14921 36737 14933 36740
rect 14967 36737 14979 36771
rect 14921 36731 14979 36737
rect 11609 36703 11667 36709
rect 11609 36700 11621 36703
rect 7576 36672 11621 36700
rect 11609 36669 11621 36672
rect 11655 36700 11667 36703
rect 12084 36700 12112 36731
rect 11655 36672 12112 36700
rect 14936 36700 14964 36731
rect 18782 36728 18788 36780
rect 18840 36728 18846 36780
rect 19245 36771 19303 36777
rect 19245 36737 19257 36771
rect 19291 36768 19303 36771
rect 22281 36771 22339 36777
rect 22281 36768 22293 36771
rect 19291 36740 22293 36768
rect 19291 36737 19303 36740
rect 19245 36731 19303 36737
rect 22281 36737 22293 36740
rect 22327 36737 22339 36771
rect 22281 36731 22339 36737
rect 19260 36700 19288 36731
rect 14936 36672 19288 36700
rect 22296 36700 22324 36731
rect 25774 36728 25780 36780
rect 25832 36728 25838 36780
rect 29656 36777 29684 36876
rect 29822 36796 29828 36848
rect 29880 36836 29886 36848
rect 30576 36836 30604 36876
rect 33778 36864 33784 36916
rect 33836 36864 33842 36916
rect 33888 36876 36952 36904
rect 33888 36836 33916 36876
rect 36924 36836 36952 36876
rect 36998 36864 37004 36916
rect 37056 36864 37062 36916
rect 40862 36864 40868 36916
rect 40920 36864 40926 36916
rect 48222 36864 48228 36916
rect 48280 36864 48286 36916
rect 51902 36864 51908 36916
rect 51960 36864 51966 36916
rect 55582 36864 55588 36916
rect 55640 36864 55646 36916
rect 29880 36808 30420 36836
rect 30576 36808 33916 36836
rect 33980 36808 35894 36836
rect 36924 36808 55214 36836
rect 29880 36796 29886 36808
rect 25961 36771 26019 36777
rect 25961 36737 25973 36771
rect 26007 36768 26019 36771
rect 29641 36771 29699 36777
rect 29641 36768 29653 36771
rect 26007 36740 29653 36768
rect 26007 36737 26019 36740
rect 25961 36731 26019 36737
rect 29641 36737 29653 36740
rect 29687 36737 29699 36771
rect 29917 36771 29975 36777
rect 29917 36768 29929 36771
rect 29641 36731 29699 36737
rect 29840 36740 29929 36768
rect 25976 36700 26004 36731
rect 22296 36672 26004 36700
rect 11655 36669 11667 36672
rect 11609 36663 11667 36669
rect 11790 36592 11796 36644
rect 11848 36632 11854 36644
rect 29840 36641 29868 36740
rect 29917 36737 29929 36740
rect 29963 36737 29975 36771
rect 29917 36731 29975 36737
rect 30392 36709 30420 36808
rect 33980 36777 34008 36808
rect 33505 36771 33563 36777
rect 33505 36737 33517 36771
rect 33551 36737 33563 36771
rect 33505 36731 33563 36737
rect 33689 36771 33747 36777
rect 33689 36737 33701 36771
rect 33735 36768 33747 36771
rect 33965 36771 34023 36777
rect 33965 36768 33977 36771
rect 33735 36740 33977 36768
rect 33735 36737 33747 36740
rect 33689 36731 33747 36737
rect 33965 36737 33977 36740
rect 34011 36737 34023 36771
rect 33965 36731 34023 36737
rect 30377 36703 30435 36709
rect 30377 36669 30389 36703
rect 30423 36669 30435 36703
rect 30377 36663 30435 36669
rect 29825 36635 29883 36641
rect 11848 36604 26234 36632
rect 11848 36592 11854 36604
rect 26206 36564 26234 36604
rect 29825 36601 29837 36635
rect 29871 36601 29883 36635
rect 29825 36595 29883 36601
rect 33520 36564 33548 36731
rect 35434 36728 35440 36780
rect 35492 36728 35498 36780
rect 35866 36768 35894 36808
rect 37185 36771 37243 36777
rect 37185 36768 37197 36771
rect 35866 36740 37197 36768
rect 37185 36737 37197 36740
rect 37231 36768 37243 36771
rect 40681 36771 40739 36777
rect 40681 36768 40693 36771
rect 37231 36740 40693 36768
rect 37231 36737 37243 36740
rect 37185 36731 37243 36737
rect 40681 36737 40693 36740
rect 40727 36768 40739 36771
rect 44361 36771 44419 36777
rect 44361 36768 44373 36771
rect 40727 36740 44373 36768
rect 40727 36737 40739 36740
rect 40681 36731 40739 36737
rect 44361 36737 44373 36740
rect 44407 36737 44419 36771
rect 44637 36771 44695 36777
rect 44637 36768 44649 36771
rect 44361 36731 44419 36737
rect 44560 36740 44649 36768
rect 35342 36660 35348 36712
rect 35400 36700 35406 36712
rect 35897 36703 35955 36709
rect 35897 36700 35909 36703
rect 35400 36672 35909 36700
rect 35400 36660 35406 36672
rect 35897 36669 35909 36672
rect 35943 36669 35955 36703
rect 35897 36663 35955 36669
rect 26206 36536 33548 36564
rect 44376 36564 44404 36731
rect 44560 36641 44588 36740
rect 44637 36737 44649 36740
rect 44683 36737 44695 36771
rect 44637 36731 44695 36737
rect 48041 36771 48099 36777
rect 48041 36737 48053 36771
rect 48087 36737 48099 36771
rect 48041 36731 48099 36737
rect 44726 36660 44732 36712
rect 44784 36700 44790 36712
rect 45097 36703 45155 36709
rect 45097 36700 45109 36703
rect 44784 36672 45109 36700
rect 44784 36660 44790 36672
rect 45097 36669 45109 36672
rect 45143 36669 45155 36703
rect 45097 36663 45155 36669
rect 44545 36635 44603 36641
rect 44545 36601 44557 36635
rect 44591 36601 44603 36635
rect 48056 36632 48084 36731
rect 50154 36728 50160 36780
rect 50212 36728 50218 36780
rect 51721 36771 51779 36777
rect 51721 36737 51733 36771
rect 51767 36737 51779 36771
rect 55186 36768 55214 36808
rect 59262 36796 59268 36848
rect 59320 36836 59326 36848
rect 59320 36808 59860 36836
rect 59320 36796 59326 36808
rect 55401 36771 55459 36777
rect 55401 36768 55413 36771
rect 55186 36740 55413 36768
rect 51721 36731 51779 36737
rect 55401 36737 55413 36740
rect 55447 36768 55459 36771
rect 58437 36771 58495 36777
rect 58437 36768 58449 36771
rect 55447 36740 58449 36768
rect 55447 36737 55459 36740
rect 55401 36731 55459 36737
rect 58437 36737 58449 36740
rect 58483 36737 58495 36771
rect 58437 36731 58495 36737
rect 59357 36771 59415 36777
rect 59357 36737 59369 36771
rect 59403 36737 59415 36771
rect 59357 36731 59415 36737
rect 50062 36660 50068 36712
rect 50120 36700 50126 36712
rect 50617 36703 50675 36709
rect 50617 36700 50629 36703
rect 50120 36672 50629 36700
rect 50120 36660 50126 36672
rect 50617 36669 50629 36672
rect 50663 36669 50675 36703
rect 50617 36663 50675 36669
rect 51736 36632 51764 36731
rect 44545 36595 44603 36601
rect 45526 36604 51764 36632
rect 58621 36635 58679 36641
rect 45526 36564 45554 36604
rect 58621 36601 58633 36635
rect 58667 36632 58679 36635
rect 59372 36632 59400 36731
rect 59832 36709 59860 36808
rect 59817 36703 59875 36709
rect 59817 36669 59829 36703
rect 59863 36669 59875 36703
rect 59817 36663 59875 36669
rect 58667 36604 59400 36632
rect 58667 36601 58679 36604
rect 58621 36595 58679 36601
rect 44376 36536 45554 36564
rect 2024 36474 77924 36496
rect 2024 36422 5134 36474
rect 5186 36422 5198 36474
rect 5250 36422 5262 36474
rect 5314 36422 5326 36474
rect 5378 36422 5390 36474
rect 5442 36422 35854 36474
rect 35906 36422 35918 36474
rect 35970 36422 35982 36474
rect 36034 36422 36046 36474
rect 36098 36422 36110 36474
rect 36162 36422 66574 36474
rect 66626 36422 66638 36474
rect 66690 36422 66702 36474
rect 66754 36422 66766 36474
rect 66818 36422 66830 36474
rect 66882 36422 77924 36474
rect 2024 36400 77924 36422
rect 25774 36320 25780 36372
rect 25832 36360 25838 36372
rect 33226 36360 33232 36372
rect 25832 36332 33232 36360
rect 25832 36320 25838 36332
rect 33226 36320 33232 36332
rect 33284 36320 33290 36372
rect 2024 35930 77924 35952
rect 2024 35878 5794 35930
rect 5846 35878 5858 35930
rect 5910 35878 5922 35930
rect 5974 35878 5986 35930
rect 6038 35878 6050 35930
rect 6102 35878 36514 35930
rect 36566 35878 36578 35930
rect 36630 35878 36642 35930
rect 36694 35878 36706 35930
rect 36758 35878 36770 35930
rect 36822 35878 67234 35930
rect 67286 35878 67298 35930
rect 67350 35878 67362 35930
rect 67414 35878 67426 35930
rect 67478 35878 67490 35930
rect 67542 35878 77924 35930
rect 2024 35856 77924 35878
rect 2024 35386 77924 35408
rect 2024 35334 5134 35386
rect 5186 35334 5198 35386
rect 5250 35334 5262 35386
rect 5314 35334 5326 35386
rect 5378 35334 5390 35386
rect 5442 35334 35854 35386
rect 35906 35334 35918 35386
rect 35970 35334 35982 35386
rect 36034 35334 36046 35386
rect 36098 35334 36110 35386
rect 36162 35334 66574 35386
rect 66626 35334 66638 35386
rect 66690 35334 66702 35386
rect 66754 35334 66766 35386
rect 66818 35334 66830 35386
rect 66882 35334 77924 35386
rect 2024 35312 77924 35334
rect 2024 34842 77924 34864
rect 2024 34790 5794 34842
rect 5846 34790 5858 34842
rect 5910 34790 5922 34842
rect 5974 34790 5986 34842
rect 6038 34790 6050 34842
rect 6102 34790 36514 34842
rect 36566 34790 36578 34842
rect 36630 34790 36642 34842
rect 36694 34790 36706 34842
rect 36758 34790 36770 34842
rect 36822 34790 67234 34842
rect 67286 34790 67298 34842
rect 67350 34790 67362 34842
rect 67414 34790 67426 34842
rect 67478 34790 67490 34842
rect 67542 34790 77924 34842
rect 2024 34768 77924 34790
rect 2024 34298 77924 34320
rect 2024 34246 5134 34298
rect 5186 34246 5198 34298
rect 5250 34246 5262 34298
rect 5314 34246 5326 34298
rect 5378 34246 5390 34298
rect 5442 34246 35854 34298
rect 35906 34246 35918 34298
rect 35970 34246 35982 34298
rect 36034 34246 36046 34298
rect 36098 34246 36110 34298
rect 36162 34246 66574 34298
rect 66626 34246 66638 34298
rect 66690 34246 66702 34298
rect 66754 34246 66766 34298
rect 66818 34246 66830 34298
rect 66882 34246 77924 34298
rect 2024 34224 77924 34246
rect 2024 33754 77924 33776
rect 2024 33702 5794 33754
rect 5846 33702 5858 33754
rect 5910 33702 5922 33754
rect 5974 33702 5986 33754
rect 6038 33702 6050 33754
rect 6102 33702 36514 33754
rect 36566 33702 36578 33754
rect 36630 33702 36642 33754
rect 36694 33702 36706 33754
rect 36758 33702 36770 33754
rect 36822 33702 67234 33754
rect 67286 33702 67298 33754
rect 67350 33702 67362 33754
rect 67414 33702 67426 33754
rect 67478 33702 67490 33754
rect 67542 33702 77924 33754
rect 2024 33680 77924 33702
rect 2024 33210 77924 33232
rect 2024 33158 5134 33210
rect 5186 33158 5198 33210
rect 5250 33158 5262 33210
rect 5314 33158 5326 33210
rect 5378 33158 5390 33210
rect 5442 33158 35854 33210
rect 35906 33158 35918 33210
rect 35970 33158 35982 33210
rect 36034 33158 36046 33210
rect 36098 33158 36110 33210
rect 36162 33158 66574 33210
rect 66626 33158 66638 33210
rect 66690 33158 66702 33210
rect 66754 33158 66766 33210
rect 66818 33158 66830 33210
rect 66882 33158 77924 33210
rect 2024 33136 77924 33158
rect 2024 32666 77924 32688
rect 2024 32614 5794 32666
rect 5846 32614 5858 32666
rect 5910 32614 5922 32666
rect 5974 32614 5986 32666
rect 6038 32614 6050 32666
rect 6102 32614 36514 32666
rect 36566 32614 36578 32666
rect 36630 32614 36642 32666
rect 36694 32614 36706 32666
rect 36758 32614 36770 32666
rect 36822 32614 67234 32666
rect 67286 32614 67298 32666
rect 67350 32614 67362 32666
rect 67414 32614 67426 32666
rect 67478 32614 67490 32666
rect 67542 32614 77924 32666
rect 2024 32592 77924 32614
rect 27246 32376 27252 32428
rect 27304 32416 27310 32428
rect 50154 32416 50160 32428
rect 27304 32388 50160 32416
rect 27304 32376 27310 32388
rect 50154 32376 50160 32388
rect 50212 32376 50218 32428
rect 2024 32122 77924 32144
rect 2024 32070 5134 32122
rect 5186 32070 5198 32122
rect 5250 32070 5262 32122
rect 5314 32070 5326 32122
rect 5378 32070 5390 32122
rect 5442 32070 35854 32122
rect 35906 32070 35918 32122
rect 35970 32070 35982 32122
rect 36034 32070 36046 32122
rect 36098 32070 36110 32122
rect 36162 32070 66574 32122
rect 66626 32070 66638 32122
rect 66690 32070 66702 32122
rect 66754 32070 66766 32122
rect 66818 32070 66830 32122
rect 66882 32070 77924 32122
rect 2024 32048 77924 32070
rect 2024 31578 77924 31600
rect 2024 31526 5794 31578
rect 5846 31526 5858 31578
rect 5910 31526 5922 31578
rect 5974 31526 5986 31578
rect 6038 31526 6050 31578
rect 6102 31526 36514 31578
rect 36566 31526 36578 31578
rect 36630 31526 36642 31578
rect 36694 31526 36706 31578
rect 36758 31526 36770 31578
rect 36822 31526 67234 31578
rect 67286 31526 67298 31578
rect 67350 31526 67362 31578
rect 67414 31526 67426 31578
rect 67478 31526 67490 31578
rect 67542 31526 77924 31578
rect 2024 31504 77924 31526
rect 2024 31034 77924 31056
rect 2024 30982 5134 31034
rect 5186 30982 5198 31034
rect 5250 30982 5262 31034
rect 5314 30982 5326 31034
rect 5378 30982 5390 31034
rect 5442 30982 35854 31034
rect 35906 30982 35918 31034
rect 35970 30982 35982 31034
rect 36034 30982 36046 31034
rect 36098 30982 36110 31034
rect 36162 30982 66574 31034
rect 66626 30982 66638 31034
rect 66690 30982 66702 31034
rect 66754 30982 66766 31034
rect 66818 30982 66830 31034
rect 66882 30982 77924 31034
rect 2024 30960 77924 30982
rect 2024 30490 77924 30512
rect 2024 30438 5794 30490
rect 5846 30438 5858 30490
rect 5910 30438 5922 30490
rect 5974 30438 5986 30490
rect 6038 30438 6050 30490
rect 6102 30438 36514 30490
rect 36566 30438 36578 30490
rect 36630 30438 36642 30490
rect 36694 30438 36706 30490
rect 36758 30438 36770 30490
rect 36822 30438 67234 30490
rect 67286 30438 67298 30490
rect 67350 30438 67362 30490
rect 67414 30438 67426 30490
rect 67478 30438 67490 30490
rect 67542 30438 77924 30490
rect 2024 30416 77924 30438
rect 2024 29946 77924 29968
rect 2024 29894 5134 29946
rect 5186 29894 5198 29946
rect 5250 29894 5262 29946
rect 5314 29894 5326 29946
rect 5378 29894 5390 29946
rect 5442 29894 35854 29946
rect 35906 29894 35918 29946
rect 35970 29894 35982 29946
rect 36034 29894 36046 29946
rect 36098 29894 36110 29946
rect 36162 29894 66574 29946
rect 66626 29894 66638 29946
rect 66690 29894 66702 29946
rect 66754 29894 66766 29946
rect 66818 29894 66830 29946
rect 66882 29894 77924 29946
rect 2024 29872 77924 29894
rect 24946 29588 24952 29640
rect 25004 29628 25010 29640
rect 53834 29628 53840 29640
rect 25004 29600 53840 29628
rect 25004 29588 25010 29600
rect 53834 29588 53840 29600
rect 53892 29588 53898 29640
rect 2024 29402 77924 29424
rect 2024 29350 5794 29402
rect 5846 29350 5858 29402
rect 5910 29350 5922 29402
rect 5974 29350 5986 29402
rect 6038 29350 6050 29402
rect 6102 29350 36514 29402
rect 36566 29350 36578 29402
rect 36630 29350 36642 29402
rect 36694 29350 36706 29402
rect 36758 29350 36770 29402
rect 36822 29350 67234 29402
rect 67286 29350 67298 29402
rect 67350 29350 67362 29402
rect 67414 29350 67426 29402
rect 67478 29350 67490 29402
rect 67542 29350 77924 29402
rect 2024 29328 77924 29350
rect 2024 28858 77924 28880
rect 2024 28806 5134 28858
rect 5186 28806 5198 28858
rect 5250 28806 5262 28858
rect 5314 28806 5326 28858
rect 5378 28806 5390 28858
rect 5442 28806 35854 28858
rect 35906 28806 35918 28858
rect 35970 28806 35982 28858
rect 36034 28806 36046 28858
rect 36098 28806 36110 28858
rect 36162 28806 66574 28858
rect 66626 28806 66638 28858
rect 66690 28806 66702 28858
rect 66754 28806 66766 28858
rect 66818 28806 66830 28858
rect 66882 28806 77924 28858
rect 2024 28784 77924 28806
rect 2024 28314 77924 28336
rect 2024 28262 5794 28314
rect 5846 28262 5858 28314
rect 5910 28262 5922 28314
rect 5974 28262 5986 28314
rect 6038 28262 6050 28314
rect 6102 28262 36514 28314
rect 36566 28262 36578 28314
rect 36630 28262 36642 28314
rect 36694 28262 36706 28314
rect 36758 28262 36770 28314
rect 36822 28262 67234 28314
rect 67286 28262 67298 28314
rect 67350 28262 67362 28314
rect 67414 28262 67426 28314
rect 67478 28262 67490 28314
rect 67542 28262 77924 28314
rect 2024 28240 77924 28262
rect 2024 27770 77924 27792
rect 2024 27718 5134 27770
rect 5186 27718 5198 27770
rect 5250 27718 5262 27770
rect 5314 27718 5326 27770
rect 5378 27718 5390 27770
rect 5442 27718 35854 27770
rect 35906 27718 35918 27770
rect 35970 27718 35982 27770
rect 36034 27718 36046 27770
rect 36098 27718 36110 27770
rect 36162 27718 66574 27770
rect 66626 27718 66638 27770
rect 66690 27718 66702 27770
rect 66754 27718 66766 27770
rect 66818 27718 66830 27770
rect 66882 27718 77924 27770
rect 2024 27696 77924 27718
rect 2024 27226 77924 27248
rect 2024 27174 5794 27226
rect 5846 27174 5858 27226
rect 5910 27174 5922 27226
rect 5974 27174 5986 27226
rect 6038 27174 6050 27226
rect 6102 27174 36514 27226
rect 36566 27174 36578 27226
rect 36630 27174 36642 27226
rect 36694 27174 36706 27226
rect 36758 27174 36770 27226
rect 36822 27174 67234 27226
rect 67286 27174 67298 27226
rect 67350 27174 67362 27226
rect 67414 27174 67426 27226
rect 67478 27174 67490 27226
rect 67542 27174 77924 27226
rect 2024 27152 77924 27174
rect 18782 26936 18788 26988
rect 18840 26976 18846 26988
rect 34790 26976 34796 26988
rect 18840 26948 34796 26976
rect 18840 26936 18846 26948
rect 34790 26936 34796 26948
rect 34848 26936 34854 26988
rect 26234 26868 26240 26920
rect 26292 26908 26298 26920
rect 46474 26908 46480 26920
rect 26292 26880 46480 26908
rect 26292 26868 26298 26880
rect 46474 26868 46480 26880
rect 46532 26868 46538 26920
rect 2024 26682 77924 26704
rect 2024 26630 5134 26682
rect 5186 26630 5198 26682
rect 5250 26630 5262 26682
rect 5314 26630 5326 26682
rect 5378 26630 5390 26682
rect 5442 26630 35854 26682
rect 35906 26630 35918 26682
rect 35970 26630 35982 26682
rect 36034 26630 36046 26682
rect 36098 26630 36110 26682
rect 36162 26630 66574 26682
rect 66626 26630 66638 26682
rect 66690 26630 66702 26682
rect 66754 26630 66766 26682
rect 66818 26630 66830 26682
rect 66882 26630 77924 26682
rect 2024 26608 77924 26630
rect 2024 26138 77924 26160
rect 2024 26086 5794 26138
rect 5846 26086 5858 26138
rect 5910 26086 5922 26138
rect 5974 26086 5986 26138
rect 6038 26086 6050 26138
rect 6102 26086 36514 26138
rect 36566 26086 36578 26138
rect 36630 26086 36642 26138
rect 36694 26086 36706 26138
rect 36758 26086 36770 26138
rect 36822 26086 67234 26138
rect 67286 26086 67298 26138
rect 67350 26086 67362 26138
rect 67414 26086 67426 26138
rect 67478 26086 67490 26138
rect 67542 26086 77924 26138
rect 2024 26064 77924 26086
rect 2024 25594 77924 25616
rect 2024 25542 5134 25594
rect 5186 25542 5198 25594
rect 5250 25542 5262 25594
rect 5314 25542 5326 25594
rect 5378 25542 5390 25594
rect 5442 25542 35854 25594
rect 35906 25542 35918 25594
rect 35970 25542 35982 25594
rect 36034 25542 36046 25594
rect 36098 25542 36110 25594
rect 36162 25542 66574 25594
rect 66626 25542 66638 25594
rect 66690 25542 66702 25594
rect 66754 25542 66766 25594
rect 66818 25542 66830 25594
rect 66882 25542 77924 25594
rect 2024 25520 77924 25542
rect 2024 25050 77924 25072
rect 2024 24998 5794 25050
rect 5846 24998 5858 25050
rect 5910 24998 5922 25050
rect 5974 24998 5986 25050
rect 6038 24998 6050 25050
rect 6102 24998 36514 25050
rect 36566 24998 36578 25050
rect 36630 24998 36642 25050
rect 36694 24998 36706 25050
rect 36758 24998 36770 25050
rect 36822 24998 67234 25050
rect 67286 24998 67298 25050
rect 67350 24998 67362 25050
rect 67414 24998 67426 25050
rect 67478 24998 67490 25050
rect 67542 24998 77924 25050
rect 2024 24976 77924 24998
rect 2024 24506 77924 24528
rect 2024 24454 5134 24506
rect 5186 24454 5198 24506
rect 5250 24454 5262 24506
rect 5314 24454 5326 24506
rect 5378 24454 5390 24506
rect 5442 24454 35854 24506
rect 35906 24454 35918 24506
rect 35970 24454 35982 24506
rect 36034 24454 36046 24506
rect 36098 24454 36110 24506
rect 36162 24454 66574 24506
rect 66626 24454 66638 24506
rect 66690 24454 66702 24506
rect 66754 24454 66766 24506
rect 66818 24454 66830 24506
rect 66882 24454 77924 24506
rect 2024 24432 77924 24454
rect 21910 24148 21916 24200
rect 21968 24188 21974 24200
rect 33318 24188 33324 24200
rect 21968 24160 33324 24188
rect 21968 24148 21974 24160
rect 33318 24148 33324 24160
rect 33376 24148 33382 24200
rect 3510 24080 3516 24132
rect 3568 24120 3574 24132
rect 35342 24120 35348 24132
rect 3568 24092 35348 24120
rect 3568 24080 3574 24092
rect 35342 24080 35348 24092
rect 35400 24080 35406 24132
rect 2024 23962 77924 23984
rect 2024 23910 5794 23962
rect 5846 23910 5858 23962
rect 5910 23910 5922 23962
rect 5974 23910 5986 23962
rect 6038 23910 6050 23962
rect 6102 23910 36514 23962
rect 36566 23910 36578 23962
rect 36630 23910 36642 23962
rect 36694 23910 36706 23962
rect 36758 23910 36770 23962
rect 36822 23910 67234 23962
rect 67286 23910 67298 23962
rect 67350 23910 67362 23962
rect 67414 23910 67426 23962
rect 67478 23910 67490 23962
rect 67542 23910 77924 23962
rect 2024 23888 77924 23910
rect 2024 23418 77924 23440
rect 2024 23366 5134 23418
rect 5186 23366 5198 23418
rect 5250 23366 5262 23418
rect 5314 23366 5326 23418
rect 5378 23366 5390 23418
rect 5442 23366 35854 23418
rect 35906 23366 35918 23418
rect 35970 23366 35982 23418
rect 36034 23366 36046 23418
rect 36098 23366 36110 23418
rect 36162 23366 66574 23418
rect 66626 23366 66638 23418
rect 66690 23366 66702 23418
rect 66754 23366 66766 23418
rect 66818 23366 66830 23418
rect 66882 23366 77924 23418
rect 2024 23344 77924 23366
rect 2024 22874 77924 22896
rect 2024 22822 5794 22874
rect 5846 22822 5858 22874
rect 5910 22822 5922 22874
rect 5974 22822 5986 22874
rect 6038 22822 6050 22874
rect 6102 22822 36514 22874
rect 36566 22822 36578 22874
rect 36630 22822 36642 22874
rect 36694 22822 36706 22874
rect 36758 22822 36770 22874
rect 36822 22822 67234 22874
rect 67286 22822 67298 22874
rect 67350 22822 67362 22874
rect 67414 22822 67426 22874
rect 67478 22822 67490 22874
rect 67542 22822 77924 22874
rect 2024 22800 77924 22822
rect 2024 22330 77924 22352
rect 2024 22278 5134 22330
rect 5186 22278 5198 22330
rect 5250 22278 5262 22330
rect 5314 22278 5326 22330
rect 5378 22278 5390 22330
rect 5442 22278 35854 22330
rect 35906 22278 35918 22330
rect 35970 22278 35982 22330
rect 36034 22278 36046 22330
rect 36098 22278 36110 22330
rect 36162 22278 66574 22330
rect 66626 22278 66638 22330
rect 66690 22278 66702 22330
rect 66754 22278 66766 22330
rect 66818 22278 66830 22330
rect 66882 22278 77924 22330
rect 2024 22256 77924 22278
rect 2024 21786 77924 21808
rect 2024 21734 5794 21786
rect 5846 21734 5858 21786
rect 5910 21734 5922 21786
rect 5974 21734 5986 21786
rect 6038 21734 6050 21786
rect 6102 21734 36514 21786
rect 36566 21734 36578 21786
rect 36630 21734 36642 21786
rect 36694 21734 36706 21786
rect 36758 21734 36770 21786
rect 36822 21734 67234 21786
rect 67286 21734 67298 21786
rect 67350 21734 67362 21786
rect 67414 21734 67426 21786
rect 67478 21734 67490 21786
rect 67542 21734 77924 21786
rect 2024 21712 77924 21734
rect 28718 21360 28724 21412
rect 28776 21400 28782 21412
rect 39114 21400 39120 21412
rect 28776 21372 39120 21400
rect 28776 21360 28782 21372
rect 39114 21360 39120 21372
rect 39172 21360 39178 21412
rect 2024 21242 77924 21264
rect 2024 21190 5134 21242
rect 5186 21190 5198 21242
rect 5250 21190 5262 21242
rect 5314 21190 5326 21242
rect 5378 21190 5390 21242
rect 5442 21190 35854 21242
rect 35906 21190 35918 21242
rect 35970 21190 35982 21242
rect 36034 21190 36046 21242
rect 36098 21190 36110 21242
rect 36162 21190 66574 21242
rect 66626 21190 66638 21242
rect 66690 21190 66702 21242
rect 66754 21190 66766 21242
rect 66818 21190 66830 21242
rect 66882 21190 77924 21242
rect 2024 21168 77924 21190
rect 2024 20698 77924 20720
rect 2024 20646 5794 20698
rect 5846 20646 5858 20698
rect 5910 20646 5922 20698
rect 5974 20646 5986 20698
rect 6038 20646 6050 20698
rect 6102 20646 36514 20698
rect 36566 20646 36578 20698
rect 36630 20646 36642 20698
rect 36694 20646 36706 20698
rect 36758 20646 36770 20698
rect 36822 20646 67234 20698
rect 67286 20646 67298 20698
rect 67350 20646 67362 20698
rect 67414 20646 67426 20698
rect 67478 20646 67490 20698
rect 67542 20646 77924 20698
rect 2024 20624 77924 20646
rect 2024 20154 77924 20176
rect 2024 20102 5134 20154
rect 5186 20102 5198 20154
rect 5250 20102 5262 20154
rect 5314 20102 5326 20154
rect 5378 20102 5390 20154
rect 5442 20102 35854 20154
rect 35906 20102 35918 20154
rect 35970 20102 35982 20154
rect 36034 20102 36046 20154
rect 36098 20102 36110 20154
rect 36162 20102 66574 20154
rect 66626 20102 66638 20154
rect 66690 20102 66702 20154
rect 66754 20102 66766 20154
rect 66818 20102 66830 20154
rect 66882 20102 77924 20154
rect 2024 20080 77924 20102
rect 2024 19610 77924 19632
rect 2024 19558 5794 19610
rect 5846 19558 5858 19610
rect 5910 19558 5922 19610
rect 5974 19558 5986 19610
rect 6038 19558 6050 19610
rect 6102 19558 36514 19610
rect 36566 19558 36578 19610
rect 36630 19558 36642 19610
rect 36694 19558 36706 19610
rect 36758 19558 36770 19610
rect 36822 19558 67234 19610
rect 67286 19558 67298 19610
rect 67350 19558 67362 19610
rect 67414 19558 67426 19610
rect 67478 19558 67490 19610
rect 67542 19558 77924 19610
rect 2024 19536 77924 19558
rect 2024 19066 77924 19088
rect 2024 19014 5134 19066
rect 5186 19014 5198 19066
rect 5250 19014 5262 19066
rect 5314 19014 5326 19066
rect 5378 19014 5390 19066
rect 5442 19014 35854 19066
rect 35906 19014 35918 19066
rect 35970 19014 35982 19066
rect 36034 19014 36046 19066
rect 36098 19014 36110 19066
rect 36162 19014 66574 19066
rect 66626 19014 66638 19066
rect 66690 19014 66702 19066
rect 66754 19014 66766 19066
rect 66818 19014 66830 19066
rect 66882 19014 77924 19066
rect 2024 18992 77924 19014
rect 2024 18522 77924 18544
rect 2024 18470 5794 18522
rect 5846 18470 5858 18522
rect 5910 18470 5922 18522
rect 5974 18470 5986 18522
rect 6038 18470 6050 18522
rect 6102 18470 36514 18522
rect 36566 18470 36578 18522
rect 36630 18470 36642 18522
rect 36694 18470 36706 18522
rect 36758 18470 36770 18522
rect 36822 18470 67234 18522
rect 67286 18470 67298 18522
rect 67350 18470 67362 18522
rect 67414 18470 67426 18522
rect 67478 18470 67490 18522
rect 67542 18470 77924 18522
rect 2024 18448 77924 18470
rect 2024 17978 77924 18000
rect 2024 17926 5134 17978
rect 5186 17926 5198 17978
rect 5250 17926 5262 17978
rect 5314 17926 5326 17978
rect 5378 17926 5390 17978
rect 5442 17926 35854 17978
rect 35906 17926 35918 17978
rect 35970 17926 35982 17978
rect 36034 17926 36046 17978
rect 36098 17926 36110 17978
rect 36162 17926 66574 17978
rect 66626 17926 66638 17978
rect 66690 17926 66702 17978
rect 66754 17926 66766 17978
rect 66818 17926 66830 17978
rect 66882 17926 77924 17978
rect 2024 17904 77924 17926
rect 2024 17434 77924 17456
rect 2024 17382 5794 17434
rect 5846 17382 5858 17434
rect 5910 17382 5922 17434
rect 5974 17382 5986 17434
rect 6038 17382 6050 17434
rect 6102 17382 36514 17434
rect 36566 17382 36578 17434
rect 36630 17382 36642 17434
rect 36694 17382 36706 17434
rect 36758 17382 36770 17434
rect 36822 17382 67234 17434
rect 67286 17382 67298 17434
rect 67350 17382 67362 17434
rect 67414 17382 67426 17434
rect 67478 17382 67490 17434
rect 67542 17382 77924 17434
rect 2024 17360 77924 17382
rect 2024 16890 77924 16912
rect 2024 16838 5134 16890
rect 5186 16838 5198 16890
rect 5250 16838 5262 16890
rect 5314 16838 5326 16890
rect 5378 16838 5390 16890
rect 5442 16838 35854 16890
rect 35906 16838 35918 16890
rect 35970 16838 35982 16890
rect 36034 16838 36046 16890
rect 36098 16838 36110 16890
rect 36162 16838 66574 16890
rect 66626 16838 66638 16890
rect 66690 16838 66702 16890
rect 66754 16838 66766 16890
rect 66818 16838 66830 16890
rect 66882 16838 77924 16890
rect 2024 16816 77924 16838
rect 2024 16346 77924 16368
rect 2024 16294 5794 16346
rect 5846 16294 5858 16346
rect 5910 16294 5922 16346
rect 5974 16294 5986 16346
rect 6038 16294 6050 16346
rect 6102 16294 36514 16346
rect 36566 16294 36578 16346
rect 36630 16294 36642 16346
rect 36694 16294 36706 16346
rect 36758 16294 36770 16346
rect 36822 16294 67234 16346
rect 67286 16294 67298 16346
rect 67350 16294 67362 16346
rect 67414 16294 67426 16346
rect 67478 16294 67490 16346
rect 67542 16294 77924 16346
rect 2024 16272 77924 16294
rect 2024 15802 77924 15824
rect 2024 15750 5134 15802
rect 5186 15750 5198 15802
rect 5250 15750 5262 15802
rect 5314 15750 5326 15802
rect 5378 15750 5390 15802
rect 5442 15750 35854 15802
rect 35906 15750 35918 15802
rect 35970 15750 35982 15802
rect 36034 15750 36046 15802
rect 36098 15750 36110 15802
rect 36162 15750 66574 15802
rect 66626 15750 66638 15802
rect 66690 15750 66702 15802
rect 66754 15750 66766 15802
rect 66818 15750 66830 15802
rect 66882 15750 77924 15802
rect 2024 15728 77924 15750
rect 2024 15258 77924 15280
rect 2024 15206 5794 15258
rect 5846 15206 5858 15258
rect 5910 15206 5922 15258
rect 5974 15206 5986 15258
rect 6038 15206 6050 15258
rect 6102 15206 36514 15258
rect 36566 15206 36578 15258
rect 36630 15206 36642 15258
rect 36694 15206 36706 15258
rect 36758 15206 36770 15258
rect 36822 15206 67234 15258
rect 67286 15206 67298 15258
rect 67350 15206 67362 15258
rect 67414 15206 67426 15258
rect 67478 15206 67490 15258
rect 67542 15206 77924 15258
rect 2024 15184 77924 15206
rect 2024 14714 77924 14736
rect 2024 14662 5134 14714
rect 5186 14662 5198 14714
rect 5250 14662 5262 14714
rect 5314 14662 5326 14714
rect 5378 14662 5390 14714
rect 5442 14662 35854 14714
rect 35906 14662 35918 14714
rect 35970 14662 35982 14714
rect 36034 14662 36046 14714
rect 36098 14662 36110 14714
rect 36162 14662 66574 14714
rect 66626 14662 66638 14714
rect 66690 14662 66702 14714
rect 66754 14662 66766 14714
rect 66818 14662 66830 14714
rect 66882 14662 77924 14714
rect 2024 14640 77924 14662
rect 27430 14492 27436 14544
rect 27488 14532 27494 14544
rect 43346 14532 43352 14544
rect 27488 14504 43352 14532
rect 27488 14492 27494 14504
rect 43346 14492 43352 14504
rect 43404 14492 43410 14544
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 58802 14464 58808 14476
rect 24912 14436 58808 14464
rect 24912 14424 24918 14436
rect 58802 14424 58808 14436
rect 58860 14424 58866 14476
rect 2024 14170 77924 14192
rect 2024 14118 5794 14170
rect 5846 14118 5858 14170
rect 5910 14118 5922 14170
rect 5974 14118 5986 14170
rect 6038 14118 6050 14170
rect 6102 14118 36514 14170
rect 36566 14118 36578 14170
rect 36630 14118 36642 14170
rect 36694 14118 36706 14170
rect 36758 14118 36770 14170
rect 36822 14118 67234 14170
rect 67286 14118 67298 14170
rect 67350 14118 67362 14170
rect 67414 14118 67426 14170
rect 67478 14118 67490 14170
rect 67542 14118 77924 14170
rect 2024 14096 77924 14118
rect 2024 13626 77924 13648
rect 2024 13574 5134 13626
rect 5186 13574 5198 13626
rect 5250 13574 5262 13626
rect 5314 13574 5326 13626
rect 5378 13574 5390 13626
rect 5442 13574 35854 13626
rect 35906 13574 35918 13626
rect 35970 13574 35982 13626
rect 36034 13574 36046 13626
rect 36098 13574 36110 13626
rect 36162 13574 66574 13626
rect 66626 13574 66638 13626
rect 66690 13574 66702 13626
rect 66754 13574 66766 13626
rect 66818 13574 66830 13626
rect 66882 13574 77924 13626
rect 2024 13552 77924 13574
rect 2024 13082 77924 13104
rect 2024 13030 5794 13082
rect 5846 13030 5858 13082
rect 5910 13030 5922 13082
rect 5974 13030 5986 13082
rect 6038 13030 6050 13082
rect 6102 13030 36514 13082
rect 36566 13030 36578 13082
rect 36630 13030 36642 13082
rect 36694 13030 36706 13082
rect 36758 13030 36770 13082
rect 36822 13030 67234 13082
rect 67286 13030 67298 13082
rect 67350 13030 67362 13082
rect 67414 13030 67426 13082
rect 67478 13030 67490 13082
rect 67542 13030 77924 13082
rect 2024 13008 77924 13030
rect 2024 12538 77924 12560
rect 2024 12486 5134 12538
rect 5186 12486 5198 12538
rect 5250 12486 5262 12538
rect 5314 12486 5326 12538
rect 5378 12486 5390 12538
rect 5442 12486 35854 12538
rect 35906 12486 35918 12538
rect 35970 12486 35982 12538
rect 36034 12486 36046 12538
rect 36098 12486 36110 12538
rect 36162 12486 66574 12538
rect 66626 12486 66638 12538
rect 66690 12486 66702 12538
rect 66754 12486 66766 12538
rect 66818 12486 66830 12538
rect 66882 12486 77924 12538
rect 2024 12464 77924 12486
rect 28626 12180 28632 12232
rect 28684 12220 28690 12232
rect 31018 12220 31024 12232
rect 28684 12192 31024 12220
rect 28684 12180 28690 12192
rect 31018 12180 31024 12192
rect 31076 12180 31082 12232
rect 16574 12112 16580 12164
rect 16632 12152 16638 12164
rect 30006 12152 30012 12164
rect 16632 12124 30012 12152
rect 16632 12112 16638 12124
rect 30006 12112 30012 12124
rect 30064 12112 30070 12164
rect 17586 12044 17592 12096
rect 17644 12084 17650 12096
rect 25314 12084 25320 12096
rect 17644 12056 25320 12084
rect 17644 12044 17650 12056
rect 25314 12044 25320 12056
rect 25372 12044 25378 12096
rect 28902 12044 28908 12096
rect 28960 12084 28966 12096
rect 30558 12084 30564 12096
rect 28960 12056 30564 12084
rect 28960 12044 28966 12056
rect 30558 12044 30564 12056
rect 30616 12044 30622 12096
rect 2024 11994 77924 12016
rect 2024 11942 5794 11994
rect 5846 11942 5858 11994
rect 5910 11942 5922 11994
rect 5974 11942 5986 11994
rect 6038 11942 6050 11994
rect 6102 11942 36514 11994
rect 36566 11942 36578 11994
rect 36630 11942 36642 11994
rect 36694 11942 36706 11994
rect 36758 11942 36770 11994
rect 36822 11942 67234 11994
rect 67286 11942 67298 11994
rect 67350 11942 67362 11994
rect 67414 11942 67426 11994
rect 67478 11942 67490 11994
rect 67542 11942 77924 11994
rect 2024 11920 77924 11942
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 22097 11883 22155 11889
rect 22097 11880 22109 11883
rect 9272 11852 22109 11880
rect 9272 11840 9278 11852
rect 22097 11849 22109 11852
rect 22143 11880 22155 11883
rect 22462 11880 22468 11892
rect 22143 11852 22468 11880
rect 22143 11849 22155 11852
rect 22097 11843 22155 11849
rect 22462 11840 22468 11852
rect 22520 11840 22526 11892
rect 26221 11883 26279 11889
rect 26221 11849 26233 11883
rect 26267 11880 26279 11883
rect 27246 11880 27252 11892
rect 26267 11852 27252 11880
rect 26267 11849 26279 11852
rect 26221 11843 26279 11849
rect 27246 11840 27252 11852
rect 27304 11840 27310 11892
rect 27430 11840 27436 11892
rect 27488 11880 27494 11892
rect 28813 11883 28871 11889
rect 28813 11880 28825 11883
rect 27488 11852 28825 11880
rect 27488 11840 27494 11852
rect 28813 11849 28825 11852
rect 28859 11880 28871 11883
rect 28902 11880 28908 11892
rect 28859 11852 28908 11880
rect 28859 11849 28871 11852
rect 28813 11843 28871 11849
rect 28902 11840 28908 11852
rect 28960 11840 28966 11892
rect 29089 11883 29147 11889
rect 29089 11849 29101 11883
rect 29135 11880 29147 11883
rect 32122 11880 32128 11892
rect 29135 11852 32128 11880
rect 29135 11849 29147 11852
rect 29089 11843 29147 11849
rect 32122 11840 32128 11852
rect 32180 11840 32186 11892
rect 8478 11772 8484 11824
rect 8536 11812 8542 11824
rect 22002 11812 22008 11824
rect 8536 11784 22008 11812
rect 8536 11772 8542 11784
rect 22002 11772 22008 11784
rect 22060 11772 22066 11824
rect 22186 11772 22192 11824
rect 22244 11812 22250 11824
rect 23753 11815 23811 11821
rect 23753 11812 23765 11815
rect 22244 11784 23765 11812
rect 22244 11772 22250 11784
rect 23753 11781 23765 11784
rect 23799 11812 23811 11815
rect 23934 11812 23940 11824
rect 23799 11784 23940 11812
rect 23799 11781 23811 11784
rect 23753 11775 23811 11781
rect 23934 11772 23940 11784
rect 23992 11772 23998 11824
rect 26418 11772 26424 11824
rect 26476 11772 26482 11824
rect 26896 11784 29960 11812
rect 22462 11704 22468 11756
rect 22520 11704 22526 11756
rect 23661 11747 23719 11753
rect 23661 11713 23673 11747
rect 23707 11713 23719 11747
rect 23661 11707 23719 11713
rect 12618 11636 12624 11688
rect 12676 11676 12682 11688
rect 23293 11679 23351 11685
rect 23293 11676 23305 11679
rect 12676 11648 23305 11676
rect 12676 11636 12682 11648
rect 23293 11645 23305 11648
rect 23339 11676 23351 11679
rect 23676 11676 23704 11707
rect 24302 11704 24308 11756
rect 24360 11744 24366 11756
rect 24765 11747 24823 11753
rect 24765 11744 24777 11747
rect 24360 11716 24777 11744
rect 24360 11704 24366 11716
rect 24765 11713 24777 11716
rect 24811 11713 24823 11747
rect 24765 11707 24823 11713
rect 25133 11747 25191 11753
rect 25133 11713 25145 11747
rect 25179 11744 25191 11747
rect 26896 11744 26924 11784
rect 25179 11716 26924 11744
rect 26973 11747 27031 11753
rect 25179 11713 25191 11716
rect 25133 11707 25191 11713
rect 26973 11713 26985 11747
rect 27019 11713 27031 11747
rect 26973 11707 27031 11713
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 27249 11747 27307 11753
rect 27249 11713 27261 11747
rect 27295 11744 27307 11747
rect 27890 11744 27896 11756
rect 27295 11716 27896 11744
rect 27295 11713 27307 11716
rect 27249 11707 27307 11713
rect 23339 11648 23704 11676
rect 23339 11645 23351 11648
rect 23293 11639 23351 11645
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 26878 11608 26884 11620
rect 15068 11580 26884 11608
rect 15068 11568 15074 11580
rect 26878 11568 26884 11580
rect 26936 11568 26942 11620
rect 26988 11608 27016 11707
rect 27172 11676 27200 11707
rect 27890 11704 27896 11716
rect 27948 11704 27954 11756
rect 28626 11704 28632 11756
rect 28684 11704 28690 11756
rect 28889 11747 28947 11753
rect 28889 11744 28901 11747
rect 28828 11716 28901 11744
rect 27430 11676 27436 11688
rect 27172 11648 27436 11676
rect 27430 11636 27436 11648
rect 27488 11636 27494 11688
rect 28442 11636 28448 11688
rect 28500 11636 28506 11688
rect 28644 11608 28672 11704
rect 28718 11636 28724 11688
rect 28776 11676 28782 11688
rect 28828 11676 28856 11716
rect 28889 11713 28901 11716
rect 28935 11713 28947 11747
rect 28889 11707 28947 11713
rect 28997 11747 29055 11753
rect 28997 11713 29009 11747
rect 29043 11744 29055 11747
rect 29086 11744 29092 11756
rect 29043 11716 29092 11744
rect 29043 11713 29055 11716
rect 28997 11707 29055 11713
rect 29086 11704 29092 11716
rect 29144 11704 29150 11756
rect 29178 11704 29184 11756
rect 29236 11744 29242 11756
rect 29549 11747 29607 11753
rect 29549 11744 29561 11747
rect 29236 11716 29561 11744
rect 29236 11704 29242 11716
rect 29549 11713 29561 11716
rect 29595 11713 29607 11747
rect 29549 11707 29607 11713
rect 28776 11648 28856 11676
rect 29459 11679 29517 11685
rect 28776 11636 28782 11648
rect 29459 11645 29471 11679
rect 29505 11645 29517 11679
rect 29932 11676 29960 11784
rect 30006 11772 30012 11824
rect 30064 11772 30070 11824
rect 30558 11772 30564 11824
rect 30616 11772 30622 11824
rect 33226 11772 33232 11824
rect 33284 11812 33290 11824
rect 33870 11812 33876 11824
rect 33284 11784 33876 11812
rect 33284 11772 33290 11784
rect 33870 11772 33876 11784
rect 33928 11772 33934 11824
rect 30466 11704 30472 11756
rect 30524 11704 30530 11756
rect 30745 11747 30803 11753
rect 30745 11713 30757 11747
rect 30791 11744 30803 11747
rect 31018 11744 31024 11756
rect 30791 11716 31024 11744
rect 30791 11713 30803 11716
rect 30745 11707 30803 11713
rect 31018 11704 31024 11716
rect 31076 11704 31082 11756
rect 33318 11704 33324 11756
rect 33376 11704 33382 11756
rect 33413 11747 33471 11753
rect 33413 11713 33425 11747
rect 33459 11744 33471 11747
rect 33962 11744 33968 11756
rect 33459 11716 33968 11744
rect 33459 11713 33471 11716
rect 33413 11707 33471 11713
rect 33962 11704 33968 11716
rect 34020 11704 34026 11756
rect 30650 11676 30656 11688
rect 29932 11648 30656 11676
rect 29459 11639 29517 11645
rect 26988 11580 28672 11608
rect 28902 11568 28908 11620
rect 28960 11608 28966 11620
rect 29472 11608 29500 11639
rect 30650 11636 30656 11648
rect 30708 11636 30714 11688
rect 33226 11636 33232 11688
rect 33284 11676 33290 11688
rect 33336 11676 33364 11704
rect 33284 11648 33364 11676
rect 33284 11636 33290 11648
rect 28960 11580 29500 11608
rect 28960 11568 28966 11580
rect 33042 11568 33048 11620
rect 33100 11568 33106 11620
rect 22278 11500 22284 11552
rect 22336 11500 22342 11552
rect 22738 11500 22744 11552
rect 22796 11500 22802 11552
rect 23474 11500 23480 11552
rect 23532 11500 23538 11552
rect 24210 11500 24216 11552
rect 24268 11540 24274 11552
rect 24670 11540 24676 11552
rect 24268 11512 24676 11540
rect 24268 11500 24274 11512
rect 24670 11500 24676 11512
rect 24728 11500 24734 11552
rect 25222 11500 25228 11552
rect 25280 11500 25286 11552
rect 25958 11500 25964 11552
rect 26016 11540 26022 11552
rect 26053 11543 26111 11549
rect 26053 11540 26065 11543
rect 26016 11512 26065 11540
rect 26016 11500 26022 11512
rect 26053 11509 26065 11512
rect 26099 11509 26111 11543
rect 26053 11503 26111 11509
rect 26237 11543 26295 11549
rect 26237 11509 26249 11543
rect 26283 11540 26295 11543
rect 26510 11540 26516 11552
rect 26283 11512 26516 11540
rect 26283 11509 26295 11512
rect 26237 11503 26295 11509
rect 26510 11500 26516 11512
rect 26568 11500 26574 11552
rect 26602 11500 26608 11552
rect 26660 11540 26666 11552
rect 26789 11543 26847 11549
rect 26789 11540 26801 11543
rect 26660 11512 26801 11540
rect 26660 11500 26666 11512
rect 26789 11509 26801 11512
rect 26835 11509 26847 11543
rect 26789 11503 26847 11509
rect 28350 11500 28356 11552
rect 28408 11540 28414 11552
rect 29273 11543 29331 11549
rect 29273 11540 29285 11543
rect 28408 11512 29285 11540
rect 28408 11500 28414 11512
rect 29273 11509 29285 11512
rect 29319 11509 29331 11543
rect 29273 11503 29331 11509
rect 29362 11500 29368 11552
rect 29420 11540 29426 11552
rect 30101 11543 30159 11549
rect 30101 11540 30113 11543
rect 29420 11512 30113 11540
rect 29420 11500 29426 11512
rect 30101 11509 30113 11512
rect 30147 11509 30159 11543
rect 30101 11503 30159 11509
rect 30282 11500 30288 11552
rect 30340 11540 30346 11552
rect 30929 11543 30987 11549
rect 30929 11540 30941 11543
rect 30340 11512 30941 11540
rect 30340 11500 30346 11512
rect 30929 11509 30941 11512
rect 30975 11509 30987 11543
rect 30929 11503 30987 11509
rect 33597 11543 33655 11549
rect 33597 11509 33609 11543
rect 33643 11540 33655 11543
rect 35618 11540 35624 11552
rect 33643 11512 35624 11540
rect 33643 11509 33655 11512
rect 33597 11503 33655 11509
rect 35618 11500 35624 11512
rect 35676 11500 35682 11552
rect 2024 11450 77924 11472
rect 2024 11398 5134 11450
rect 5186 11398 5198 11450
rect 5250 11398 5262 11450
rect 5314 11398 5326 11450
rect 5378 11398 5390 11450
rect 5442 11398 35854 11450
rect 35906 11398 35918 11450
rect 35970 11398 35982 11450
rect 36034 11398 36046 11450
rect 36098 11398 36110 11450
rect 36162 11398 66574 11450
rect 66626 11398 66638 11450
rect 66690 11398 66702 11450
rect 66754 11398 66766 11450
rect 66818 11398 66830 11450
rect 66882 11398 77924 11450
rect 2024 11376 77924 11398
rect 14550 11296 14556 11348
rect 14608 11336 14614 11348
rect 22278 11336 22284 11348
rect 14608 11308 22284 11336
rect 14608 11296 14614 11308
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22646 11296 22652 11348
rect 22704 11336 22710 11348
rect 22925 11339 22983 11345
rect 22925 11336 22937 11339
rect 22704 11308 22937 11336
rect 22704 11296 22710 11308
rect 22925 11305 22937 11308
rect 22971 11305 22983 11339
rect 22925 11299 22983 11305
rect 23290 11296 23296 11348
rect 23348 11336 23354 11348
rect 24854 11336 24860 11348
rect 23348 11308 24860 11336
rect 23348 11296 23354 11308
rect 24854 11296 24860 11308
rect 24912 11296 24918 11348
rect 25314 11296 25320 11348
rect 25372 11296 25378 11348
rect 26050 11296 26056 11348
rect 26108 11336 26114 11348
rect 26108 11308 26832 11336
rect 26108 11296 26114 11308
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 23474 11268 23480 11280
rect 16264 11240 23480 11268
rect 16264 11228 16270 11240
rect 23474 11228 23480 11240
rect 23532 11228 23538 11280
rect 12342 11160 12348 11212
rect 12400 11200 12406 11212
rect 22462 11200 22468 11212
rect 12400 11172 22468 11200
rect 12400 11160 12406 11172
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 22738 11200 22744 11212
rect 22664 11172 22744 11200
rect 21726 11092 21732 11144
rect 21784 11092 21790 11144
rect 22557 11135 22615 11141
rect 22557 11101 22569 11135
rect 22603 11126 22615 11135
rect 22664 11126 22692 11172
rect 22738 11160 22744 11172
rect 22796 11160 22802 11212
rect 23934 11160 23940 11212
rect 23992 11160 23998 11212
rect 24210 11160 24216 11212
rect 24268 11160 24274 11212
rect 24397 11203 24455 11209
rect 24397 11169 24409 11203
rect 24443 11200 24455 11203
rect 24443 11172 24900 11200
rect 24443 11169 24455 11172
rect 24397 11163 24455 11169
rect 24872 11144 24900 11172
rect 25222 11160 25228 11212
rect 25280 11200 25286 11212
rect 25869 11203 25927 11209
rect 25869 11200 25881 11203
rect 25280 11172 25881 11200
rect 25280 11160 25286 11172
rect 25869 11169 25881 11172
rect 25915 11169 25927 11203
rect 25869 11163 25927 11169
rect 26234 11160 26240 11212
rect 26292 11160 26298 11212
rect 26804 11209 26832 11308
rect 28810 11296 28816 11348
rect 28868 11296 28874 11348
rect 31665 11339 31723 11345
rect 31665 11305 31677 11339
rect 31711 11336 31723 11339
rect 38378 11336 38384 11348
rect 31711 11308 38384 11336
rect 31711 11305 31723 11308
rect 31665 11299 31723 11305
rect 38378 11296 38384 11308
rect 38436 11296 38442 11348
rect 26878 11228 26884 11280
rect 26936 11268 26942 11280
rect 33045 11271 33103 11277
rect 33045 11268 33057 11271
rect 26936 11240 33057 11268
rect 26936 11228 26942 11240
rect 33045 11237 33057 11240
rect 33091 11237 33103 11271
rect 33045 11231 33103 11237
rect 33226 11228 33232 11280
rect 33284 11268 33290 11280
rect 33284 11240 34744 11268
rect 33284 11228 33290 11240
rect 26789 11203 26847 11209
rect 26789 11169 26801 11203
rect 26835 11169 26847 11203
rect 26789 11163 26847 11169
rect 26896 11172 28580 11200
rect 22603 11101 22692 11126
rect 22557 11098 22692 11101
rect 22557 11095 22615 11098
rect 24670 11092 24676 11144
rect 24728 11092 24734 11144
rect 24854 11092 24860 11144
rect 24912 11092 24918 11144
rect 24946 11092 24952 11144
rect 25004 11092 25010 11144
rect 25038 11092 25044 11144
rect 25096 11132 25102 11144
rect 26896 11132 26924 11172
rect 25096 11104 26924 11132
rect 25096 11092 25102 11104
rect 26970 11092 26976 11144
rect 27028 11132 27034 11144
rect 27709 11135 27767 11141
rect 27709 11132 27721 11135
rect 27028 11104 27721 11132
rect 27028 11092 27034 11104
rect 27709 11101 27721 11104
rect 27755 11101 27767 11135
rect 27709 11095 27767 11101
rect 28442 11092 28448 11144
rect 28500 11092 28506 11144
rect 28552 11132 28580 11172
rect 29178 11160 29184 11212
rect 29236 11200 29242 11212
rect 30101 11203 30159 11209
rect 30101 11200 30113 11203
rect 29236 11172 30113 11200
rect 29236 11160 29242 11172
rect 30101 11169 30113 11172
rect 30147 11169 30159 11203
rect 30101 11163 30159 11169
rect 30190 11160 30196 11212
rect 30248 11200 30254 11212
rect 32217 11203 32275 11209
rect 32217 11200 32229 11203
rect 30248 11172 32229 11200
rect 30248 11160 30254 11172
rect 32217 11169 32229 11172
rect 32263 11169 32275 11203
rect 32217 11163 32275 11169
rect 32582 11160 32588 11212
rect 32640 11200 32646 11212
rect 33781 11203 33839 11209
rect 33781 11200 33793 11203
rect 32640 11172 33793 11200
rect 32640 11160 32646 11172
rect 33781 11169 33793 11172
rect 33827 11169 33839 11203
rect 34149 11203 34207 11209
rect 34149 11200 34161 11203
rect 33781 11163 33839 11169
rect 33888 11172 34161 11200
rect 29365 11135 29423 11141
rect 29365 11132 29377 11135
rect 28552 11104 29377 11132
rect 29365 11101 29377 11104
rect 29411 11101 29423 11135
rect 29365 11095 29423 11101
rect 31386 11092 31392 11144
rect 31444 11092 31450 11144
rect 33410 11092 33416 11144
rect 33468 11132 33474 11144
rect 33597 11135 33655 11141
rect 33597 11132 33609 11135
rect 33468 11104 33609 11132
rect 33468 11092 33474 11104
rect 33597 11101 33609 11104
rect 33643 11101 33655 11135
rect 33888 11132 33916 11172
rect 34149 11169 34161 11172
rect 34195 11200 34207 11203
rect 34425 11203 34483 11209
rect 34425 11200 34437 11203
rect 34195 11172 34437 11200
rect 34195 11169 34207 11172
rect 34149 11163 34207 11169
rect 34425 11169 34437 11172
rect 34471 11169 34483 11203
rect 34425 11163 34483 11169
rect 34716 11200 34744 11240
rect 35710 11200 35716 11212
rect 34716 11172 35716 11200
rect 33597 11095 33655 11101
rect 33704 11104 33916 11132
rect 21818 11024 21824 11076
rect 21876 11024 21882 11076
rect 22370 11024 22376 11076
rect 22428 11024 22434 11076
rect 22664 11036 23060 11064
rect 17678 10956 17684 11008
rect 17736 10996 17742 11008
rect 22664 10996 22692 11036
rect 17736 10968 22692 10996
rect 17736 10956 17742 10968
rect 22738 10956 22744 11008
rect 22796 10956 22802 11008
rect 23032 10996 23060 11036
rect 23198 11024 23204 11076
rect 23256 11024 23262 11076
rect 23382 11024 23388 11076
rect 23440 11024 23446 11076
rect 23474 11024 23480 11076
rect 23532 11064 23538 11076
rect 24489 11067 24547 11073
rect 24489 11064 24501 11067
rect 23532 11036 24501 11064
rect 23532 11024 23538 11036
rect 24489 11033 24501 11036
rect 24535 11033 24547 11067
rect 24489 11027 24547 11033
rect 26878 11024 26884 11076
rect 26936 11064 26942 11076
rect 27893 11067 27951 11073
rect 27893 11064 27905 11067
rect 26936 11036 27905 11064
rect 26936 11024 26942 11036
rect 27893 11033 27905 11036
rect 27939 11033 27951 11067
rect 27893 11027 27951 11033
rect 29546 11024 29552 11076
rect 29604 11024 29610 11076
rect 30742 11024 30748 11076
rect 30800 11024 30806 11076
rect 33042 11024 33048 11076
rect 33100 11064 33106 11076
rect 33704 11064 33732 11104
rect 33962 11092 33968 11144
rect 34020 11092 34026 11144
rect 34057 11135 34115 11141
rect 34057 11101 34069 11135
rect 34103 11132 34115 11135
rect 34241 11135 34299 11141
rect 34103 11104 34137 11132
rect 34103 11101 34115 11104
rect 34057 11095 34115 11101
rect 34241 11101 34253 11135
rect 34287 11132 34299 11135
rect 34514 11132 34520 11144
rect 34287 11104 34520 11132
rect 34287 11101 34299 11104
rect 34241 11095 34299 11101
rect 33100 11036 33732 11064
rect 33100 11024 33106 11036
rect 33870 11024 33876 11076
rect 33928 11064 33934 11076
rect 34072 11064 34100 11095
rect 34514 11092 34520 11104
rect 34572 11092 34578 11144
rect 34716 11141 34744 11172
rect 35710 11160 35716 11172
rect 35768 11160 35774 11212
rect 34701 11135 34759 11141
rect 34701 11101 34713 11135
rect 34747 11101 34759 11135
rect 34701 11095 34759 11101
rect 34790 11092 34796 11144
rect 34848 11132 34854 11144
rect 37826 11132 37832 11144
rect 34848 11104 37832 11132
rect 34848 11092 34854 11104
rect 37826 11092 37832 11104
rect 37884 11092 37890 11144
rect 34609 11067 34667 11073
rect 34609 11064 34621 11067
rect 33928 11036 34621 11064
rect 33928 11024 33934 11036
rect 34609 11033 34621 11036
rect 34655 11033 34667 11067
rect 34609 11027 34667 11033
rect 34977 11067 35035 11073
rect 34977 11033 34989 11067
rect 35023 11064 35035 11067
rect 35250 11064 35256 11076
rect 35023 11036 35256 11064
rect 35023 11033 35035 11036
rect 34977 11027 35035 11033
rect 35250 11024 35256 11036
rect 35308 11024 35314 11076
rect 24026 10996 24032 11008
rect 23032 10968 24032 10996
rect 24026 10956 24032 10968
rect 24084 10956 24090 11008
rect 24118 10956 24124 11008
rect 24176 10996 24182 11008
rect 24946 10996 24952 11008
rect 24176 10968 24952 10996
rect 24176 10956 24182 10968
rect 24946 10956 24952 10968
rect 25004 10996 25010 11008
rect 25041 10999 25099 11005
rect 25041 10996 25053 10999
rect 25004 10968 25053 10996
rect 25004 10956 25010 10968
rect 25041 10965 25053 10968
rect 25087 10965 25099 10999
rect 25041 10959 25099 10965
rect 27157 10999 27215 11005
rect 27157 10965 27169 10999
rect 27203 10996 27215 10999
rect 27430 10996 27436 11008
rect 27203 10968 27436 10996
rect 27203 10965 27215 10968
rect 27157 10959 27215 10965
rect 27430 10956 27436 10968
rect 27488 10956 27494 11008
rect 2024 10906 77924 10928
rect 2024 10854 5794 10906
rect 5846 10854 5858 10906
rect 5910 10854 5922 10906
rect 5974 10854 5986 10906
rect 6038 10854 6050 10906
rect 6102 10854 36514 10906
rect 36566 10854 36578 10906
rect 36630 10854 36642 10906
rect 36694 10854 36706 10906
rect 36758 10854 36770 10906
rect 36822 10854 67234 10906
rect 67286 10854 67298 10906
rect 67350 10854 67362 10906
rect 67414 10854 67426 10906
rect 67478 10854 67490 10906
rect 67542 10854 77924 10906
rect 2024 10832 77924 10854
rect 13170 10752 13176 10804
rect 13228 10792 13234 10804
rect 24489 10795 24547 10801
rect 24489 10792 24501 10795
rect 13228 10764 24501 10792
rect 13228 10752 13234 10764
rect 24489 10761 24501 10764
rect 24535 10761 24547 10795
rect 24489 10755 24547 10761
rect 27709 10795 27767 10801
rect 27709 10761 27721 10795
rect 27755 10792 27767 10795
rect 28442 10792 28448 10804
rect 27755 10764 28448 10792
rect 27755 10761 27767 10764
rect 27709 10755 27767 10761
rect 13722 10684 13728 10736
rect 13780 10724 13786 10736
rect 13780 10696 21772 10724
rect 13780 10684 13786 10696
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 20533 10659 20591 10665
rect 20533 10656 20545 10659
rect 19392 10628 20545 10656
rect 19392 10616 19398 10628
rect 20533 10625 20545 10628
rect 20579 10625 20591 10659
rect 20533 10619 20591 10625
rect 20990 10616 20996 10668
rect 21048 10616 21054 10668
rect 21744 10665 21772 10696
rect 22554 10684 22560 10736
rect 22612 10724 22618 10736
rect 22612 10696 24256 10724
rect 22612 10684 22618 10696
rect 21545 10659 21603 10665
rect 21545 10656 21557 10659
rect 21100 10628 21557 10656
rect 15470 10548 15476 10600
rect 15528 10588 15534 10600
rect 21100 10588 21128 10628
rect 21545 10625 21557 10628
rect 21591 10625 21603 10659
rect 21545 10619 21603 10625
rect 21729 10659 21787 10665
rect 21729 10625 21741 10659
rect 21775 10656 21787 10659
rect 22741 10659 22799 10665
rect 22741 10656 22753 10659
rect 21775 10628 22753 10656
rect 21775 10625 21787 10628
rect 21729 10619 21787 10625
rect 22741 10625 22753 10628
rect 22787 10625 22799 10659
rect 22741 10619 22799 10625
rect 22922 10616 22928 10668
rect 22980 10616 22986 10668
rect 23014 10616 23020 10668
rect 23072 10656 23078 10668
rect 23661 10659 23719 10665
rect 23661 10656 23673 10659
rect 23072 10628 23673 10656
rect 23072 10616 23078 10628
rect 23661 10625 23673 10628
rect 23707 10625 23719 10659
rect 23661 10619 23719 10625
rect 15528 10560 21128 10588
rect 21269 10591 21327 10597
rect 15528 10548 15534 10560
rect 21269 10557 21281 10591
rect 21315 10588 21327 10591
rect 21315 10560 21772 10588
rect 21315 10557 21327 10560
rect 21269 10551 21327 10557
rect 17862 10480 17868 10532
rect 17920 10520 17926 10532
rect 21634 10520 21640 10532
rect 17920 10492 21640 10520
rect 17920 10480 17926 10492
rect 21634 10480 21640 10492
rect 21692 10480 21698 10532
rect 21744 10520 21772 10560
rect 22186 10548 22192 10600
rect 22244 10588 22250 10600
rect 22373 10591 22431 10597
rect 22373 10588 22385 10591
rect 22244 10560 22385 10588
rect 22244 10548 22250 10560
rect 22373 10557 22385 10560
rect 22419 10557 22431 10591
rect 23290 10588 23296 10600
rect 22373 10551 22431 10557
rect 22756 10560 23296 10588
rect 22756 10520 22784 10560
rect 23290 10548 23296 10560
rect 23348 10548 23354 10600
rect 23566 10548 23572 10600
rect 23624 10588 23630 10600
rect 24118 10588 24124 10600
rect 23624 10560 24124 10588
rect 23624 10548 23630 10560
rect 24118 10548 24124 10560
rect 24176 10548 24182 10600
rect 24228 10588 24256 10696
rect 24394 10616 24400 10668
rect 24452 10616 24458 10668
rect 24504 10656 24532 10755
rect 28442 10752 28448 10764
rect 28500 10752 28506 10804
rect 33318 10752 33324 10804
rect 33376 10752 33382 10804
rect 26786 10684 26792 10736
rect 26844 10724 26850 10736
rect 26844 10696 31754 10724
rect 26844 10684 26850 10696
rect 25225 10659 25283 10665
rect 25225 10656 25237 10659
rect 24504 10628 25237 10656
rect 25225 10625 25237 10628
rect 25271 10625 25283 10659
rect 25225 10619 25283 10625
rect 26050 10616 26056 10668
rect 26108 10656 26114 10668
rect 26237 10659 26295 10665
rect 26237 10656 26249 10659
rect 26108 10628 26249 10656
rect 26108 10616 26114 10628
rect 26237 10625 26249 10628
rect 26283 10625 26295 10659
rect 26510 10656 26516 10668
rect 26237 10619 26295 10625
rect 26344 10628 26516 10656
rect 26344 10588 26372 10628
rect 26510 10616 26516 10628
rect 26568 10656 26574 10668
rect 26605 10659 26663 10665
rect 26605 10656 26617 10659
rect 26568 10628 26617 10656
rect 26568 10616 26574 10628
rect 26605 10625 26617 10628
rect 26651 10625 26663 10659
rect 26605 10619 26663 10625
rect 28074 10616 28080 10668
rect 28132 10616 28138 10668
rect 31726 10656 31754 10696
rect 32033 10659 32091 10665
rect 32033 10656 32045 10659
rect 28184 10628 31064 10656
rect 31726 10628 32045 10656
rect 24228 10560 26372 10588
rect 26418 10548 26424 10600
rect 26476 10548 26482 10600
rect 27062 10548 27068 10600
rect 27120 10548 27126 10600
rect 21744 10492 22784 10520
rect 18966 10412 18972 10464
rect 19024 10452 19030 10464
rect 20625 10455 20683 10461
rect 20625 10452 20637 10455
rect 19024 10424 20637 10452
rect 19024 10412 19030 10424
rect 20625 10421 20637 10424
rect 20671 10421 20683 10455
rect 20625 10415 20683 10421
rect 20809 10455 20867 10461
rect 20809 10421 20821 10455
rect 20855 10452 20867 10455
rect 20898 10452 20904 10464
rect 20855 10424 20904 10452
rect 20855 10421 20867 10424
rect 20809 10415 20867 10421
rect 20898 10412 20904 10424
rect 20956 10412 20962 10464
rect 21174 10412 21180 10464
rect 21232 10412 21238 10464
rect 21450 10412 21456 10464
rect 21508 10452 21514 10464
rect 21744 10452 21772 10492
rect 22830 10480 22836 10532
rect 22888 10520 22894 10532
rect 23845 10523 23903 10529
rect 23845 10520 23857 10523
rect 22888 10492 23857 10520
rect 22888 10480 22894 10492
rect 23845 10489 23857 10492
rect 23891 10489 23903 10523
rect 24762 10520 24768 10532
rect 23845 10483 23903 10489
rect 24044 10492 24768 10520
rect 21508 10424 21772 10452
rect 21508 10412 21514 10424
rect 21818 10412 21824 10464
rect 21876 10412 21882 10464
rect 23106 10412 23112 10464
rect 23164 10412 23170 10464
rect 24044 10461 24072 10492
rect 24762 10480 24768 10492
rect 24820 10480 24826 10532
rect 26510 10480 26516 10532
rect 26568 10520 26574 10532
rect 28184 10520 28212 10628
rect 28810 10548 28816 10600
rect 28868 10548 28874 10600
rect 29733 10591 29791 10597
rect 29733 10588 29745 10591
rect 29012 10560 29745 10588
rect 26568 10492 28212 10520
rect 26568 10480 26574 10492
rect 29012 10464 29040 10560
rect 29733 10557 29745 10560
rect 29779 10557 29791 10591
rect 29733 10551 29791 10557
rect 30466 10548 30472 10600
rect 30524 10588 30530 10600
rect 30929 10591 30987 10597
rect 30929 10588 30941 10591
rect 30524 10560 30941 10588
rect 30524 10548 30530 10560
rect 30929 10557 30941 10560
rect 30975 10557 30987 10591
rect 31036 10588 31064 10628
rect 32033 10625 32045 10628
rect 32079 10625 32091 10659
rect 33336 10656 33364 10752
rect 34057 10659 34115 10665
rect 34057 10656 34069 10659
rect 33336 10628 34069 10656
rect 32033 10619 32091 10625
rect 34057 10625 34069 10628
rect 34103 10625 34115 10659
rect 34057 10619 34115 10625
rect 31036 10560 31754 10588
rect 30929 10551 30987 10557
rect 30837 10523 30895 10529
rect 30837 10489 30849 10523
rect 30883 10520 30895 10523
rect 31386 10520 31392 10532
rect 30883 10492 31392 10520
rect 30883 10489 30895 10492
rect 30837 10483 30895 10489
rect 31386 10480 31392 10492
rect 31444 10480 31450 10532
rect 31726 10520 31754 10560
rect 32766 10548 32772 10600
rect 32824 10548 32830 10600
rect 33137 10591 33195 10597
rect 33137 10557 33149 10591
rect 33183 10588 33195 10591
rect 33318 10588 33324 10600
rect 33183 10560 33324 10588
rect 33183 10557 33195 10560
rect 33137 10551 33195 10557
rect 33318 10548 33324 10560
rect 33376 10548 33382 10600
rect 34790 10548 34796 10600
rect 34848 10548 34854 10600
rect 35526 10548 35532 10600
rect 35584 10548 35590 10600
rect 33505 10523 33563 10529
rect 33505 10520 33517 10523
rect 31726 10492 33517 10520
rect 33505 10489 33517 10492
rect 33551 10489 33563 10523
rect 33505 10483 33563 10489
rect 34974 10480 34980 10532
rect 35032 10480 35038 10532
rect 24029 10455 24087 10461
rect 24029 10421 24041 10455
rect 24075 10421 24087 10455
rect 24029 10415 24087 10421
rect 24118 10412 24124 10464
rect 24176 10452 24182 10464
rect 24673 10455 24731 10461
rect 24673 10452 24685 10455
rect 24176 10424 24685 10452
rect 24176 10412 24182 10424
rect 24673 10421 24685 10424
rect 24719 10421 24731 10455
rect 24673 10415 24731 10421
rect 25222 10412 25228 10464
rect 25280 10452 25286 10464
rect 25501 10455 25559 10461
rect 25501 10452 25513 10455
rect 25280 10424 25513 10452
rect 25280 10412 25286 10424
rect 25501 10421 25513 10424
rect 25547 10421 25559 10455
rect 25501 10415 25559 10421
rect 26789 10455 26847 10461
rect 26789 10421 26801 10455
rect 26835 10452 26847 10455
rect 27522 10452 27528 10464
rect 26835 10424 27528 10452
rect 26835 10421 26847 10424
rect 26789 10415 26847 10421
rect 27522 10412 27528 10424
rect 27580 10412 27586 10464
rect 27614 10412 27620 10464
rect 27672 10452 27678 10464
rect 27893 10455 27951 10461
rect 27893 10452 27905 10455
rect 27672 10424 27905 10452
rect 27672 10412 27678 10424
rect 27893 10421 27905 10424
rect 27939 10421 27951 10455
rect 27893 10415 27951 10421
rect 28258 10412 28264 10464
rect 28316 10412 28322 10464
rect 28994 10412 29000 10464
rect 29052 10412 29058 10464
rect 29181 10455 29239 10461
rect 29181 10421 29193 10455
rect 29227 10452 29239 10455
rect 29270 10452 29276 10464
rect 29227 10424 29276 10452
rect 29227 10421 29239 10424
rect 29181 10415 29239 10421
rect 29270 10412 29276 10424
rect 29328 10412 29334 10464
rect 29546 10412 29552 10464
rect 29604 10452 29610 10464
rect 29917 10455 29975 10461
rect 29917 10452 29929 10455
rect 29604 10424 29929 10452
rect 29604 10412 29610 10424
rect 29917 10421 29929 10424
rect 29963 10421 29975 10455
rect 29917 10415 29975 10421
rect 31478 10412 31484 10464
rect 31536 10412 31542 10464
rect 31570 10412 31576 10464
rect 31628 10452 31634 10464
rect 32217 10455 32275 10461
rect 32217 10452 32229 10455
rect 31628 10424 32229 10452
rect 31628 10412 31634 10424
rect 32217 10421 32229 10424
rect 32263 10421 32275 10455
rect 32217 10415 32275 10421
rect 33134 10412 33140 10464
rect 33192 10452 33198 10464
rect 34241 10455 34299 10461
rect 34241 10452 34253 10455
rect 33192 10424 34253 10452
rect 33192 10412 33198 10424
rect 34241 10421 34253 10424
rect 34287 10421 34299 10455
rect 34241 10415 34299 10421
rect 2024 10362 77924 10384
rect 2024 10310 5134 10362
rect 5186 10310 5198 10362
rect 5250 10310 5262 10362
rect 5314 10310 5326 10362
rect 5378 10310 5390 10362
rect 5442 10310 35854 10362
rect 35906 10310 35918 10362
rect 35970 10310 35982 10362
rect 36034 10310 36046 10362
rect 36098 10310 36110 10362
rect 36162 10310 66574 10362
rect 66626 10310 66638 10362
rect 66690 10310 66702 10362
rect 66754 10310 66766 10362
rect 66818 10310 66830 10362
rect 66882 10310 77924 10362
rect 2024 10288 77924 10310
rect 14918 10208 14924 10260
rect 14976 10248 14982 10260
rect 23106 10248 23112 10260
rect 14976 10220 23112 10248
rect 14976 10208 14982 10220
rect 23106 10208 23112 10220
rect 23164 10208 23170 10260
rect 24026 10208 24032 10260
rect 24084 10248 24090 10260
rect 26329 10251 26387 10257
rect 26329 10248 26341 10251
rect 24084 10220 26341 10248
rect 24084 10208 24090 10220
rect 26329 10217 26341 10220
rect 26375 10217 26387 10251
rect 26329 10211 26387 10217
rect 27062 10208 27068 10260
rect 27120 10248 27126 10260
rect 27157 10251 27215 10257
rect 27157 10248 27169 10251
rect 27120 10220 27169 10248
rect 27120 10208 27126 10220
rect 27157 10217 27169 10220
rect 27203 10248 27215 10251
rect 30374 10248 30380 10260
rect 27203 10220 30380 10248
rect 27203 10217 27215 10220
rect 27157 10211 27215 10217
rect 30374 10208 30380 10220
rect 30432 10208 30438 10260
rect 17402 10140 17408 10192
rect 17460 10180 17466 10192
rect 20257 10183 20315 10189
rect 20257 10180 20269 10183
rect 17460 10152 20269 10180
rect 17460 10140 17466 10152
rect 20257 10149 20269 10152
rect 20303 10149 20315 10183
rect 20257 10143 20315 10149
rect 20622 10140 20628 10192
rect 20680 10180 20686 10192
rect 31478 10180 31484 10192
rect 20680 10152 31484 10180
rect 20680 10140 20686 10152
rect 31478 10140 31484 10152
rect 31536 10140 31542 10192
rect 32950 10180 32956 10192
rect 31726 10152 32956 10180
rect 19150 10072 19156 10124
rect 19208 10112 19214 10124
rect 21361 10115 21419 10121
rect 21361 10112 21373 10115
rect 19208 10084 21373 10112
rect 19208 10072 19214 10084
rect 21361 10081 21373 10084
rect 21407 10081 21419 10115
rect 22373 10115 22431 10121
rect 22373 10112 22385 10115
rect 21361 10075 21419 10081
rect 21468 10084 22385 10112
rect 19610 10004 19616 10056
rect 19668 10004 19674 10056
rect 19702 10004 19708 10056
rect 19760 10044 19766 10056
rect 19889 10047 19947 10053
rect 19889 10044 19901 10047
rect 19760 10016 19901 10044
rect 19760 10004 19766 10016
rect 19889 10013 19901 10016
rect 19935 10013 19947 10047
rect 19889 10007 19947 10013
rect 20438 10004 20444 10056
rect 20496 10044 20502 10056
rect 20533 10047 20591 10053
rect 20533 10044 20545 10047
rect 20496 10016 20545 10044
rect 20496 10004 20502 10016
rect 20533 10013 20545 10016
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 19794 9936 19800 9988
rect 19852 9976 19858 9988
rect 21468 9976 21496 10084
rect 22373 10081 22385 10084
rect 22419 10081 22431 10115
rect 22373 10075 22431 10081
rect 22738 10072 22744 10124
rect 22796 10112 22802 10124
rect 22925 10115 22983 10121
rect 22925 10112 22937 10115
rect 22796 10084 22937 10112
rect 22796 10072 22802 10084
rect 22925 10081 22937 10084
rect 22971 10081 22983 10115
rect 22925 10075 22983 10081
rect 23198 10072 23204 10124
rect 23256 10112 23262 10124
rect 23661 10115 23719 10121
rect 23661 10112 23673 10115
rect 23256 10084 23673 10112
rect 23256 10072 23262 10084
rect 23661 10081 23673 10084
rect 23707 10081 23719 10115
rect 23661 10075 23719 10081
rect 26237 10115 26295 10121
rect 26237 10081 26249 10115
rect 26283 10112 26295 10115
rect 26326 10112 26332 10124
rect 26283 10084 26332 10112
rect 26283 10081 26295 10084
rect 26237 10075 26295 10081
rect 26326 10072 26332 10084
rect 26384 10072 26390 10124
rect 27706 10072 27712 10124
rect 27764 10112 27770 10124
rect 28905 10115 28963 10121
rect 28905 10112 28917 10115
rect 27764 10084 28917 10112
rect 27764 10072 27770 10084
rect 28905 10081 28917 10084
rect 28951 10081 28963 10115
rect 28905 10075 28963 10081
rect 29546 10072 29552 10124
rect 29604 10072 29610 10124
rect 21634 10004 21640 10056
rect 21692 10044 21698 10056
rect 22097 10047 22155 10053
rect 22097 10044 22109 10047
rect 21692 10016 22109 10044
rect 21692 10004 21698 10016
rect 22097 10013 22109 10016
rect 22143 10013 22155 10047
rect 22097 10007 22155 10013
rect 23290 10004 23296 10056
rect 23348 10004 23354 10056
rect 24486 10004 24492 10056
rect 24544 10004 24550 10056
rect 26973 10047 27031 10053
rect 26973 10013 26985 10047
rect 27019 10040 27031 10047
rect 27430 10044 27436 10056
rect 27080 10040 27436 10044
rect 27019 10016 27436 10040
rect 27019 10013 27108 10016
rect 26973 10012 27108 10013
rect 26973 10007 27031 10012
rect 27430 10004 27436 10016
rect 27488 10004 27494 10056
rect 27982 10004 27988 10056
rect 28040 10004 28046 10056
rect 28169 10047 28227 10053
rect 28169 10013 28181 10047
rect 28215 10013 28227 10047
rect 28169 10007 28227 10013
rect 29733 10047 29791 10053
rect 29733 10013 29745 10047
rect 29779 10044 29791 10047
rect 29822 10044 29828 10056
rect 29779 10016 29828 10044
rect 29779 10013 29791 10016
rect 29733 10007 29791 10013
rect 19852 9948 21496 9976
rect 23385 9979 23443 9985
rect 19852 9936 19858 9948
rect 23385 9945 23397 9979
rect 23431 9976 23443 9979
rect 23569 9979 23627 9985
rect 23431 9948 23520 9976
rect 23431 9945 23443 9948
rect 23385 9939 23443 9945
rect 23492 9920 23520 9948
rect 23569 9945 23581 9979
rect 23615 9976 23627 9979
rect 23750 9976 23756 9988
rect 23615 9948 23756 9976
rect 23615 9945 23627 9948
rect 23569 9939 23627 9945
rect 23750 9936 23756 9948
rect 23808 9976 23814 9988
rect 23808 9948 27568 9976
rect 23808 9936 23814 9948
rect 27540 9920 27568 9948
rect 27614 9936 27620 9988
rect 27672 9976 27678 9988
rect 28184 9976 28212 10007
rect 29822 10004 29828 10016
rect 29880 10004 29886 10056
rect 31110 10004 31116 10056
rect 31168 10044 31174 10056
rect 31297 10047 31355 10053
rect 31297 10044 31309 10047
rect 31168 10016 31309 10044
rect 31168 10004 31174 10016
rect 31297 10013 31309 10016
rect 31343 10013 31355 10047
rect 31297 10007 31355 10013
rect 31726 9976 31754 10152
rect 32950 10140 32956 10152
rect 33008 10140 33014 10192
rect 33594 10140 33600 10192
rect 33652 10140 33658 10192
rect 31938 10004 31944 10056
rect 31996 10044 32002 10056
rect 32585 10047 32643 10053
rect 32585 10044 32597 10047
rect 31996 10016 32597 10044
rect 31996 10004 32002 10016
rect 32585 10013 32597 10016
rect 32631 10013 32643 10047
rect 32585 10007 32643 10013
rect 33410 10004 33416 10056
rect 33468 10004 33474 10056
rect 34238 10004 34244 10056
rect 34296 10004 34302 10056
rect 34882 10004 34888 10056
rect 34940 10004 34946 10056
rect 36354 10004 36360 10056
rect 36412 10044 36418 10056
rect 36449 10047 36507 10053
rect 36449 10044 36461 10047
rect 36412 10016 36461 10044
rect 36412 10004 36418 10016
rect 36449 10013 36461 10016
rect 36495 10013 36507 10047
rect 36449 10007 36507 10013
rect 36630 10004 36636 10056
rect 36688 10004 36694 10056
rect 37277 10047 37335 10053
rect 37277 10013 37289 10047
rect 37323 10044 37335 10047
rect 37642 10044 37648 10056
rect 37323 10016 37648 10044
rect 37323 10013 37335 10016
rect 37277 10007 37335 10013
rect 37642 10004 37648 10016
rect 37700 10004 37706 10056
rect 27672 9948 28212 9976
rect 28276 9948 31754 9976
rect 27672 9936 27678 9948
rect 19426 9868 19432 9920
rect 19484 9868 19490 9920
rect 19518 9868 19524 9920
rect 19576 9908 19582 9920
rect 19705 9911 19763 9917
rect 19705 9908 19717 9911
rect 19576 9880 19717 9908
rect 19576 9868 19582 9880
rect 19705 9877 19717 9880
rect 19751 9877 19763 9911
rect 19705 9871 19763 9877
rect 20806 9868 20812 9920
rect 20864 9868 20870 9920
rect 21542 9868 21548 9920
rect 21600 9868 21606 9920
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 23014 9908 23020 9920
rect 22152 9880 23020 9908
rect 22152 9868 22158 9880
rect 23014 9868 23020 9880
rect 23072 9908 23078 9920
rect 23109 9911 23167 9917
rect 23109 9908 23121 9911
rect 23072 9880 23121 9908
rect 23072 9868 23078 9880
rect 23109 9877 23121 9880
rect 23155 9877 23167 9911
rect 23109 9871 23167 9877
rect 23290 9868 23296 9920
rect 23348 9868 23354 9920
rect 23474 9868 23480 9920
rect 23532 9868 23538 9920
rect 24305 9911 24363 9917
rect 24305 9877 24317 9911
rect 24351 9908 24363 9911
rect 24578 9908 24584 9920
rect 24351 9880 24584 9908
rect 24351 9877 24363 9880
rect 24305 9871 24363 9877
rect 24578 9868 24584 9880
rect 24636 9868 24642 9920
rect 24670 9868 24676 9920
rect 24728 9908 24734 9920
rect 25041 9911 25099 9917
rect 25041 9908 25053 9911
rect 24728 9880 25053 9908
rect 24728 9868 24734 9880
rect 25041 9877 25053 9880
rect 25087 9877 25099 9911
rect 25041 9871 25099 9877
rect 25130 9868 25136 9920
rect 25188 9908 25194 9920
rect 25593 9911 25651 9917
rect 25593 9908 25605 9911
rect 25188 9880 25605 9908
rect 25188 9868 25194 9880
rect 25593 9877 25605 9880
rect 25639 9877 25651 9911
rect 25593 9871 25651 9877
rect 27246 9868 27252 9920
rect 27304 9908 27310 9920
rect 27433 9911 27491 9917
rect 27433 9908 27445 9911
rect 27304 9880 27445 9908
rect 27304 9868 27310 9880
rect 27433 9877 27445 9880
rect 27479 9877 27491 9911
rect 27433 9871 27491 9877
rect 27522 9868 27528 9920
rect 27580 9908 27586 9920
rect 28276 9908 28304 9948
rect 27580 9880 28304 9908
rect 27580 9868 27586 9880
rect 28718 9868 28724 9920
rect 28776 9908 28782 9920
rect 28813 9911 28871 9917
rect 28813 9908 28825 9911
rect 28776 9880 28825 9908
rect 28776 9868 28782 9880
rect 28813 9877 28825 9880
rect 28859 9877 28871 9911
rect 28813 9871 28871 9877
rect 30006 9868 30012 9920
rect 30064 9908 30070 9920
rect 30285 9911 30343 9917
rect 30285 9908 30297 9911
rect 30064 9880 30297 9908
rect 30064 9868 30070 9880
rect 30285 9877 30297 9880
rect 30331 9877 30343 9911
rect 30285 9871 30343 9877
rect 30558 9868 30564 9920
rect 30616 9868 30622 9920
rect 31846 9868 31852 9920
rect 31904 9908 31910 9920
rect 32033 9911 32091 9917
rect 32033 9908 32045 9911
rect 31904 9880 32045 9908
rect 31904 9868 31910 9880
rect 32033 9877 32045 9880
rect 32079 9877 32091 9911
rect 32033 9871 32091 9877
rect 32858 9868 32864 9920
rect 32916 9868 32922 9920
rect 34330 9868 34336 9920
rect 34388 9868 34394 9920
rect 35894 9868 35900 9920
rect 35952 9868 35958 9920
rect 2024 9818 77924 9840
rect 2024 9766 5794 9818
rect 5846 9766 5858 9818
rect 5910 9766 5922 9818
rect 5974 9766 5986 9818
rect 6038 9766 6050 9818
rect 6102 9766 36514 9818
rect 36566 9766 36578 9818
rect 36630 9766 36642 9818
rect 36694 9766 36706 9818
rect 36758 9766 36770 9818
rect 36822 9766 67234 9818
rect 67286 9766 67298 9818
rect 67350 9766 67362 9818
rect 67414 9766 67426 9818
rect 67478 9766 67490 9818
rect 67542 9766 77924 9818
rect 2024 9744 77924 9766
rect 13262 9664 13268 9716
rect 13320 9704 13326 9716
rect 16574 9704 16580 9716
rect 13320 9676 16580 9704
rect 13320 9664 13326 9676
rect 16574 9664 16580 9676
rect 16632 9664 16638 9716
rect 21726 9664 21732 9716
rect 21784 9704 21790 9716
rect 26418 9704 26424 9716
rect 21784 9676 26424 9704
rect 21784 9664 21790 9676
rect 26418 9664 26424 9676
rect 26476 9664 26482 9716
rect 31938 9704 31944 9716
rect 26528 9676 31944 9704
rect 18782 9596 18788 9648
rect 18840 9636 18846 9648
rect 20901 9639 20959 9645
rect 20901 9636 20913 9639
rect 18840 9608 20913 9636
rect 18840 9596 18846 9608
rect 20901 9605 20913 9608
rect 20947 9605 20959 9639
rect 20901 9599 20959 9605
rect 21082 9596 21088 9648
rect 21140 9636 21146 9648
rect 21140 9608 24256 9636
rect 21140 9596 21146 9608
rect 19245 9571 19303 9577
rect 19245 9537 19257 9571
rect 19291 9568 19303 9571
rect 19426 9568 19432 9580
rect 19291 9540 19432 9568
rect 19291 9537 19303 9540
rect 19245 9531 19303 9537
rect 19426 9528 19432 9540
rect 19484 9528 19490 9580
rect 22189 9571 22247 9577
rect 22189 9568 22201 9571
rect 19536 9540 22201 9568
rect 18506 9460 18512 9512
rect 18564 9500 18570 9512
rect 19536 9500 19564 9540
rect 22189 9537 22201 9540
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 22554 9528 22560 9580
rect 22612 9568 22618 9580
rect 23382 9568 23388 9580
rect 22612 9540 23388 9568
rect 22612 9528 22618 9540
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 24228 9577 24256 9608
rect 25590 9596 25596 9648
rect 25648 9636 25654 9648
rect 26528 9636 26556 9676
rect 31938 9664 31944 9676
rect 31996 9664 32002 9716
rect 34793 9707 34851 9713
rect 34793 9673 34805 9707
rect 34839 9704 34851 9707
rect 34882 9704 34888 9716
rect 34839 9676 34888 9704
rect 34839 9673 34851 9676
rect 34793 9667 34851 9673
rect 34882 9664 34888 9676
rect 34940 9664 34946 9716
rect 25648 9608 26556 9636
rect 27341 9639 27399 9645
rect 25648 9596 25654 9608
rect 27341 9605 27353 9639
rect 27387 9636 27399 9639
rect 28074 9636 28080 9648
rect 27387 9608 28080 9636
rect 27387 9605 27399 9608
rect 27341 9599 27399 9605
rect 28074 9596 28080 9608
rect 28132 9596 28138 9648
rect 31662 9636 31668 9648
rect 28184 9608 31668 9636
rect 24213 9571 24271 9577
rect 24213 9537 24225 9571
rect 24259 9537 24271 9571
rect 24213 9531 24271 9537
rect 25130 9528 25136 9580
rect 25188 9528 25194 9580
rect 25314 9528 25320 9580
rect 25372 9528 25378 9580
rect 26602 9528 26608 9580
rect 26660 9528 26666 9580
rect 26789 9571 26847 9577
rect 26789 9537 26801 9571
rect 26835 9568 26847 9571
rect 26878 9568 26884 9580
rect 26835 9540 26884 9568
rect 26835 9537 26847 9540
rect 26789 9531 26847 9537
rect 26878 9528 26884 9540
rect 26936 9528 26942 9580
rect 27433 9571 27491 9577
rect 27433 9537 27445 9571
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 18564 9472 19564 9500
rect 18564 9460 18570 9472
rect 19886 9460 19892 9512
rect 19944 9460 19950 9512
rect 20714 9460 20720 9512
rect 20772 9460 20778 9512
rect 21545 9503 21603 9509
rect 21545 9469 21557 9503
rect 21591 9500 21603 9503
rect 21726 9500 21732 9512
rect 21591 9472 21732 9500
rect 21591 9469 21603 9472
rect 21545 9463 21603 9469
rect 21726 9460 21732 9472
rect 21784 9460 21790 9512
rect 22465 9503 22523 9509
rect 22465 9469 22477 9503
rect 22511 9500 22523 9503
rect 22738 9500 22744 9512
rect 22511 9472 22744 9500
rect 22511 9469 22523 9472
rect 22465 9463 22523 9469
rect 22738 9460 22744 9472
rect 22796 9460 22802 9512
rect 23477 9503 23535 9509
rect 23477 9469 23489 9503
rect 23523 9469 23535 9503
rect 23477 9463 23535 9469
rect 19242 9392 19248 9444
rect 19300 9432 19306 9444
rect 20073 9435 20131 9441
rect 20073 9432 20085 9435
rect 19300 9404 20085 9432
rect 19300 9392 19306 9404
rect 20073 9401 20085 9404
rect 20119 9401 20131 9435
rect 20073 9395 20131 9401
rect 20254 9392 20260 9444
rect 20312 9432 20318 9444
rect 21637 9435 21695 9441
rect 21637 9432 21649 9435
rect 20312 9404 21649 9432
rect 20312 9392 20318 9404
rect 21637 9401 21649 9404
rect 21683 9401 21695 9435
rect 21637 9395 21695 9401
rect 22002 9392 22008 9444
rect 22060 9432 22066 9444
rect 23492 9432 23520 9463
rect 25958 9460 25964 9512
rect 26016 9460 26022 9512
rect 27448 9500 27476 9531
rect 27890 9528 27896 9580
rect 27948 9568 27954 9580
rect 27985 9571 28043 9577
rect 27985 9568 27997 9571
rect 27948 9540 27997 9568
rect 27948 9528 27954 9540
rect 27985 9537 27997 9540
rect 28031 9537 28043 9571
rect 27985 9531 28043 9537
rect 28184 9500 28212 9608
rect 31662 9596 31668 9608
rect 31720 9596 31726 9648
rect 35618 9596 35624 9648
rect 35676 9636 35682 9648
rect 35676 9608 37688 9636
rect 35676 9596 35682 9608
rect 28442 9528 28448 9580
rect 28500 9568 28506 9580
rect 28721 9571 28779 9577
rect 28721 9568 28733 9571
rect 28500 9540 28733 9568
rect 28500 9528 28506 9540
rect 28721 9537 28733 9540
rect 28767 9537 28779 9571
rect 28721 9531 28779 9537
rect 29549 9571 29607 9577
rect 29549 9537 29561 9571
rect 29595 9568 29607 9571
rect 30742 9568 30748 9580
rect 29595 9540 30748 9568
rect 29595 9537 29607 9540
rect 29549 9531 29607 9537
rect 30742 9528 30748 9540
rect 30800 9528 30806 9580
rect 32398 9568 32404 9580
rect 30852 9540 32404 9568
rect 27448 9472 28212 9500
rect 23750 9432 23756 9444
rect 22060 9404 23520 9432
rect 23584 9404 23756 9432
rect 22060 9392 22066 9404
rect 18598 9324 18604 9376
rect 18656 9324 18662 9376
rect 18690 9324 18696 9376
rect 18748 9364 18754 9376
rect 19337 9367 19395 9373
rect 19337 9364 19349 9367
rect 18748 9336 19349 9364
rect 18748 9324 18754 9336
rect 19337 9333 19349 9336
rect 19383 9333 19395 9367
rect 19337 9327 19395 9333
rect 20806 9324 20812 9376
rect 20864 9364 20870 9376
rect 22925 9367 22983 9373
rect 22925 9364 22937 9367
rect 20864 9336 22937 9364
rect 20864 9324 20870 9336
rect 22925 9333 22937 9336
rect 22971 9333 22983 9367
rect 22925 9327 22983 9333
rect 23474 9324 23480 9376
rect 23532 9364 23538 9376
rect 23584 9364 23612 9404
rect 23750 9392 23756 9404
rect 23808 9392 23814 9444
rect 24210 9392 24216 9444
rect 24268 9432 24274 9444
rect 24762 9432 24768 9444
rect 24268 9404 24768 9432
rect 24268 9392 24274 9404
rect 24762 9392 24768 9404
rect 24820 9432 24826 9444
rect 27448 9432 27476 9472
rect 28626 9460 28632 9512
rect 28684 9460 28690 9512
rect 30098 9460 30104 9512
rect 30156 9460 30162 9512
rect 30190 9460 30196 9512
rect 30248 9500 30254 9512
rect 30377 9503 30435 9509
rect 30377 9500 30389 9503
rect 30248 9472 30389 9500
rect 30248 9460 30254 9472
rect 30377 9469 30389 9472
rect 30423 9469 30435 9503
rect 30377 9463 30435 9469
rect 24820 9404 27476 9432
rect 27617 9435 27675 9441
rect 24820 9392 24826 9404
rect 27617 9401 27629 9435
rect 27663 9432 27675 9435
rect 27890 9432 27896 9444
rect 27663 9404 27896 9432
rect 27663 9401 27675 9404
rect 27617 9395 27675 9401
rect 27890 9392 27896 9404
rect 27948 9432 27954 9444
rect 30852 9432 30880 9540
rect 32398 9528 32404 9540
rect 32456 9528 32462 9580
rect 33505 9571 33563 9577
rect 33505 9537 33517 9571
rect 33551 9568 33563 9571
rect 34330 9568 34336 9580
rect 33551 9540 34336 9568
rect 33551 9537 33563 9540
rect 33505 9531 33563 9537
rect 34330 9528 34336 9540
rect 34388 9528 34394 9580
rect 34698 9528 34704 9580
rect 34756 9568 34762 9580
rect 35805 9571 35863 9577
rect 35805 9568 35817 9571
rect 34756 9540 35817 9568
rect 34756 9528 34762 9540
rect 35805 9537 35817 9540
rect 35851 9537 35863 9571
rect 35805 9531 35863 9537
rect 37366 9528 37372 9580
rect 37424 9568 37430 9580
rect 37660 9577 37688 9608
rect 37553 9571 37611 9577
rect 37553 9568 37565 9571
rect 37424 9540 37565 9568
rect 37424 9528 37430 9540
rect 37553 9537 37565 9540
rect 37599 9537 37611 9571
rect 37553 9531 37611 9537
rect 37645 9571 37703 9577
rect 37645 9537 37657 9571
rect 37691 9537 37703 9571
rect 37645 9531 37703 9537
rect 37826 9528 37832 9580
rect 37884 9528 37890 9580
rect 31202 9460 31208 9512
rect 31260 9460 31266 9512
rect 31570 9460 31576 9512
rect 31628 9500 31634 9512
rect 31849 9503 31907 9509
rect 31849 9500 31861 9503
rect 31628 9472 31861 9500
rect 31628 9460 31634 9472
rect 31849 9469 31861 9472
rect 31895 9469 31907 9503
rect 31849 9463 31907 9469
rect 34149 9503 34207 9509
rect 34149 9469 34161 9503
rect 34195 9469 34207 9503
rect 34149 9463 34207 9469
rect 34164 9432 34192 9463
rect 34882 9460 34888 9512
rect 34940 9500 34946 9512
rect 35069 9503 35127 9509
rect 35069 9500 35081 9503
rect 34940 9472 35081 9500
rect 34940 9460 34946 9472
rect 35069 9469 35081 9472
rect 35115 9469 35127 9503
rect 35069 9463 35127 9469
rect 35713 9503 35771 9509
rect 35713 9469 35725 9503
rect 35759 9500 35771 9503
rect 36357 9503 36415 9509
rect 36357 9500 36369 9503
rect 35759 9472 36369 9500
rect 35759 9469 35771 9472
rect 35713 9463 35771 9469
rect 36357 9469 36369 9472
rect 36403 9469 36415 9503
rect 36357 9463 36415 9469
rect 37277 9503 37335 9509
rect 37277 9469 37289 9503
rect 37323 9469 37335 9503
rect 37277 9463 37335 9469
rect 38841 9503 38899 9509
rect 38841 9469 38853 9503
rect 38887 9500 38899 9503
rect 40034 9500 40040 9512
rect 38887 9472 40040 9500
rect 38887 9469 38899 9472
rect 38841 9463 38899 9469
rect 27948 9404 30880 9432
rect 30944 9404 34192 9432
rect 27948 9392 27954 9404
rect 23532 9336 23612 9364
rect 23532 9324 23538 9336
rect 23658 9324 23664 9376
rect 23716 9324 23722 9376
rect 23842 9324 23848 9376
rect 23900 9364 23906 9376
rect 24489 9367 24547 9373
rect 24489 9364 24501 9367
rect 23900 9336 24501 9364
rect 23900 9324 23906 9336
rect 24489 9333 24501 9336
rect 24535 9333 24547 9367
rect 24489 9327 24547 9333
rect 25866 9324 25872 9376
rect 25924 9324 25930 9376
rect 27338 9324 27344 9376
rect 27396 9364 27402 9376
rect 27798 9364 27804 9376
rect 27396 9336 27804 9364
rect 27396 9324 27402 9336
rect 27798 9324 27804 9336
rect 27856 9324 27862 9376
rect 29365 9367 29423 9373
rect 29365 9333 29377 9367
rect 29411 9364 29423 9367
rect 29454 9364 29460 9376
rect 29411 9336 29460 9364
rect 29411 9333 29423 9336
rect 29365 9327 29423 9333
rect 29454 9324 29460 9336
rect 29512 9324 29518 9376
rect 30190 9324 30196 9376
rect 30248 9324 30254 9376
rect 30834 9324 30840 9376
rect 30892 9364 30898 9376
rect 30944 9364 30972 9404
rect 34330 9392 34336 9444
rect 34388 9432 34394 9444
rect 36541 9435 36599 9441
rect 36541 9432 36553 9435
rect 34388 9404 36553 9432
rect 34388 9392 34394 9404
rect 36541 9401 36553 9404
rect 36587 9432 36599 9435
rect 37292 9432 37320 9463
rect 40034 9460 40040 9472
rect 40092 9460 40098 9512
rect 36587 9404 37320 9432
rect 36587 9401 36599 9404
rect 36541 9395 36599 9401
rect 37734 9392 37740 9444
rect 37792 9392 37798 9444
rect 30892 9336 30972 9364
rect 31021 9367 31079 9373
rect 30892 9324 30898 9336
rect 31021 9333 31033 9367
rect 31067 9364 31079 9367
rect 31478 9364 31484 9376
rect 31067 9336 31484 9364
rect 31067 9333 31079 9336
rect 31021 9327 31079 9333
rect 31478 9324 31484 9336
rect 31536 9324 31542 9376
rect 31757 9367 31815 9373
rect 31757 9333 31769 9367
rect 31803 9364 31815 9367
rect 32306 9364 32312 9376
rect 31803 9336 32312 9364
rect 31803 9333 31815 9336
rect 31757 9327 31815 9333
rect 32306 9324 32312 9336
rect 32364 9324 32370 9376
rect 32493 9367 32551 9373
rect 32493 9333 32505 9367
rect 32539 9364 32551 9367
rect 32674 9364 32680 9376
rect 32539 9336 32680 9364
rect 32539 9333 32551 9336
rect 32493 9327 32551 9333
rect 32674 9324 32680 9336
rect 32732 9324 32738 9376
rect 34054 9324 34060 9376
rect 34112 9324 34118 9376
rect 34882 9324 34888 9376
rect 34940 9324 34946 9376
rect 36725 9367 36783 9373
rect 36725 9333 36737 9367
rect 36771 9364 36783 9367
rect 37182 9364 37188 9376
rect 36771 9336 37188 9364
rect 36771 9333 36783 9336
rect 36725 9327 36783 9333
rect 37182 9324 37188 9336
rect 37240 9324 37246 9376
rect 38010 9324 38016 9376
rect 38068 9324 38074 9376
rect 38194 9324 38200 9376
rect 38252 9324 38258 9376
rect 2024 9274 77924 9296
rect 2024 9222 5134 9274
rect 5186 9222 5198 9274
rect 5250 9222 5262 9274
rect 5314 9222 5326 9274
rect 5378 9222 5390 9274
rect 5442 9222 35854 9274
rect 35906 9222 35918 9274
rect 35970 9222 35982 9274
rect 36034 9222 36046 9274
rect 36098 9222 36110 9274
rect 36162 9222 66574 9274
rect 66626 9222 66638 9274
rect 66690 9222 66702 9274
rect 66754 9222 66766 9274
rect 66818 9222 66830 9274
rect 66882 9222 77924 9274
rect 2024 9200 77924 9222
rect 11698 9120 11704 9172
rect 11756 9120 11762 9172
rect 15562 9120 15568 9172
rect 15620 9160 15626 9172
rect 15620 9132 17356 9160
rect 15620 9120 15626 9132
rect 10594 9052 10600 9104
rect 10652 9092 10658 9104
rect 17129 9095 17187 9101
rect 17129 9092 17141 9095
rect 10652 9064 17141 9092
rect 10652 9052 10658 9064
rect 17129 9061 17141 9064
rect 17175 9061 17187 9095
rect 17328 9092 17356 9132
rect 19150 9120 19156 9172
rect 19208 9160 19214 9172
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 19208 9132 19257 9160
rect 19208 9120 19214 9132
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 19245 9123 19303 9129
rect 20990 9120 20996 9172
rect 21048 9160 21054 9172
rect 21269 9163 21327 9169
rect 21269 9160 21281 9163
rect 21048 9132 21281 9160
rect 21048 9120 21054 9132
rect 21269 9129 21281 9132
rect 21315 9129 21327 9163
rect 21269 9123 21327 9129
rect 22189 9163 22247 9169
rect 22189 9129 22201 9163
rect 22235 9160 22247 9163
rect 24670 9160 24676 9172
rect 22235 9132 24676 9160
rect 22235 9129 22247 9132
rect 22189 9123 22247 9129
rect 24670 9120 24676 9132
rect 24728 9120 24734 9172
rect 27430 9120 27436 9172
rect 27488 9160 27494 9172
rect 27488 9132 27844 9160
rect 27488 9120 27494 9132
rect 19334 9092 19340 9104
rect 17328 9064 19340 9092
rect 17129 9055 17187 9061
rect 19334 9052 19340 9064
rect 19392 9052 19398 9104
rect 20349 9095 20407 9101
rect 20349 9061 20361 9095
rect 20395 9092 20407 9095
rect 21634 9092 21640 9104
rect 20395 9064 21640 9092
rect 20395 9061 20407 9064
rect 20349 9055 20407 9061
rect 21634 9052 21640 9064
rect 21692 9092 21698 9104
rect 24394 9092 24400 9104
rect 21692 9064 24400 9092
rect 21692 9052 21698 9064
rect 24394 9052 24400 9064
rect 24452 9052 24458 9104
rect 25501 9095 25559 9101
rect 25501 9061 25513 9095
rect 25547 9092 25559 9095
rect 27816 9092 27844 9132
rect 28626 9120 28632 9172
rect 28684 9120 28690 9172
rect 28810 9120 28816 9172
rect 28868 9160 28874 9172
rect 29641 9163 29699 9169
rect 29641 9160 29653 9163
rect 28868 9132 29653 9160
rect 28868 9120 28874 9132
rect 29641 9129 29653 9132
rect 29687 9129 29699 9163
rect 29641 9123 29699 9129
rect 29914 9120 29920 9172
rect 29972 9160 29978 9172
rect 32217 9163 32275 9169
rect 32217 9160 32229 9163
rect 29972 9132 32229 9160
rect 29972 9120 29978 9132
rect 32217 9129 32229 9132
rect 32263 9129 32275 9163
rect 32217 9123 32275 9129
rect 32398 9120 32404 9172
rect 32456 9160 32462 9172
rect 32766 9160 32772 9172
rect 32456 9132 32772 9160
rect 32456 9120 32462 9132
rect 32766 9120 32772 9132
rect 32824 9160 32830 9172
rect 34514 9160 34520 9172
rect 32824 9132 34520 9160
rect 32824 9120 32830 9132
rect 34514 9120 34520 9132
rect 34572 9160 34578 9172
rect 35802 9160 35808 9172
rect 34572 9132 35808 9160
rect 34572 9120 34578 9132
rect 31570 9092 31576 9104
rect 25547 9064 27200 9092
rect 27816 9064 31576 9092
rect 25547 9061 25559 9064
rect 25501 9055 25559 9061
rect 15930 8984 15936 9036
rect 15988 9024 15994 9036
rect 17681 9027 17739 9033
rect 17681 9024 17693 9027
rect 15988 8996 17693 9024
rect 15988 8984 15994 8996
rect 17681 8993 17693 8996
rect 17727 8993 17739 9027
rect 17681 8987 17739 8993
rect 18322 8984 18328 9036
rect 18380 9024 18386 9036
rect 18509 9027 18567 9033
rect 18509 9024 18521 9027
rect 18380 8996 18521 9024
rect 18380 8984 18386 8996
rect 18509 8993 18521 8996
rect 18555 8993 18567 9027
rect 18509 8987 18567 8993
rect 19150 8984 19156 9036
rect 19208 9024 19214 9036
rect 21085 9027 21143 9033
rect 21085 9024 21097 9027
rect 19208 8996 21097 9024
rect 19208 8984 19214 8996
rect 21085 8993 21097 8996
rect 21131 8993 21143 9027
rect 21085 8987 21143 8993
rect 21266 8984 21272 9036
rect 21324 9024 21330 9036
rect 23569 9027 23627 9033
rect 23569 9024 23581 9027
rect 21324 8996 23581 9024
rect 21324 8984 21330 8996
rect 23569 8993 23581 8996
rect 23615 8993 23627 9027
rect 23569 8987 23627 8993
rect 25685 9027 25743 9033
rect 25685 8993 25697 9027
rect 25731 9024 25743 9027
rect 27065 9027 27123 9033
rect 27065 9024 27077 9027
rect 25731 8996 27077 9024
rect 25731 8993 25743 8996
rect 25685 8987 25743 8993
rect 27065 8993 27077 8996
rect 27111 8993 27123 9027
rect 27065 8987 27123 8993
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11296 8928 11621 8956
rect 11296 8916 11302 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 16485 8959 16543 8965
rect 16485 8956 16497 8959
rect 11609 8919 11667 8925
rect 12406 8928 16497 8956
rect 8846 8848 8852 8900
rect 8904 8888 8910 8900
rect 12406 8888 12434 8928
rect 16485 8925 16497 8928
rect 16531 8925 16543 8959
rect 16485 8919 16543 8925
rect 18414 8916 18420 8968
rect 18472 8956 18478 8968
rect 18601 8959 18659 8965
rect 18601 8956 18613 8959
rect 18472 8928 18613 8956
rect 18472 8916 18478 8928
rect 18601 8925 18613 8928
rect 18647 8925 18659 8959
rect 18601 8919 18659 8925
rect 18874 8916 18880 8968
rect 18932 8956 18938 8968
rect 19337 8959 19395 8965
rect 19337 8956 19349 8959
rect 18932 8928 19349 8956
rect 18932 8916 18938 8928
rect 19337 8925 19349 8928
rect 19383 8925 19395 8959
rect 19337 8919 19395 8925
rect 19610 8916 19616 8968
rect 19668 8956 19674 8968
rect 19794 8956 19800 8968
rect 19668 8928 19800 8956
rect 19668 8916 19674 8928
rect 19794 8916 19800 8928
rect 19852 8916 19858 8968
rect 20162 8916 20168 8968
rect 20220 8956 20226 8968
rect 20257 8959 20315 8965
rect 20257 8956 20269 8959
rect 20220 8928 20269 8956
rect 20220 8916 20226 8928
rect 20257 8925 20269 8928
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 20438 8916 20444 8968
rect 20496 8956 20502 8968
rect 21450 8956 21456 8968
rect 20496 8928 21456 8956
rect 20496 8916 20502 8928
rect 21450 8916 21456 8928
rect 21508 8916 21514 8968
rect 21818 8916 21824 8968
rect 21876 8916 21882 8968
rect 22005 8959 22063 8965
rect 22005 8925 22017 8959
rect 22051 8956 22063 8959
rect 22189 8959 22247 8965
rect 22051 8928 22140 8956
rect 22051 8925 22063 8928
rect 22005 8919 22063 8925
rect 8904 8860 12434 8888
rect 8904 8848 8910 8860
rect 16666 8848 16672 8900
rect 16724 8888 16730 8900
rect 20533 8891 20591 8897
rect 20533 8888 20545 8891
rect 16724 8860 20545 8888
rect 16724 8848 16730 8860
rect 20533 8857 20545 8860
rect 20579 8857 20591 8891
rect 20533 8851 20591 8857
rect 3234 8780 3240 8832
rect 3292 8820 3298 8832
rect 15933 8823 15991 8829
rect 15933 8820 15945 8823
rect 3292 8792 15945 8820
rect 3292 8780 3298 8792
rect 15933 8789 15945 8792
rect 15979 8789 15991 8823
rect 15933 8783 15991 8789
rect 17865 8823 17923 8829
rect 17865 8789 17877 8823
rect 17911 8820 17923 8823
rect 18230 8820 18236 8832
rect 17911 8792 18236 8820
rect 17911 8789 17923 8792
rect 17865 8783 17923 8789
rect 18230 8780 18236 8792
rect 18288 8780 18294 8832
rect 19794 8780 19800 8832
rect 19852 8820 19858 8832
rect 19981 8823 20039 8829
rect 19981 8820 19993 8823
rect 19852 8792 19993 8820
rect 19852 8780 19858 8792
rect 19981 8789 19993 8792
rect 20027 8789 20039 8823
rect 19981 8783 20039 8789
rect 21358 8780 21364 8832
rect 21416 8820 21422 8832
rect 22002 8820 22008 8832
rect 21416 8792 22008 8820
rect 21416 8780 21422 8792
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 22112 8820 22140 8928
rect 22189 8925 22201 8959
rect 22235 8925 22247 8959
rect 22189 8919 22247 8925
rect 22204 8888 22232 8919
rect 22554 8916 22560 8968
rect 22612 8916 22618 8968
rect 22646 8916 22652 8968
rect 22704 8916 22710 8968
rect 22741 8959 22799 8965
rect 22741 8925 22753 8959
rect 22787 8956 22799 8959
rect 22830 8956 22836 8968
rect 22787 8928 22836 8956
rect 22787 8925 22799 8928
rect 22741 8919 22799 8925
rect 22830 8916 22836 8928
rect 22888 8916 22894 8968
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8956 22983 8959
rect 23290 8956 23296 8968
rect 22971 8928 23296 8956
rect 22971 8925 22983 8928
rect 22925 8919 22983 8925
rect 23290 8916 23296 8928
rect 23348 8916 23354 8968
rect 23750 8916 23756 8968
rect 23808 8916 23814 8968
rect 24210 8956 24216 8968
rect 23860 8928 24216 8956
rect 22204 8860 22876 8888
rect 22848 8832 22876 8860
rect 23014 8848 23020 8900
rect 23072 8848 23078 8900
rect 23106 8848 23112 8900
rect 23164 8888 23170 8900
rect 23860 8888 23888 8928
rect 24210 8916 24216 8928
rect 24268 8956 24274 8968
rect 24673 8959 24731 8965
rect 24673 8956 24685 8959
rect 24268 8928 24685 8956
rect 24268 8916 24274 8928
rect 24673 8925 24685 8928
rect 24719 8925 24731 8959
rect 24673 8919 24731 8925
rect 24762 8916 24768 8968
rect 24820 8916 24826 8968
rect 25314 8916 25320 8968
rect 25372 8916 25378 8968
rect 26421 8959 26479 8965
rect 26421 8925 26433 8959
rect 26467 8925 26479 8959
rect 27172 8956 27200 9064
rect 31570 9052 31576 9064
rect 31628 9052 31634 9104
rect 31662 9052 31668 9104
rect 31720 9092 31726 9104
rect 34422 9092 34428 9104
rect 31720 9064 34428 9092
rect 31720 9052 31726 9064
rect 34422 9052 34428 9064
rect 34480 9052 34486 9104
rect 27798 8984 27804 9036
rect 27856 9024 27862 9036
rect 27985 9027 28043 9033
rect 27985 9024 27997 9027
rect 27856 8996 27997 9024
rect 27856 8984 27862 8996
rect 27985 8993 27997 8996
rect 28031 8993 28043 9027
rect 27985 8987 28043 8993
rect 29457 9027 29515 9033
rect 29457 8993 29469 9027
rect 29503 9024 29515 9027
rect 30282 9024 30288 9036
rect 29503 8996 30288 9024
rect 29503 8993 29515 8996
rect 29457 8987 29515 8993
rect 30282 8984 30288 8996
rect 30340 8984 30346 9036
rect 32769 9027 32827 9033
rect 32769 9024 32781 9027
rect 31312 8996 32781 9024
rect 27617 8959 27675 8965
rect 27617 8956 27629 8959
rect 27172 8928 27629 8956
rect 26421 8919 26479 8925
rect 27617 8925 27629 8928
rect 27663 8925 27675 8959
rect 27617 8919 27675 8925
rect 23164 8860 23888 8888
rect 23164 8848 23170 8860
rect 23934 8848 23940 8900
rect 23992 8888 23998 8900
rect 24489 8891 24547 8897
rect 24489 8888 24501 8891
rect 23992 8860 24501 8888
rect 23992 8848 23998 8860
rect 24489 8857 24501 8860
rect 24535 8857 24547 8891
rect 26436 8888 26464 8919
rect 28074 8916 28080 8968
rect 28132 8956 28138 8968
rect 28905 8959 28963 8965
rect 28905 8956 28917 8959
rect 28132 8928 28917 8956
rect 28132 8916 28138 8928
rect 28905 8925 28917 8928
rect 28951 8925 28963 8959
rect 28905 8919 28963 8925
rect 29546 8916 29552 8968
rect 29604 8956 29610 8968
rect 30193 8959 30251 8965
rect 30193 8956 30205 8959
rect 29604 8928 30205 8956
rect 29604 8916 29610 8928
rect 30193 8925 30205 8928
rect 30239 8925 30251 8959
rect 30193 8919 30251 8925
rect 30558 8916 30564 8968
rect 30616 8956 30622 8968
rect 31312 8965 31340 8996
rect 32769 8993 32781 8996
rect 32815 9024 32827 9027
rect 33042 9024 33048 9036
rect 32815 8996 33048 9024
rect 32815 8993 32827 8996
rect 32769 8987 32827 8993
rect 33042 8984 33048 8996
rect 33100 8984 33106 9036
rect 34606 8984 34612 9036
rect 34664 8984 34670 9036
rect 31297 8959 31355 8965
rect 31297 8956 31309 8959
rect 30616 8928 31309 8956
rect 30616 8916 30622 8928
rect 31297 8925 31309 8928
rect 31343 8925 31355 8959
rect 31297 8919 31355 8925
rect 31389 8959 31447 8965
rect 31389 8925 31401 8959
rect 31435 8956 31447 8959
rect 31570 8956 31576 8968
rect 31435 8928 31576 8956
rect 31435 8925 31447 8928
rect 31389 8919 31447 8925
rect 31570 8916 31576 8928
rect 31628 8916 31634 8968
rect 33962 8916 33968 8968
rect 34020 8916 34026 8968
rect 34716 8956 34744 9132
rect 35802 9120 35808 9132
rect 35860 9160 35866 9172
rect 37734 9160 37740 9172
rect 35860 9132 37740 9160
rect 35860 9120 35866 9132
rect 37734 9120 37740 9132
rect 37792 9120 37798 9172
rect 34974 9092 34980 9104
rect 34900 9064 34980 9092
rect 34900 9024 34928 9064
rect 34974 9052 34980 9064
rect 35032 9052 35038 9104
rect 35437 9095 35495 9101
rect 35437 9061 35449 9095
rect 35483 9092 35495 9095
rect 36170 9092 36176 9104
rect 35483 9064 36176 9092
rect 35483 9061 35495 9064
rect 35437 9055 35495 9061
rect 36170 9052 36176 9064
rect 36228 9052 36234 9104
rect 36817 9027 36875 9033
rect 36817 9024 36829 9027
rect 34900 8996 34954 9024
rect 34926 8965 34954 8996
rect 34793 8959 34851 8965
rect 34793 8956 34805 8959
rect 34716 8928 34805 8956
rect 34793 8925 34805 8928
rect 34839 8925 34851 8959
rect 34793 8919 34851 8925
rect 34885 8959 34954 8965
rect 34885 8925 34897 8959
rect 34931 8930 34954 8959
rect 34992 8996 36829 9024
rect 34931 8925 34943 8930
rect 34885 8919 34943 8925
rect 28258 8888 28264 8900
rect 24489 8851 24547 8857
rect 25884 8860 26372 8888
rect 26436 8860 28264 8888
rect 25884 8832 25912 8860
rect 22186 8820 22192 8832
rect 22112 8792 22192 8820
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 22278 8780 22284 8832
rect 22336 8780 22342 8832
rect 22830 8780 22836 8832
rect 22888 8780 22894 8832
rect 24210 8780 24216 8832
rect 24268 8820 24274 8832
rect 24397 8823 24455 8829
rect 24397 8820 24409 8823
rect 24268 8792 24409 8820
rect 24268 8780 24274 8792
rect 24397 8789 24409 8792
rect 24443 8789 24455 8823
rect 24397 8783 24455 8789
rect 25130 8780 25136 8832
rect 25188 8780 25194 8832
rect 25866 8780 25872 8832
rect 25924 8780 25930 8832
rect 26234 8780 26240 8832
rect 26292 8780 26298 8832
rect 26344 8820 26372 8860
rect 28258 8848 28264 8860
rect 28316 8848 28322 8900
rect 30926 8848 30932 8900
rect 30984 8848 30990 8900
rect 31662 8848 31668 8900
rect 31720 8848 31726 8900
rect 31757 8891 31815 8897
rect 31757 8857 31769 8891
rect 31803 8888 31815 8891
rect 32398 8888 32404 8900
rect 31803 8860 32404 8888
rect 31803 8857 31815 8860
rect 31757 8851 31815 8857
rect 32398 8848 32404 8860
rect 32456 8848 32462 8900
rect 33042 8848 33048 8900
rect 33100 8888 33106 8900
rect 34992 8888 35020 8996
rect 36817 8993 36829 8996
rect 36863 8993 36875 9027
rect 36817 8987 36875 8993
rect 38746 8984 38752 9036
rect 38804 9024 38810 9036
rect 40037 9027 40095 9033
rect 40037 9024 40049 9027
rect 38804 8996 40049 9024
rect 38804 8984 38810 8996
rect 40037 8993 40049 8996
rect 40083 8993 40095 9027
rect 40037 8987 40095 8993
rect 35158 8916 35164 8968
rect 35216 8916 35222 8968
rect 35250 8916 35256 8968
rect 35308 8916 35314 8968
rect 35802 8916 35808 8968
rect 35860 8916 35866 8968
rect 35989 8959 36047 8965
rect 35989 8925 36001 8959
rect 36035 8925 36047 8959
rect 35989 8919 36047 8925
rect 33100 8860 35020 8888
rect 33100 8848 33106 8860
rect 35066 8848 35072 8900
rect 35124 8848 35130 8900
rect 36004 8888 36032 8919
rect 36354 8916 36360 8968
rect 36412 8956 36418 8968
rect 36633 8959 36691 8965
rect 36633 8956 36645 8959
rect 36412 8928 36645 8956
rect 36412 8916 36418 8928
rect 36633 8925 36645 8928
rect 36679 8925 36691 8959
rect 36633 8919 36691 8925
rect 36998 8916 37004 8968
rect 37056 8956 37062 8968
rect 37369 8959 37427 8965
rect 37369 8956 37381 8959
rect 37056 8928 37381 8956
rect 37056 8916 37062 8928
rect 37369 8925 37381 8928
rect 37415 8925 37427 8959
rect 37369 8919 37427 8925
rect 38194 8916 38200 8968
rect 38252 8916 38258 8968
rect 38841 8959 38899 8965
rect 38841 8925 38853 8959
rect 38887 8956 38899 8959
rect 39485 8959 39543 8965
rect 39485 8956 39497 8959
rect 38887 8928 39497 8956
rect 38887 8925 38899 8928
rect 38841 8919 38899 8925
rect 39485 8925 39497 8928
rect 39531 8925 39543 8959
rect 39485 8919 39543 8925
rect 38654 8888 38660 8900
rect 36004 8860 38660 8888
rect 38654 8848 38660 8860
rect 38712 8848 38718 8900
rect 26602 8820 26608 8832
rect 26344 8792 26608 8820
rect 26602 8780 26608 8792
rect 26660 8780 26666 8832
rect 26973 8823 27031 8829
rect 26973 8789 26985 8823
rect 27019 8820 27031 8823
rect 28166 8820 28172 8832
rect 27019 8792 28172 8820
rect 27019 8789 27031 8792
rect 26973 8783 27031 8789
rect 28166 8780 28172 8792
rect 28224 8780 28230 8832
rect 31110 8780 31116 8832
rect 31168 8780 31174 8832
rect 33226 8780 33232 8832
rect 33284 8820 33290 8832
rect 33321 8823 33379 8829
rect 33321 8820 33333 8823
rect 33284 8792 33333 8820
rect 33284 8780 33290 8792
rect 33321 8789 33333 8792
rect 33367 8789 33379 8823
rect 33321 8783 33379 8789
rect 33502 8780 33508 8832
rect 33560 8820 33566 8832
rect 34057 8823 34115 8829
rect 34057 8820 34069 8823
rect 33560 8792 34069 8820
rect 33560 8780 33566 8792
rect 34057 8789 34069 8792
rect 34103 8789 34115 8823
rect 34057 8783 34115 8789
rect 34146 8780 34152 8832
rect 34204 8820 34210 8832
rect 35621 8823 35679 8829
rect 35621 8820 35633 8823
rect 34204 8792 35633 8820
rect 34204 8780 34210 8792
rect 35621 8789 35633 8792
rect 35667 8789 35679 8823
rect 35621 8783 35679 8789
rect 36081 8823 36139 8829
rect 36081 8789 36093 8823
rect 36127 8820 36139 8823
rect 36906 8820 36912 8832
rect 36127 8792 36912 8820
rect 36127 8789 36139 8792
rect 36081 8783 36139 8789
rect 36906 8780 36912 8792
rect 36964 8780 36970 8832
rect 37458 8780 37464 8832
rect 37516 8820 37522 8832
rect 37553 8823 37611 8829
rect 37553 8820 37565 8823
rect 37516 8792 37565 8820
rect 37516 8780 37522 8792
rect 37553 8789 37565 8792
rect 37599 8789 37611 8823
rect 37553 8783 37611 8789
rect 39393 8823 39451 8829
rect 39393 8789 39405 8823
rect 39439 8820 39451 8823
rect 39758 8820 39764 8832
rect 39439 8792 39764 8820
rect 39439 8789 39451 8792
rect 39393 8783 39451 8789
rect 39758 8780 39764 8792
rect 39816 8780 39822 8832
rect 2024 8730 77924 8752
rect 2024 8678 5794 8730
rect 5846 8678 5858 8730
rect 5910 8678 5922 8730
rect 5974 8678 5986 8730
rect 6038 8678 6050 8730
rect 6102 8678 36514 8730
rect 36566 8678 36578 8730
rect 36630 8678 36642 8730
rect 36694 8678 36706 8730
rect 36758 8678 36770 8730
rect 36822 8678 67234 8730
rect 67286 8678 67298 8730
rect 67350 8678 67362 8730
rect 67414 8678 67426 8730
rect 67478 8678 67490 8730
rect 67542 8678 77924 8730
rect 2024 8656 77924 8678
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 18690 8616 18696 8628
rect 11756 8588 18696 8616
rect 11756 8576 11762 8588
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 18874 8576 18880 8628
rect 18932 8576 18938 8628
rect 21358 8616 21364 8628
rect 18984 8588 21364 8616
rect 18138 8508 18144 8560
rect 18196 8508 18202 8560
rect 13998 8440 14004 8492
rect 14056 8480 14062 8492
rect 14056 8452 16988 8480
rect 14056 8440 14062 8452
rect 14642 8372 14648 8424
rect 14700 8412 14706 8424
rect 16025 8415 16083 8421
rect 16025 8412 16037 8415
rect 14700 8384 16037 8412
rect 14700 8372 14706 8384
rect 16025 8381 16037 8384
rect 16071 8381 16083 8415
rect 16025 8375 16083 8381
rect 16669 8415 16727 8421
rect 16669 8381 16681 8415
rect 16715 8412 16727 8415
rect 16850 8412 16856 8424
rect 16715 8384 16856 8412
rect 16715 8381 16727 8384
rect 16669 8375 16727 8381
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 3970 8304 3976 8356
rect 4028 8344 4034 8356
rect 16761 8347 16819 8353
rect 16761 8344 16773 8347
rect 4028 8316 16773 8344
rect 4028 8304 4034 8316
rect 16761 8313 16773 8316
rect 16807 8313 16819 8347
rect 16960 8344 16988 8452
rect 17770 8440 17776 8492
rect 17828 8440 17834 8492
rect 18046 8440 18052 8492
rect 18104 8480 18110 8492
rect 18984 8480 19012 8588
rect 21358 8576 21364 8588
rect 21416 8576 21422 8628
rect 21821 8619 21879 8625
rect 21821 8585 21833 8619
rect 21867 8616 21879 8619
rect 22554 8616 22560 8628
rect 21867 8588 22560 8616
rect 21867 8585 21879 8588
rect 21821 8579 21879 8585
rect 22554 8576 22560 8588
rect 22612 8576 22618 8628
rect 22830 8576 22836 8628
rect 22888 8616 22894 8628
rect 23382 8616 23388 8628
rect 22888 8588 23388 8616
rect 22888 8576 22894 8588
rect 23382 8576 23388 8588
rect 23440 8576 23446 8628
rect 24302 8576 24308 8628
rect 24360 8616 24366 8628
rect 29914 8616 29920 8628
rect 24360 8588 29920 8616
rect 24360 8576 24366 8588
rect 29914 8576 29920 8588
rect 29972 8576 29978 8628
rect 30098 8576 30104 8628
rect 30156 8616 30162 8628
rect 30650 8616 30656 8628
rect 30156 8588 30656 8616
rect 30156 8576 30162 8588
rect 21542 8548 21548 8560
rect 19628 8520 21548 8548
rect 19628 8489 19656 8520
rect 21542 8508 21548 8520
rect 21600 8508 21606 8560
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 22646 8548 22652 8560
rect 21784 8520 22652 8548
rect 21784 8508 21790 8520
rect 22646 8508 22652 8520
rect 22704 8508 22710 8560
rect 23842 8508 23848 8560
rect 23900 8508 23906 8560
rect 24210 8508 24216 8560
rect 24268 8508 24274 8560
rect 25866 8508 25872 8560
rect 25924 8548 25930 8560
rect 25961 8551 26019 8557
rect 25961 8548 25973 8551
rect 25924 8520 25973 8548
rect 25924 8508 25930 8520
rect 25961 8517 25973 8520
rect 26007 8517 26019 8551
rect 25961 8511 26019 8517
rect 26234 8508 26240 8560
rect 26292 8548 26298 8560
rect 26292 8520 27108 8548
rect 26292 8508 26298 8520
rect 18104 8452 19012 8480
rect 19613 8483 19671 8489
rect 18104 8440 18110 8452
rect 19613 8449 19625 8483
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 19978 8440 19984 8492
rect 20036 8480 20042 8492
rect 20993 8483 21051 8489
rect 20993 8480 21005 8483
rect 20036 8452 21005 8480
rect 20036 8440 20042 8452
rect 20993 8449 21005 8452
rect 21039 8449 21051 8483
rect 20993 8443 21051 8449
rect 22005 8483 22063 8489
rect 22005 8449 22017 8483
rect 22051 8480 22063 8483
rect 22278 8480 22284 8492
rect 22051 8452 22284 8480
rect 22051 8449 22063 8452
rect 22005 8443 22063 8449
rect 22278 8440 22284 8452
rect 22336 8440 22342 8492
rect 22554 8440 22560 8492
rect 22612 8440 22618 8492
rect 22830 8440 22836 8492
rect 22888 8440 22894 8492
rect 23753 8483 23811 8489
rect 23753 8449 23765 8483
rect 23799 8480 23811 8483
rect 23860 8480 23888 8508
rect 26418 8480 26424 8492
rect 23799 8452 23888 8480
rect 25346 8452 26424 8480
rect 23799 8449 23811 8452
rect 23753 8443 23811 8449
rect 26418 8440 26424 8452
rect 26476 8440 26482 8492
rect 27080 8489 27108 8520
rect 27522 8508 27528 8560
rect 27580 8548 27586 8560
rect 27985 8551 28043 8557
rect 27985 8548 27997 8551
rect 27580 8520 27997 8548
rect 27580 8508 27586 8520
rect 27985 8517 27997 8520
rect 28031 8517 28043 8551
rect 30190 8548 30196 8560
rect 27985 8511 28043 8517
rect 29564 8520 30196 8548
rect 26789 8483 26847 8489
rect 26789 8480 26801 8483
rect 26528 8452 26801 8480
rect 17034 8372 17040 8424
rect 17092 8412 17098 8424
rect 17313 8415 17371 8421
rect 17313 8412 17325 8415
rect 17092 8384 17325 8412
rect 17092 8372 17098 8384
rect 17313 8381 17325 8384
rect 17359 8381 17371 8415
rect 17313 8375 17371 8381
rect 18325 8415 18383 8421
rect 18325 8381 18337 8415
rect 18371 8381 18383 8415
rect 18325 8375 18383 8381
rect 16960 8316 18092 8344
rect 16761 8307 16819 8313
rect 15194 8236 15200 8288
rect 15252 8276 15258 8288
rect 17862 8276 17868 8288
rect 15252 8248 17868 8276
rect 15252 8236 15258 8248
rect 17862 8236 17868 8248
rect 17920 8236 17926 8288
rect 18064 8276 18092 8316
rect 18138 8304 18144 8356
rect 18196 8344 18202 8356
rect 18340 8344 18368 8375
rect 20254 8372 20260 8424
rect 20312 8372 20318 8424
rect 20346 8372 20352 8424
rect 20404 8412 20410 8424
rect 21177 8415 21235 8421
rect 21177 8412 21189 8415
rect 20404 8384 21189 8412
rect 20404 8372 20410 8384
rect 21177 8381 21189 8384
rect 21223 8381 21235 8415
rect 23201 8415 23259 8421
rect 23201 8412 23213 8415
rect 21177 8375 21235 8381
rect 22066 8384 23213 8412
rect 18196 8316 18368 8344
rect 18196 8304 18202 8316
rect 18874 8304 18880 8356
rect 18932 8344 18938 8356
rect 20441 8347 20499 8353
rect 20441 8344 20453 8347
rect 18932 8316 20453 8344
rect 18932 8304 18938 8316
rect 20441 8313 20453 8316
rect 20487 8313 20499 8347
rect 20441 8307 20499 8313
rect 22066 8288 22094 8384
rect 23201 8381 23213 8384
rect 23247 8381 23259 8415
rect 23201 8375 23259 8381
rect 23937 8415 23995 8421
rect 23937 8381 23949 8415
rect 23983 8381 23995 8415
rect 23937 8375 23995 8381
rect 22370 8304 22376 8356
rect 22428 8344 22434 8356
rect 23952 8344 23980 8375
rect 25958 8372 25964 8424
rect 26016 8412 26022 8424
rect 26528 8412 26556 8452
rect 26789 8449 26801 8452
rect 26835 8449 26847 8483
rect 26789 8443 26847 8449
rect 26973 8483 27031 8489
rect 26973 8449 26985 8483
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27065 8483 27123 8489
rect 27065 8449 27077 8483
rect 27111 8449 27123 8483
rect 27065 8443 27123 8449
rect 26016 8384 26556 8412
rect 26016 8372 26022 8384
rect 26602 8372 26608 8424
rect 26660 8372 26666 8424
rect 26988 8412 27016 8443
rect 27798 8440 27804 8492
rect 27856 8480 27862 8492
rect 27893 8483 27951 8489
rect 27893 8480 27905 8483
rect 27856 8452 27905 8480
rect 27856 8440 27862 8452
rect 27893 8449 27905 8452
rect 27939 8449 27951 8483
rect 27893 8443 27951 8449
rect 28077 8483 28135 8489
rect 28077 8449 28089 8483
rect 28123 8480 28135 8483
rect 28123 8452 28488 8480
rect 28123 8449 28135 8452
rect 28077 8443 28135 8449
rect 28460 8424 28488 8452
rect 28534 8440 28540 8492
rect 28592 8480 28598 8492
rect 28721 8483 28779 8489
rect 28721 8480 28733 8483
rect 28592 8452 28733 8480
rect 28592 8440 28598 8452
rect 28721 8449 28733 8452
rect 28767 8449 28779 8483
rect 28721 8443 28779 8449
rect 29454 8440 29460 8492
rect 29512 8440 29518 8492
rect 27154 8412 27160 8424
rect 26988 8384 27160 8412
rect 27154 8372 27160 8384
rect 27212 8372 27218 8424
rect 27706 8372 27712 8424
rect 27764 8372 27770 8424
rect 28442 8372 28448 8424
rect 28500 8372 28506 8424
rect 22428 8316 23980 8344
rect 22428 8304 22434 8316
rect 25774 8304 25780 8356
rect 25832 8344 25838 8356
rect 26789 8347 26847 8353
rect 26789 8344 26801 8347
rect 25832 8316 26801 8344
rect 25832 8304 25838 8316
rect 26789 8313 26801 8316
rect 26835 8313 26847 8347
rect 26789 8307 26847 8313
rect 26878 8304 26884 8356
rect 26936 8344 26942 8356
rect 28169 8347 28227 8353
rect 28169 8344 28181 8347
rect 26936 8316 28181 8344
rect 26936 8304 26942 8316
rect 28169 8313 28181 8316
rect 28215 8313 28227 8347
rect 28169 8307 28227 8313
rect 29454 8304 29460 8356
rect 29512 8344 29518 8356
rect 29564 8344 29592 8520
rect 30190 8508 30196 8520
rect 30248 8508 30254 8560
rect 30300 8548 30328 8588
rect 30650 8576 30656 8588
rect 30708 8576 30714 8628
rect 32214 8576 32220 8628
rect 32272 8616 32278 8628
rect 32651 8619 32709 8625
rect 32651 8616 32663 8619
rect 32272 8588 32663 8616
rect 32272 8576 32278 8588
rect 32651 8585 32663 8588
rect 32697 8585 32709 8619
rect 32651 8579 32709 8585
rect 35250 8576 35256 8628
rect 35308 8616 35314 8628
rect 35894 8616 35900 8628
rect 35308 8588 35900 8616
rect 35308 8576 35314 8588
rect 35894 8576 35900 8588
rect 35952 8576 35958 8628
rect 30300 8520 30406 8548
rect 31294 8508 31300 8560
rect 31352 8548 31358 8560
rect 31665 8551 31723 8557
rect 31665 8548 31677 8551
rect 31352 8520 31677 8548
rect 31352 8508 31358 8520
rect 31665 8517 31677 8520
rect 31711 8517 31723 8551
rect 31665 8511 31723 8517
rect 29641 8415 29699 8421
rect 29641 8381 29653 8415
rect 29687 8381 29699 8415
rect 29641 8375 29699 8381
rect 29512 8316 29592 8344
rect 29512 8304 29518 8316
rect 29656 8288 29684 8375
rect 29914 8372 29920 8424
rect 29972 8372 29978 8424
rect 31680 8412 31708 8511
rect 32030 8508 32036 8560
rect 32088 8548 32094 8560
rect 32861 8551 32919 8557
rect 32861 8548 32873 8551
rect 32088 8520 32873 8548
rect 32088 8508 32094 8520
rect 32861 8517 32873 8520
rect 32907 8517 32919 8551
rect 32861 8511 32919 8517
rect 33686 8508 33692 8560
rect 33744 8548 33750 8560
rect 35066 8548 35072 8560
rect 33744 8520 35072 8548
rect 33744 8508 33750 8520
rect 35066 8508 35072 8520
rect 35124 8548 35130 8560
rect 35434 8548 35440 8560
rect 35124 8520 35440 8548
rect 35124 8508 35130 8520
rect 35434 8508 35440 8520
rect 35492 8508 35498 8560
rect 37550 8508 37556 8560
rect 37608 8548 37614 8560
rect 38197 8551 38255 8557
rect 38197 8548 38209 8551
rect 37608 8520 38209 8548
rect 37608 8508 37614 8520
rect 38197 8517 38209 8520
rect 38243 8517 38255 8551
rect 38197 8511 38255 8517
rect 32214 8440 32220 8492
rect 32272 8480 32278 8492
rect 33597 8483 33655 8489
rect 33597 8480 33609 8483
rect 32272 8452 33609 8480
rect 32272 8440 32278 8452
rect 33597 8449 33609 8452
rect 33643 8449 33655 8483
rect 33597 8443 33655 8449
rect 33778 8440 33784 8492
rect 33836 8480 33842 8492
rect 34885 8483 34943 8489
rect 34885 8480 34897 8483
rect 33836 8452 34897 8480
rect 33836 8440 33842 8452
rect 34885 8449 34897 8452
rect 34931 8449 34943 8483
rect 34885 8443 34943 8449
rect 36262 8440 36268 8492
rect 36320 8480 36326 8492
rect 36722 8480 36728 8492
rect 36320 8452 36728 8480
rect 36320 8440 36326 8452
rect 36722 8440 36728 8452
rect 36780 8440 36786 8492
rect 39758 8440 39764 8492
rect 39816 8440 39822 8492
rect 32309 8415 32367 8421
rect 32309 8412 32321 8415
rect 31680 8384 32321 8412
rect 32309 8381 32321 8384
rect 32355 8381 32367 8415
rect 32309 8375 32367 8381
rect 32398 8372 32404 8424
rect 32456 8412 32462 8424
rect 33045 8415 33103 8421
rect 33045 8412 33057 8415
rect 32456 8384 33057 8412
rect 32456 8372 32462 8384
rect 33045 8381 33057 8384
rect 33091 8381 33103 8415
rect 33045 8375 33103 8381
rect 33226 8372 33232 8424
rect 33284 8412 33290 8424
rect 34057 8415 34115 8421
rect 34057 8412 34069 8415
rect 33284 8384 34069 8412
rect 33284 8372 33290 8384
rect 34057 8381 34069 8384
rect 34103 8381 34115 8415
rect 34057 8375 34115 8381
rect 34606 8372 34612 8424
rect 34664 8372 34670 8424
rect 35158 8372 35164 8424
rect 35216 8372 35222 8424
rect 35710 8372 35716 8424
rect 35768 8412 35774 8424
rect 36909 8415 36967 8421
rect 36909 8412 36921 8415
rect 35768 8384 36921 8412
rect 35768 8372 35774 8384
rect 36909 8381 36921 8384
rect 36955 8412 36967 8415
rect 37553 8415 37611 8421
rect 37553 8412 37565 8415
rect 36955 8384 37565 8412
rect 36955 8381 36967 8384
rect 36909 8375 36967 8381
rect 37553 8381 37565 8384
rect 37599 8381 37611 8415
rect 37553 8375 37611 8381
rect 38841 8415 38899 8421
rect 38841 8381 38853 8415
rect 38887 8412 38899 8415
rect 38933 8415 38991 8421
rect 38933 8412 38945 8415
rect 38887 8384 38945 8412
rect 38887 8381 38899 8384
rect 38841 8375 38899 8381
rect 38933 8381 38945 8384
rect 38979 8412 38991 8415
rect 38979 8384 39344 8412
rect 38979 8381 38991 8384
rect 38933 8375 38991 8381
rect 30926 8304 30932 8356
rect 30984 8344 30990 8356
rect 37001 8347 37059 8353
rect 30984 8316 32996 8344
rect 30984 8304 30990 8316
rect 18969 8279 19027 8285
rect 18969 8276 18981 8279
rect 18064 8248 18981 8276
rect 18969 8245 18981 8248
rect 19015 8245 19027 8279
rect 18969 8239 19027 8245
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 19705 8279 19763 8285
rect 19705 8276 19717 8279
rect 19392 8248 19717 8276
rect 19392 8236 19398 8248
rect 19705 8245 19717 8248
rect 19751 8245 19763 8279
rect 19705 8239 19763 8245
rect 22002 8236 22008 8288
rect 22060 8248 22094 8288
rect 22060 8236 22066 8248
rect 22278 8236 22284 8288
rect 22336 8276 22342 8288
rect 22925 8279 22983 8285
rect 22925 8276 22937 8279
rect 22336 8248 22937 8276
rect 22336 8236 22342 8248
rect 22925 8245 22937 8248
rect 22971 8276 22983 8279
rect 23106 8276 23112 8288
rect 22971 8248 23112 8276
rect 22971 8245 22983 8248
rect 22925 8239 22983 8245
rect 23106 8236 23112 8248
rect 23164 8276 23170 8288
rect 23842 8276 23848 8288
rect 23164 8248 23848 8276
rect 23164 8236 23170 8248
rect 23842 8236 23848 8248
rect 23900 8236 23906 8288
rect 26050 8236 26056 8288
rect 26108 8236 26114 8288
rect 26326 8236 26332 8288
rect 26384 8276 26390 8288
rect 28074 8276 28080 8288
rect 26384 8248 28080 8276
rect 26384 8236 26390 8248
rect 28074 8236 28080 8248
rect 28132 8236 28138 8288
rect 28258 8236 28264 8288
rect 28316 8276 28322 8288
rect 28905 8279 28963 8285
rect 28905 8276 28917 8279
rect 28316 8248 28917 8276
rect 28316 8236 28322 8248
rect 28905 8245 28917 8248
rect 28951 8245 28963 8279
rect 28905 8239 28963 8245
rect 29638 8236 29644 8288
rect 29696 8276 29702 8288
rect 30944 8276 30972 8304
rect 32968 8288 32996 8316
rect 37001 8313 37013 8347
rect 37047 8344 37059 8347
rect 37274 8344 37280 8356
rect 37047 8316 37280 8344
rect 37047 8313 37059 8316
rect 37001 8307 37059 8313
rect 37274 8304 37280 8316
rect 37332 8304 37338 8356
rect 39206 8304 39212 8356
rect 39264 8304 39270 8356
rect 39316 8344 39344 8384
rect 39390 8372 39396 8424
rect 39448 8412 39454 8424
rect 39945 8415 40003 8421
rect 39945 8412 39957 8415
rect 39448 8384 39957 8412
rect 39448 8372 39454 8384
rect 39945 8381 39957 8384
rect 39991 8381 40003 8415
rect 39945 8375 40003 8381
rect 39850 8344 39856 8356
rect 39316 8316 39856 8344
rect 39850 8304 39856 8316
rect 39908 8304 39914 8356
rect 40589 8347 40647 8353
rect 40589 8313 40601 8347
rect 40635 8344 40647 8347
rect 41414 8344 41420 8356
rect 40635 8316 41420 8344
rect 40635 8313 40647 8316
rect 40589 8307 40647 8313
rect 41414 8304 41420 8316
rect 41472 8304 41478 8356
rect 29696 8248 30972 8276
rect 29696 8236 29702 8248
rect 31018 8236 31024 8288
rect 31076 8276 31082 8288
rect 31294 8276 31300 8288
rect 31076 8248 31300 8276
rect 31076 8236 31082 8248
rect 31294 8236 31300 8248
rect 31352 8236 31358 8288
rect 31754 8236 31760 8288
rect 31812 8236 31818 8288
rect 32490 8236 32496 8288
rect 32548 8236 32554 8288
rect 32674 8236 32680 8288
rect 32732 8236 32738 8288
rect 32950 8236 32956 8288
rect 33008 8236 33014 8288
rect 33134 8236 33140 8288
rect 33192 8276 33198 8288
rect 35526 8276 35532 8288
rect 33192 8248 35532 8276
rect 33192 8236 33198 8248
rect 35526 8236 35532 8248
rect 35584 8236 35590 8288
rect 36722 8236 36728 8288
rect 36780 8276 36786 8288
rect 39022 8276 39028 8288
rect 36780 8248 39028 8276
rect 36780 8236 36786 8248
rect 39022 8236 39028 8248
rect 39080 8236 39086 8288
rect 2024 8186 77924 8208
rect 2024 8134 5134 8186
rect 5186 8134 5198 8186
rect 5250 8134 5262 8186
rect 5314 8134 5326 8186
rect 5378 8134 5390 8186
rect 5442 8134 35854 8186
rect 35906 8134 35918 8186
rect 35970 8134 35982 8186
rect 36034 8134 36046 8186
rect 36098 8134 36110 8186
rect 36162 8134 66574 8186
rect 66626 8134 66638 8186
rect 66690 8134 66702 8186
rect 66754 8134 66766 8186
rect 66818 8134 66830 8186
rect 66882 8134 77924 8186
rect 2024 8112 77924 8134
rect 10502 8032 10508 8084
rect 10560 8072 10566 8084
rect 16574 8072 16580 8084
rect 10560 8044 16580 8072
rect 10560 8032 10566 8044
rect 16574 8032 16580 8044
rect 16632 8032 16638 8084
rect 16684 8044 19840 8072
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 12768 7976 15516 8004
rect 12768 7964 12774 7976
rect 15488 7936 15516 7976
rect 15654 7964 15660 8016
rect 15712 7964 15718 8016
rect 16684 8004 16712 8044
rect 16224 7976 16712 8004
rect 17037 8007 17095 8013
rect 16224 7936 16252 7976
rect 17037 7973 17049 8007
rect 17083 8004 17095 8007
rect 19702 8004 19708 8016
rect 17083 7976 19708 8004
rect 17083 7973 17095 7976
rect 17037 7967 17095 7973
rect 19702 7964 19708 7976
rect 19760 7964 19766 8016
rect 19812 8004 19840 8044
rect 19978 8032 19984 8084
rect 20036 8032 20042 8084
rect 20165 8075 20223 8081
rect 20165 8072 20177 8075
rect 20088 8044 20177 8072
rect 20088 8004 20116 8044
rect 20165 8041 20177 8044
rect 20211 8041 20223 8075
rect 20165 8035 20223 8041
rect 20533 8075 20591 8081
rect 20533 8041 20545 8075
rect 20579 8072 20591 8075
rect 21082 8072 21088 8084
rect 20579 8044 21088 8072
rect 20579 8041 20591 8044
rect 20533 8035 20591 8041
rect 21082 8032 21088 8044
rect 21140 8032 21146 8084
rect 21266 8032 21272 8084
rect 21324 8032 21330 8084
rect 24489 8075 24547 8081
rect 24489 8072 24501 8075
rect 22066 8044 24501 8072
rect 19812 7976 20116 8004
rect 20254 7964 20260 8016
rect 20312 8004 20318 8016
rect 22066 8004 22094 8044
rect 24489 8041 24501 8044
rect 24535 8041 24547 8075
rect 24489 8035 24547 8041
rect 25130 8032 25136 8084
rect 25188 8072 25194 8084
rect 25317 8075 25375 8081
rect 25317 8072 25329 8075
rect 25188 8044 25329 8072
rect 25188 8032 25194 8044
rect 25317 8041 25329 8044
rect 25363 8041 25375 8075
rect 25317 8035 25375 8041
rect 25406 8032 25412 8084
rect 25464 8072 25470 8084
rect 25682 8072 25688 8084
rect 25464 8044 25688 8072
rect 25464 8032 25470 8044
rect 25682 8032 25688 8044
rect 25740 8072 25746 8084
rect 27154 8072 27160 8084
rect 25740 8044 27160 8072
rect 25740 8032 25746 8044
rect 27154 8032 27160 8044
rect 27212 8032 27218 8084
rect 27338 8032 27344 8084
rect 27396 8032 27402 8084
rect 29549 8075 29607 8081
rect 29549 8041 29561 8075
rect 29595 8072 29607 8075
rect 29914 8072 29920 8084
rect 29595 8044 29920 8072
rect 29595 8041 29607 8044
rect 29549 8035 29607 8041
rect 29914 8032 29920 8044
rect 29972 8032 29978 8084
rect 31110 8072 31116 8084
rect 30024 8044 31116 8072
rect 20312 7976 22094 8004
rect 20312 7964 20318 7976
rect 23474 7964 23480 8016
rect 23532 8004 23538 8016
rect 23532 7976 24256 8004
rect 23532 7964 23538 7976
rect 15488 7908 16252 7936
rect 16298 7896 16304 7948
rect 16356 7936 16362 7948
rect 16393 7939 16451 7945
rect 16393 7936 16405 7939
rect 16356 7908 16405 7936
rect 16356 7896 16362 7908
rect 16393 7905 16405 7908
rect 16439 7905 16451 7939
rect 16393 7899 16451 7905
rect 16482 7896 16488 7948
rect 16540 7936 16546 7948
rect 17865 7939 17923 7945
rect 17865 7936 17877 7939
rect 16540 7908 17877 7936
rect 16540 7896 16546 7908
rect 17865 7905 17877 7908
rect 17911 7905 17923 7939
rect 17865 7899 17923 7905
rect 18693 7939 18751 7945
rect 18693 7905 18705 7939
rect 18739 7936 18751 7939
rect 18782 7936 18788 7948
rect 18739 7908 18788 7936
rect 18739 7905 18751 7908
rect 18693 7899 18751 7905
rect 18782 7896 18788 7908
rect 18840 7896 18846 7948
rect 21361 7939 21419 7945
rect 21361 7936 21373 7939
rect 18892 7908 21373 7936
rect 14090 7828 14096 7880
rect 14148 7828 14154 7880
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7837 15071 7871
rect 15013 7831 15071 7837
rect 14366 7760 14372 7812
rect 14424 7800 14430 7812
rect 15028 7800 15056 7831
rect 15194 7828 15200 7880
rect 15252 7828 15258 7880
rect 15286 7828 15292 7880
rect 15344 7828 15350 7880
rect 16209 7871 16267 7877
rect 16209 7837 16221 7871
rect 16255 7837 16267 7871
rect 16209 7831 16267 7837
rect 15838 7800 15844 7812
rect 14424 7772 15844 7800
rect 14424 7760 14430 7772
rect 15838 7760 15844 7772
rect 15896 7760 15902 7812
rect 14458 7692 14464 7744
rect 14516 7732 14522 7744
rect 14737 7735 14795 7741
rect 14737 7732 14749 7735
rect 14516 7704 14749 7732
rect 14516 7692 14522 7704
rect 14737 7701 14749 7704
rect 14783 7701 14795 7735
rect 14737 7695 14795 7701
rect 15010 7692 15016 7744
rect 15068 7732 15074 7744
rect 15105 7735 15163 7741
rect 15105 7732 15117 7735
rect 15068 7704 15117 7732
rect 15068 7692 15074 7704
rect 15105 7701 15117 7704
rect 15151 7701 15163 7735
rect 15105 7695 15163 7701
rect 15473 7735 15531 7741
rect 15473 7701 15485 7735
rect 15519 7732 15531 7735
rect 16224 7732 16252 7831
rect 17126 7828 17132 7880
rect 17184 7828 17190 7880
rect 18892 7868 18920 7908
rect 21361 7905 21373 7908
rect 21407 7905 21419 7939
rect 21361 7899 21419 7905
rect 22002 7896 22008 7948
rect 22060 7896 22066 7948
rect 22097 7939 22155 7945
rect 22097 7905 22109 7939
rect 22143 7936 22155 7939
rect 22370 7936 22376 7948
rect 22143 7908 22376 7936
rect 22143 7905 22155 7908
rect 22097 7899 22155 7905
rect 22370 7896 22376 7908
rect 22428 7896 22434 7948
rect 23566 7896 23572 7948
rect 23624 7936 23630 7948
rect 24121 7939 24179 7945
rect 24121 7936 24133 7939
rect 23624 7908 24133 7936
rect 23624 7896 23630 7908
rect 24121 7905 24133 7908
rect 24167 7905 24179 7939
rect 24121 7899 24179 7905
rect 24228 7936 24256 7976
rect 25866 7964 25872 8016
rect 25924 8004 25930 8016
rect 28169 8007 28227 8013
rect 28169 8004 28181 8007
rect 25924 7976 28181 8004
rect 25924 7964 25930 7976
rect 28169 7973 28181 7976
rect 28215 7973 28227 8007
rect 28169 7967 28227 7973
rect 24762 7936 24768 7948
rect 24228 7908 24768 7936
rect 17696 7840 18920 7868
rect 16482 7760 16488 7812
rect 16540 7800 16546 7812
rect 17696 7800 17724 7840
rect 19150 7828 19156 7880
rect 19208 7868 19214 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 19208 7840 19257 7868
rect 19208 7828 19214 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 19426 7828 19432 7880
rect 19484 7828 19490 7880
rect 20162 7828 20168 7880
rect 20220 7828 20226 7880
rect 20254 7828 20260 7880
rect 20312 7828 20318 7880
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7868 20775 7871
rect 21174 7868 21180 7880
rect 20763 7840 21180 7868
rect 20763 7837 20775 7840
rect 20717 7831 20775 7837
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 24228 7877 24256 7908
rect 24762 7896 24768 7908
rect 24820 7896 24826 7948
rect 25133 7939 25191 7945
rect 25133 7905 25145 7939
rect 25179 7936 25191 7939
rect 26050 7936 26056 7948
rect 25179 7908 26056 7936
rect 25179 7905 25191 7908
rect 25133 7899 25191 7905
rect 26050 7896 26056 7908
rect 26108 7896 26114 7948
rect 26789 7939 26847 7945
rect 26789 7905 26801 7939
rect 26835 7936 26847 7939
rect 26878 7936 26884 7948
rect 26835 7908 26884 7936
rect 26835 7905 26847 7908
rect 26789 7899 26847 7905
rect 26878 7896 26884 7908
rect 26936 7896 26942 7948
rect 28813 7939 28871 7945
rect 28813 7905 28825 7939
rect 28859 7936 28871 7939
rect 30024 7936 30052 8044
rect 31110 8032 31116 8044
rect 31168 8032 31174 8084
rect 33686 8032 33692 8084
rect 33744 8072 33750 8084
rect 33744 8044 34376 8072
rect 33744 8032 33750 8044
rect 31754 8004 31760 8016
rect 30300 7976 31760 8004
rect 30300 7945 30328 7976
rect 31754 7964 31760 7976
rect 31812 7964 31818 8016
rect 33410 7964 33416 8016
rect 33468 8004 33474 8016
rect 34241 8007 34299 8013
rect 34241 8004 34253 8007
rect 33468 7976 34253 8004
rect 33468 7964 33474 7976
rect 34241 7973 34253 7976
rect 34287 7973 34299 8007
rect 34348 8004 34376 8044
rect 35158 8032 35164 8084
rect 35216 8072 35222 8084
rect 35437 8075 35495 8081
rect 35437 8072 35449 8075
rect 35216 8044 35449 8072
rect 35216 8032 35222 8044
rect 35437 8041 35449 8044
rect 35483 8041 35495 8075
rect 35437 8035 35495 8041
rect 35544 8044 39620 8072
rect 35544 8004 35572 8044
rect 34348 7976 35572 8004
rect 34241 7967 34299 7973
rect 28859 7908 30052 7936
rect 30285 7939 30343 7945
rect 28859 7905 28871 7908
rect 28813 7899 28871 7905
rect 30285 7905 30297 7939
rect 30331 7905 30343 7939
rect 31662 7936 31668 7948
rect 30285 7899 30343 7905
rect 30392 7908 31668 7936
rect 24213 7871 24271 7877
rect 24213 7837 24225 7871
rect 24259 7837 24271 7871
rect 24213 7831 24271 7837
rect 24397 7871 24455 7877
rect 24397 7837 24409 7871
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 16540 7772 17724 7800
rect 17773 7803 17831 7809
rect 16540 7760 16546 7772
rect 17773 7769 17785 7803
rect 17819 7800 17831 7803
rect 19702 7800 19708 7812
rect 17819 7772 19708 7800
rect 17819 7769 17831 7772
rect 17773 7763 17831 7769
rect 19702 7760 19708 7772
rect 19760 7760 19766 7812
rect 21358 7760 21364 7812
rect 21416 7800 21422 7812
rect 22373 7803 22431 7809
rect 21416 7772 21680 7800
rect 21416 7760 21422 7772
rect 15519 7704 16252 7732
rect 15519 7701 15531 7704
rect 15473 7695 15531 7701
rect 18506 7692 18512 7744
rect 18564 7692 18570 7744
rect 18690 7692 18696 7744
rect 18748 7732 18754 7744
rect 21542 7732 21548 7744
rect 18748 7704 21548 7732
rect 18748 7692 18754 7704
rect 21542 7692 21548 7704
rect 21600 7692 21606 7744
rect 21652 7732 21680 7772
rect 22373 7769 22385 7803
rect 22419 7800 22431 7803
rect 22462 7800 22468 7812
rect 22419 7772 22468 7800
rect 22419 7769 22431 7772
rect 22373 7763 22431 7769
rect 22462 7760 22468 7772
rect 22520 7760 22526 7812
rect 22572 7772 22862 7800
rect 22572 7732 22600 7772
rect 23842 7760 23848 7812
rect 23900 7800 23906 7812
rect 24412 7800 24440 7831
rect 25314 7828 25320 7880
rect 25372 7868 25378 7880
rect 25501 7871 25559 7877
rect 25501 7868 25513 7871
rect 25372 7840 25513 7868
rect 25372 7828 25378 7840
rect 25501 7837 25513 7840
rect 25547 7837 25559 7871
rect 25501 7831 25559 7837
rect 25593 7871 25651 7877
rect 25593 7837 25605 7871
rect 25639 7868 25651 7871
rect 25682 7868 25688 7880
rect 25639 7840 25688 7868
rect 25639 7837 25651 7840
rect 25593 7831 25651 7837
rect 25682 7828 25688 7840
rect 25740 7828 25746 7880
rect 25774 7828 25780 7880
rect 25832 7828 25838 7880
rect 25869 7871 25927 7877
rect 25869 7837 25881 7871
rect 25915 7837 25927 7871
rect 25869 7831 25927 7837
rect 25961 7871 26019 7877
rect 25961 7837 25973 7871
rect 26007 7868 26019 7871
rect 26694 7868 26700 7880
rect 26007 7840 26700 7868
rect 26007 7837 26019 7840
rect 25961 7831 26019 7837
rect 25884 7800 25912 7831
rect 26694 7828 26700 7840
rect 26752 7828 26758 7880
rect 27062 7828 27068 7880
rect 27120 7868 27126 7880
rect 27433 7871 27491 7877
rect 27433 7868 27445 7871
rect 27120 7840 27445 7868
rect 27120 7828 27126 7840
rect 27433 7837 27445 7840
rect 27479 7837 27491 7871
rect 27433 7831 27491 7837
rect 28902 7828 28908 7880
rect 28960 7828 28966 7880
rect 30392 7868 30420 7908
rect 31662 7896 31668 7908
rect 31720 7896 31726 7948
rect 32125 7939 32183 7945
rect 32125 7905 32137 7939
rect 32171 7936 32183 7939
rect 32950 7936 32956 7948
rect 32171 7908 32956 7936
rect 32171 7905 32183 7908
rect 32125 7899 32183 7905
rect 32950 7896 32956 7908
rect 33008 7896 33014 7948
rect 33594 7896 33600 7948
rect 33652 7936 33658 7948
rect 34793 7939 34851 7945
rect 34793 7936 34805 7939
rect 33652 7908 34805 7936
rect 33652 7896 33658 7908
rect 34793 7905 34805 7908
rect 34839 7905 34851 7939
rect 34793 7899 34851 7905
rect 35250 7896 35256 7948
rect 35308 7936 35314 7948
rect 35989 7939 36047 7945
rect 35308 7908 35848 7936
rect 35308 7896 35314 7908
rect 29840 7840 30420 7868
rect 23900 7772 25912 7800
rect 28077 7803 28135 7809
rect 23900 7760 23906 7772
rect 28077 7769 28089 7803
rect 28123 7800 28135 7803
rect 29840 7800 29868 7840
rect 30466 7828 30472 7880
rect 30524 7828 30530 7880
rect 30650 7828 30656 7880
rect 30708 7828 30714 7880
rect 30837 7871 30895 7877
rect 30837 7837 30849 7871
rect 30883 7868 30895 7871
rect 31110 7868 31116 7880
rect 30883 7840 31116 7868
rect 30883 7837 30895 7840
rect 30837 7831 30895 7837
rect 31110 7828 31116 7840
rect 31168 7828 31174 7880
rect 31481 7871 31539 7877
rect 31481 7837 31493 7871
rect 31527 7837 31539 7871
rect 31481 7831 31539 7837
rect 28123 7772 29868 7800
rect 28123 7769 28135 7772
rect 28077 7763 28135 7769
rect 30282 7760 30288 7812
rect 30340 7800 30346 7812
rect 31496 7800 31524 7831
rect 34238 7828 34244 7880
rect 34296 7868 34302 7880
rect 34425 7871 34483 7877
rect 34425 7868 34437 7871
rect 34296 7840 34437 7868
rect 34296 7828 34302 7840
rect 34425 7837 34437 7840
rect 34471 7837 34483 7871
rect 34425 7831 34483 7837
rect 34701 7871 34759 7877
rect 34701 7837 34713 7871
rect 34747 7868 34759 7871
rect 35158 7868 35164 7880
rect 34747 7840 35164 7868
rect 34747 7837 34759 7840
rect 34701 7831 34759 7837
rect 35158 7828 35164 7840
rect 35216 7828 35222 7880
rect 35618 7828 35624 7880
rect 35676 7828 35682 7880
rect 35820 7877 35848 7908
rect 35989 7905 36001 7939
rect 36035 7936 36047 7939
rect 37826 7936 37832 7948
rect 36035 7908 37832 7936
rect 36035 7905 36047 7908
rect 35989 7899 36047 7905
rect 37826 7896 37832 7908
rect 37884 7896 37890 7948
rect 37918 7896 37924 7948
rect 37976 7936 37982 7948
rect 39592 7945 39620 8044
rect 38013 7939 38071 7945
rect 38013 7936 38025 7939
rect 37976 7908 38025 7936
rect 37976 7896 37982 7908
rect 38013 7905 38025 7908
rect 38059 7936 38071 7939
rect 38105 7939 38163 7945
rect 38105 7936 38117 7939
rect 38059 7908 38117 7936
rect 38059 7905 38071 7908
rect 38013 7899 38071 7905
rect 38105 7905 38117 7908
rect 38151 7905 38163 7939
rect 38105 7899 38163 7905
rect 39577 7939 39635 7945
rect 39577 7905 39589 7939
rect 39623 7905 39635 7939
rect 39577 7899 39635 7905
rect 41414 7896 41420 7948
rect 41472 7896 41478 7948
rect 35805 7871 35863 7877
rect 35805 7837 35817 7871
rect 35851 7837 35863 7871
rect 35805 7831 35863 7837
rect 38838 7828 38844 7880
rect 38896 7828 38902 7880
rect 40221 7871 40279 7877
rect 40221 7837 40233 7871
rect 40267 7868 40279 7871
rect 46474 7868 46480 7880
rect 40267 7840 46480 7868
rect 40267 7837 40279 7840
rect 40221 7831 40279 7837
rect 46474 7828 46480 7840
rect 46532 7828 46538 7880
rect 30340 7772 31524 7800
rect 30340 7760 30346 7772
rect 32398 7760 32404 7812
rect 32456 7760 32462 7812
rect 32508 7772 32890 7800
rect 21652 7704 22600 7732
rect 24026 7692 24032 7744
rect 24084 7732 24090 7744
rect 24305 7735 24363 7741
rect 24305 7732 24317 7735
rect 24084 7704 24317 7732
rect 24084 7692 24090 7704
rect 24305 7701 24317 7704
rect 24351 7701 24363 7735
rect 24305 7695 24363 7701
rect 25314 7692 25320 7744
rect 25372 7732 25378 7744
rect 25774 7732 25780 7744
rect 25372 7704 25780 7732
rect 25372 7692 25378 7704
rect 25774 7692 25780 7704
rect 25832 7732 25838 7744
rect 25958 7732 25964 7744
rect 25832 7704 25964 7732
rect 25832 7692 25838 7704
rect 25958 7692 25964 7704
rect 26016 7692 26022 7744
rect 26602 7692 26608 7744
rect 26660 7692 26666 7744
rect 26878 7692 26884 7744
rect 26936 7732 26942 7744
rect 27154 7732 27160 7744
rect 26936 7704 27160 7732
rect 26936 7692 26942 7704
rect 27154 7692 27160 7704
rect 27212 7692 27218 7744
rect 29086 7692 29092 7744
rect 29144 7732 29150 7744
rect 29641 7735 29699 7741
rect 29641 7732 29653 7735
rect 29144 7704 29653 7732
rect 29144 7692 29150 7704
rect 29641 7701 29653 7704
rect 29687 7701 29699 7735
rect 29641 7695 29699 7701
rect 29730 7692 29736 7744
rect 29788 7732 29794 7744
rect 30929 7735 30987 7741
rect 30929 7732 30941 7735
rect 29788 7704 30941 7732
rect 29788 7692 29794 7704
rect 30929 7701 30941 7704
rect 30975 7701 30987 7735
rect 30929 7695 30987 7701
rect 31018 7692 31024 7744
rect 31076 7732 31082 7744
rect 32508 7732 32536 7772
rect 33870 7760 33876 7812
rect 33928 7800 33934 7812
rect 34149 7803 34207 7809
rect 34149 7800 34161 7803
rect 33928 7772 34161 7800
rect 33928 7760 33934 7772
rect 34149 7769 34161 7772
rect 34195 7769 34207 7803
rect 34149 7763 34207 7769
rect 34330 7760 34336 7812
rect 34388 7800 34394 7812
rect 35713 7803 35771 7809
rect 35713 7800 35725 7803
rect 34388 7772 35725 7800
rect 34388 7760 34394 7772
rect 35713 7769 35725 7772
rect 35759 7769 35771 7803
rect 35713 7763 35771 7769
rect 35894 7760 35900 7812
rect 35952 7800 35958 7812
rect 36265 7803 36323 7809
rect 36265 7800 36277 7803
rect 35952 7772 36277 7800
rect 35952 7760 35958 7772
rect 36265 7769 36277 7772
rect 36311 7769 36323 7803
rect 36265 7763 36323 7769
rect 36722 7760 36728 7812
rect 36780 7760 36786 7812
rect 37918 7760 37924 7812
rect 37976 7800 37982 7812
rect 41230 7800 41236 7812
rect 37976 7772 41236 7800
rect 37976 7760 37982 7772
rect 41230 7760 41236 7772
rect 41288 7760 41294 7812
rect 41598 7760 41604 7812
rect 41656 7760 41662 7812
rect 31076 7704 32536 7732
rect 31076 7692 31082 7704
rect 34514 7692 34520 7744
rect 34572 7732 34578 7744
rect 34609 7735 34667 7741
rect 34609 7732 34621 7735
rect 34572 7704 34621 7732
rect 34572 7692 34578 7704
rect 34609 7701 34621 7704
rect 34655 7701 34667 7735
rect 34609 7695 34667 7701
rect 38286 7692 38292 7744
rect 38344 7732 38350 7744
rect 38749 7735 38807 7741
rect 38749 7732 38761 7735
rect 38344 7704 38761 7732
rect 38344 7692 38350 7704
rect 38749 7701 38761 7704
rect 38795 7701 38807 7735
rect 38749 7695 38807 7701
rect 39114 7692 39120 7744
rect 39172 7732 39178 7744
rect 39485 7735 39543 7741
rect 39485 7732 39497 7735
rect 39172 7704 39497 7732
rect 39172 7692 39178 7704
rect 39485 7701 39497 7704
rect 39531 7701 39543 7735
rect 39485 7695 39543 7701
rect 40126 7692 40132 7744
rect 40184 7732 40190 7744
rect 40773 7735 40831 7741
rect 40773 7732 40785 7735
rect 40184 7704 40785 7732
rect 40184 7692 40190 7704
rect 40773 7701 40785 7704
rect 40819 7701 40831 7735
rect 40773 7695 40831 7701
rect 41782 7692 41788 7744
rect 41840 7732 41846 7744
rect 41877 7735 41935 7741
rect 41877 7732 41889 7735
rect 41840 7704 41889 7732
rect 41840 7692 41846 7704
rect 41877 7701 41889 7704
rect 41923 7701 41935 7735
rect 41877 7695 41935 7701
rect 2024 7642 77924 7664
rect 2024 7590 5794 7642
rect 5846 7590 5858 7642
rect 5910 7590 5922 7642
rect 5974 7590 5986 7642
rect 6038 7590 6050 7642
rect 6102 7590 36514 7642
rect 36566 7590 36578 7642
rect 36630 7590 36642 7642
rect 36694 7590 36706 7642
rect 36758 7590 36770 7642
rect 36822 7590 67234 7642
rect 67286 7590 67298 7642
rect 67350 7590 67362 7642
rect 67414 7590 67426 7642
rect 67478 7590 67490 7642
rect 67542 7590 77924 7642
rect 2024 7568 77924 7590
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 15286 7528 15292 7540
rect 11931 7500 15292 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 15930 7488 15936 7540
rect 15988 7488 15994 7540
rect 16114 7488 16120 7540
rect 16172 7528 16178 7540
rect 17589 7531 17647 7537
rect 17589 7528 17601 7531
rect 16172 7500 17601 7528
rect 16172 7488 16178 7500
rect 17589 7497 17601 7500
rect 17635 7497 17647 7531
rect 17589 7491 17647 7497
rect 18598 7488 18604 7540
rect 18656 7528 18662 7540
rect 18877 7531 18935 7537
rect 18877 7528 18889 7531
rect 18656 7500 18889 7528
rect 18656 7488 18662 7500
rect 18877 7497 18889 7500
rect 18923 7497 18935 7531
rect 18877 7491 18935 7497
rect 20990 7488 20996 7540
rect 21048 7528 21054 7540
rect 21085 7531 21143 7537
rect 21085 7528 21097 7531
rect 21048 7500 21097 7528
rect 21048 7488 21054 7500
rect 21085 7497 21097 7500
rect 21131 7497 21143 7531
rect 21085 7491 21143 7497
rect 21174 7488 21180 7540
rect 21232 7488 21238 7540
rect 22278 7528 22284 7540
rect 21744 7500 22284 7528
rect 8938 7420 8944 7472
rect 8996 7460 9002 7472
rect 8996 7432 14596 7460
rect 8996 7420 9002 7432
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 13725 7395 13783 7401
rect 13725 7392 13737 7395
rect 6788 7364 13737 7392
rect 6788 7352 6794 7364
rect 13725 7361 13737 7364
rect 13771 7361 13783 7395
rect 13725 7355 13783 7361
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 9180 7296 11253 7324
rect 9180 7284 9186 7296
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 11241 7287 11299 7293
rect 13354 7284 13360 7336
rect 13412 7284 13418 7336
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 12066 7256 12072 7268
rect 7616 7228 12072 7256
rect 7616 7216 7622 7228
rect 12066 7216 12072 7228
rect 12124 7216 12130 7268
rect 12158 7216 12164 7268
rect 12216 7256 12222 7268
rect 14108 7256 14136 7355
rect 14366 7352 14372 7404
rect 14424 7352 14430 7404
rect 14568 7401 14596 7432
rect 15378 7420 15384 7472
rect 15436 7460 15442 7472
rect 19518 7460 19524 7472
rect 15436 7432 19524 7460
rect 15436 7420 15442 7432
rect 19518 7420 19524 7432
rect 19576 7420 19582 7472
rect 21450 7460 21456 7472
rect 20640 7432 21456 7460
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 14553 7395 14611 7401
rect 14553 7361 14565 7395
rect 14599 7361 14611 7395
rect 14553 7355 14611 7361
rect 14476 7324 14504 7355
rect 15102 7352 15108 7404
rect 15160 7392 15166 7404
rect 16482 7392 16488 7404
rect 15160 7364 16488 7392
rect 15160 7352 15166 7364
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 16574 7352 16580 7404
rect 16632 7352 16638 7404
rect 17402 7352 17408 7404
rect 17460 7352 17466 7404
rect 17773 7395 17831 7401
rect 17773 7361 17785 7395
rect 17819 7361 17831 7395
rect 17773 7355 17831 7361
rect 15194 7324 15200 7336
rect 14476 7296 15200 7324
rect 15194 7284 15200 7296
rect 15252 7284 15258 7336
rect 15286 7284 15292 7336
rect 15344 7284 15350 7336
rect 15378 7284 15384 7336
rect 15436 7324 15442 7336
rect 16025 7327 16083 7333
rect 16025 7324 16037 7327
rect 15436 7296 16037 7324
rect 15436 7284 15442 7296
rect 16025 7293 16037 7296
rect 16071 7293 16083 7327
rect 17788 7324 17816 7355
rect 17862 7352 17868 7404
rect 17920 7352 17926 7404
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7392 18199 7395
rect 19334 7392 19340 7404
rect 18187 7364 19340 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 19334 7352 19340 7364
rect 19392 7352 19398 7404
rect 20162 7352 20168 7404
rect 20220 7392 20226 7404
rect 20640 7401 20668 7432
rect 21450 7420 21456 7432
rect 21508 7420 21514 7472
rect 20441 7395 20499 7401
rect 20441 7392 20453 7395
rect 20220 7364 20453 7392
rect 20220 7352 20226 7364
rect 20441 7361 20453 7364
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 20589 7395 20668 7401
rect 20589 7361 20601 7395
rect 20635 7364 20668 7395
rect 20717 7395 20775 7401
rect 20635 7361 20647 7364
rect 20589 7355 20647 7361
rect 20717 7361 20729 7395
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 16025 7287 16083 7293
rect 16500 7296 17816 7324
rect 18325 7327 18383 7333
rect 16500 7268 16528 7296
rect 18325 7293 18337 7327
rect 18371 7324 18383 7327
rect 18782 7324 18788 7336
rect 18371 7296 18788 7324
rect 18371 7293 18383 7296
rect 18325 7287 18383 7293
rect 18782 7284 18788 7296
rect 18840 7284 18846 7336
rect 18966 7284 18972 7336
rect 19024 7284 19030 7336
rect 19705 7327 19763 7333
rect 19705 7293 19717 7327
rect 19751 7293 19763 7327
rect 20732 7324 20760 7355
rect 20806 7352 20812 7404
rect 20864 7352 20870 7404
rect 20947 7395 21005 7401
rect 20947 7361 20959 7395
rect 20993 7392 21005 7395
rect 21744 7392 21772 7500
rect 22278 7488 22284 7500
rect 22336 7488 22342 7540
rect 22557 7531 22615 7537
rect 22557 7497 22569 7531
rect 22603 7528 22615 7531
rect 24302 7528 24308 7540
rect 22603 7500 24308 7528
rect 22603 7497 22615 7500
rect 22557 7491 22615 7497
rect 24302 7488 24308 7500
rect 24360 7488 24366 7540
rect 24949 7531 25007 7537
rect 24949 7497 24961 7531
rect 24995 7528 25007 7531
rect 27614 7528 27620 7540
rect 24995 7500 27620 7528
rect 24995 7497 25007 7500
rect 24949 7491 25007 7497
rect 27614 7488 27620 7500
rect 27672 7488 27678 7540
rect 27709 7531 27767 7537
rect 27709 7497 27721 7531
rect 27755 7528 27767 7531
rect 28902 7528 28908 7540
rect 27755 7500 28908 7528
rect 27755 7497 27767 7500
rect 27709 7491 27767 7497
rect 28902 7488 28908 7500
rect 28960 7488 28966 7540
rect 30098 7488 30104 7540
rect 30156 7528 30162 7540
rect 30926 7528 30932 7540
rect 30156 7500 30932 7528
rect 30156 7488 30162 7500
rect 22462 7460 22468 7472
rect 22020 7432 22468 7460
rect 22020 7401 22048 7432
rect 22462 7420 22468 7432
rect 22520 7420 22526 7472
rect 24762 7420 24768 7472
rect 24820 7460 24826 7472
rect 25317 7463 25375 7469
rect 25317 7460 25329 7463
rect 24820 7432 25329 7460
rect 24820 7420 24826 7432
rect 25317 7429 25329 7432
rect 25363 7429 25375 7463
rect 25317 7423 25375 7429
rect 26878 7420 26884 7472
rect 26936 7460 26942 7472
rect 27065 7463 27123 7469
rect 27065 7460 27077 7463
rect 26936 7432 27077 7460
rect 26936 7420 26942 7432
rect 27065 7429 27077 7432
rect 27111 7429 27123 7463
rect 27065 7423 27123 7429
rect 27433 7463 27491 7469
rect 27433 7429 27445 7463
rect 27479 7460 27491 7463
rect 28258 7460 28264 7472
rect 27479 7432 28264 7460
rect 27479 7429 27491 7432
rect 27433 7423 27491 7429
rect 28258 7420 28264 7432
rect 28316 7420 28322 7472
rect 28813 7463 28871 7469
rect 28813 7429 28825 7463
rect 28859 7460 28871 7463
rect 30009 7463 30067 7469
rect 30009 7460 30021 7463
rect 28859 7432 30021 7460
rect 28859 7429 28871 7432
rect 28813 7423 28871 7429
rect 30009 7429 30021 7432
rect 30055 7429 30067 7463
rect 30395 7460 30423 7500
rect 30926 7488 30932 7500
rect 30984 7488 30990 7540
rect 31018 7488 31024 7540
rect 31076 7528 31082 7540
rect 31076 7500 32168 7528
rect 31076 7488 31082 7500
rect 30395 7432 30498 7460
rect 30009 7423 30067 7429
rect 31754 7420 31760 7472
rect 31812 7420 31818 7472
rect 32140 7460 32168 7500
rect 32214 7488 32220 7540
rect 32272 7488 32278 7540
rect 33965 7531 34023 7537
rect 32324 7500 33088 7528
rect 32324 7460 32352 7500
rect 32140 7432 32352 7460
rect 32398 7420 32404 7472
rect 32456 7420 32462 7472
rect 32674 7420 32680 7472
rect 32732 7460 32738 7472
rect 32858 7460 32864 7472
rect 32732 7432 32864 7460
rect 32732 7420 32738 7432
rect 32858 7420 32864 7432
rect 32916 7420 32922 7472
rect 20993 7364 21772 7392
rect 21821 7395 21879 7401
rect 20993 7361 21005 7364
rect 20947 7355 21005 7361
rect 21821 7361 21833 7395
rect 21867 7392 21879 7395
rect 22005 7395 22063 7401
rect 21867 7364 21968 7392
rect 21867 7361 21879 7364
rect 21821 7355 21879 7361
rect 21174 7324 21180 7336
rect 20732 7296 21180 7324
rect 19705 7287 19763 7293
rect 12216 7228 14136 7256
rect 12216 7216 12222 7228
rect 14826 7216 14832 7268
rect 14884 7256 14890 7268
rect 16114 7256 16120 7268
rect 14884 7228 16120 7256
rect 14884 7216 14890 7228
rect 16114 7216 16120 7228
rect 16172 7216 16178 7268
rect 16482 7216 16488 7268
rect 16540 7216 16546 7268
rect 16758 7216 16764 7268
rect 16816 7216 16822 7268
rect 17678 7216 17684 7268
rect 17736 7256 17742 7268
rect 19720 7256 19748 7287
rect 21174 7284 21180 7296
rect 21232 7284 21238 7336
rect 21940 7324 21968 7364
rect 22005 7361 22017 7395
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22370 7352 22376 7404
rect 22428 7392 22434 7404
rect 23474 7392 23480 7404
rect 22428 7364 23480 7392
rect 22428 7352 22434 7364
rect 23474 7352 23480 7364
rect 23532 7392 23538 7404
rect 25041 7395 25099 7401
rect 25041 7392 25053 7395
rect 23532 7364 25053 7392
rect 23532 7352 23538 7364
rect 25041 7361 25053 7364
rect 25087 7361 25099 7395
rect 25041 7355 25099 7361
rect 23201 7327 23259 7333
rect 23201 7324 23213 7327
rect 21940 7296 23213 7324
rect 23201 7293 23213 7296
rect 23247 7293 23259 7327
rect 23201 7287 23259 7293
rect 23566 7284 23572 7336
rect 23624 7324 23630 7336
rect 23750 7324 23756 7336
rect 23624 7296 23756 7324
rect 23624 7284 23630 7296
rect 23750 7284 23756 7296
rect 23808 7284 23814 7336
rect 24305 7327 24363 7333
rect 24305 7293 24317 7327
rect 24351 7293 24363 7327
rect 25056 7324 25084 7355
rect 26418 7352 26424 7404
rect 26476 7352 26482 7404
rect 26896 7392 26924 7420
rect 26528 7364 26924 7392
rect 26528 7336 26556 7364
rect 27154 7352 27160 7404
rect 27212 7352 27218 7404
rect 27341 7395 27399 7401
rect 27341 7361 27353 7395
rect 27387 7392 27399 7395
rect 27525 7395 27583 7401
rect 27387 7364 27476 7392
rect 27387 7361 27399 7364
rect 27341 7355 27399 7361
rect 25958 7324 25964 7336
rect 25056 7296 25964 7324
rect 24305 7287 24363 7293
rect 20990 7256 20996 7268
rect 17736 7228 19748 7256
rect 20272 7228 20996 7256
rect 17736 7216 17742 7228
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 9732 7160 12817 7188
rect 9732 7148 9738 7160
rect 12805 7157 12817 7160
rect 12851 7157 12863 7191
rect 12805 7151 12863 7157
rect 13538 7148 13544 7200
rect 13596 7148 13602 7200
rect 15197 7191 15255 7197
rect 15197 7157 15209 7191
rect 15243 7188 15255 7191
rect 15930 7188 15936 7200
rect 15243 7160 15936 7188
rect 15243 7157 15255 7160
rect 15197 7151 15255 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 18049 7191 18107 7197
rect 18049 7157 18061 7191
rect 18095 7188 18107 7191
rect 18598 7188 18604 7200
rect 18095 7160 18604 7188
rect 18095 7157 18107 7160
rect 18049 7151 18107 7157
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 19613 7191 19671 7197
rect 19613 7157 19625 7191
rect 19659 7188 19671 7191
rect 20272 7188 20300 7228
rect 20990 7216 20996 7228
rect 21048 7216 21054 7268
rect 21542 7216 21548 7268
rect 21600 7256 21606 7268
rect 24320 7256 24348 7287
rect 25958 7284 25964 7296
rect 26016 7284 26022 7336
rect 26510 7284 26516 7336
rect 26568 7284 26574 7336
rect 21600 7228 21772 7256
rect 21600 7216 21606 7228
rect 19659 7160 20300 7188
rect 20349 7191 20407 7197
rect 19659 7157 19671 7160
rect 19613 7151 19671 7157
rect 20349 7157 20361 7191
rect 20395 7188 20407 7191
rect 20806 7188 20812 7200
rect 20395 7160 20812 7188
rect 20395 7157 20407 7160
rect 20349 7151 20407 7157
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 21744 7188 21772 7228
rect 23308 7228 24348 7256
rect 27448 7256 27476 7364
rect 27525 7361 27537 7395
rect 27571 7392 27583 7395
rect 27890 7392 27896 7404
rect 27571 7364 27896 7392
rect 27571 7361 27583 7364
rect 27525 7355 27583 7361
rect 27890 7352 27896 7364
rect 27948 7352 27954 7404
rect 29638 7352 29644 7404
rect 29696 7392 29702 7404
rect 29733 7395 29791 7401
rect 29733 7392 29745 7395
rect 29696 7364 29745 7392
rect 29696 7352 29702 7364
rect 29733 7361 29745 7364
rect 29779 7361 29791 7395
rect 29733 7355 29791 7361
rect 31662 7352 31668 7404
rect 31720 7392 31726 7404
rect 31849 7395 31907 7401
rect 31849 7392 31861 7395
rect 31720 7364 31861 7392
rect 31720 7352 31726 7364
rect 31849 7361 31861 7364
rect 31895 7361 31907 7395
rect 31849 7355 31907 7361
rect 31938 7352 31944 7404
rect 31996 7352 32002 7404
rect 32125 7395 32183 7401
rect 32125 7361 32137 7395
rect 32171 7392 32183 7395
rect 32214 7392 32220 7404
rect 32171 7364 32220 7392
rect 32171 7361 32183 7364
rect 32125 7355 32183 7361
rect 32214 7352 32220 7364
rect 32272 7352 32278 7404
rect 32416 7392 32444 7420
rect 32324 7364 32444 7392
rect 32493 7395 32551 7401
rect 28261 7327 28319 7333
rect 28261 7293 28273 7327
rect 28307 7324 28319 7327
rect 28350 7324 28356 7336
rect 28307 7296 28356 7324
rect 28307 7293 28319 7296
rect 28261 7287 28319 7293
rect 28350 7284 28356 7296
rect 28408 7284 28414 7336
rect 28810 7284 28816 7336
rect 28868 7324 28874 7336
rect 28905 7327 28963 7333
rect 28905 7324 28917 7327
rect 28868 7296 28917 7324
rect 28868 7284 28874 7296
rect 28905 7293 28917 7296
rect 28951 7293 28963 7327
rect 28905 7287 28963 7293
rect 29549 7327 29607 7333
rect 29549 7293 29561 7327
rect 29595 7324 29607 7327
rect 30466 7324 30472 7336
rect 29595 7296 30472 7324
rect 29595 7293 29607 7296
rect 29549 7287 29607 7293
rect 30466 7284 30472 7296
rect 30524 7284 30530 7336
rect 31018 7284 31024 7336
rect 31076 7324 31082 7336
rect 31570 7324 31576 7336
rect 31076 7296 31576 7324
rect 31076 7284 31082 7296
rect 31570 7284 31576 7296
rect 31628 7324 31634 7336
rect 32324 7324 32352 7364
rect 32493 7361 32505 7395
rect 32539 7392 32551 7395
rect 32582 7392 32588 7404
rect 32539 7364 32588 7392
rect 32539 7361 32551 7364
rect 32493 7355 32551 7361
rect 32582 7352 32588 7364
rect 32640 7352 32646 7404
rect 33060 7401 33088 7500
rect 33965 7497 33977 7531
rect 34011 7528 34023 7531
rect 34606 7528 34612 7540
rect 34011 7500 34612 7528
rect 34011 7497 34023 7500
rect 33965 7491 34023 7497
rect 34606 7488 34612 7500
rect 34664 7488 34670 7540
rect 34885 7531 34943 7537
rect 34885 7497 34897 7531
rect 34931 7528 34943 7531
rect 34974 7528 34980 7540
rect 34931 7500 34980 7528
rect 34931 7497 34943 7500
rect 34885 7491 34943 7497
rect 34974 7488 34980 7500
rect 35032 7488 35038 7540
rect 35250 7488 35256 7540
rect 35308 7488 35314 7540
rect 35526 7488 35532 7540
rect 35584 7488 35590 7540
rect 35894 7488 35900 7540
rect 35952 7488 35958 7540
rect 36446 7488 36452 7540
rect 36504 7528 36510 7540
rect 36504 7500 38148 7528
rect 36504 7488 36510 7500
rect 34422 7420 34428 7472
rect 34480 7460 34486 7472
rect 35069 7463 35127 7469
rect 35069 7460 35081 7463
rect 34480 7432 35081 7460
rect 34480 7420 34486 7432
rect 35069 7429 35081 7432
rect 35115 7460 35127 7463
rect 35268 7460 35296 7488
rect 35437 7463 35495 7469
rect 35437 7460 35449 7463
rect 35115 7432 35204 7460
rect 35268 7432 35449 7460
rect 35115 7429 35127 7432
rect 35069 7423 35127 7429
rect 33045 7395 33103 7401
rect 33045 7361 33057 7395
rect 33091 7361 33103 7395
rect 33045 7355 33103 7361
rect 33134 7352 33140 7404
rect 33192 7392 33198 7404
rect 33229 7395 33287 7401
rect 33229 7392 33241 7395
rect 33192 7364 33241 7392
rect 33192 7352 33198 7364
rect 33229 7361 33241 7364
rect 33275 7361 33287 7395
rect 33229 7355 33287 7361
rect 33870 7352 33876 7404
rect 33928 7392 33934 7404
rect 34609 7395 34667 7401
rect 34609 7392 34621 7395
rect 33928 7364 34621 7392
rect 33928 7352 33934 7364
rect 34609 7361 34621 7364
rect 34655 7361 34667 7395
rect 34609 7355 34667 7361
rect 34790 7352 34796 7404
rect 34848 7352 34854 7404
rect 35176 7401 35204 7432
rect 35437 7429 35449 7432
rect 35483 7429 35495 7463
rect 35437 7423 35495 7429
rect 35161 7395 35219 7401
rect 35161 7361 35173 7395
rect 35207 7361 35219 7395
rect 35161 7355 35219 7361
rect 35253 7395 35311 7401
rect 35253 7361 35265 7395
rect 35299 7392 35311 7395
rect 35342 7392 35348 7404
rect 35299 7364 35348 7392
rect 35299 7361 35311 7364
rect 35253 7355 35311 7361
rect 35342 7352 35348 7364
rect 35400 7352 35406 7404
rect 35544 7401 35572 7488
rect 38010 7460 38016 7472
rect 36556 7432 38016 7460
rect 35529 7395 35587 7401
rect 35529 7361 35541 7395
rect 35575 7361 35587 7395
rect 35529 7355 35587 7361
rect 35621 7395 35679 7401
rect 35621 7361 35633 7395
rect 35667 7392 35679 7395
rect 35710 7392 35716 7404
rect 35667 7364 35716 7392
rect 35667 7361 35679 7364
rect 35621 7355 35679 7361
rect 35710 7352 35716 7364
rect 35768 7352 35774 7404
rect 36556 7401 36584 7432
rect 38010 7420 38016 7432
rect 38068 7420 38074 7472
rect 38120 7460 38148 7500
rect 40034 7488 40040 7540
rect 40092 7528 40098 7540
rect 42061 7531 42119 7537
rect 42061 7528 42073 7531
rect 40092 7500 42073 7528
rect 40092 7488 40098 7500
rect 42061 7497 42073 7500
rect 42107 7497 42119 7531
rect 42061 7491 42119 7497
rect 38120 7432 41184 7460
rect 36541 7395 36599 7401
rect 36541 7361 36553 7395
rect 36587 7361 36599 7395
rect 36541 7355 36599 7361
rect 37274 7352 37280 7404
rect 37332 7352 37338 7404
rect 38286 7352 38292 7404
rect 38344 7352 38350 7404
rect 41156 7401 41184 7432
rect 41230 7420 41236 7472
rect 41288 7460 41294 7472
rect 41288 7432 41414 7460
rect 41288 7420 41294 7432
rect 40221 7395 40279 7401
rect 40221 7392 40233 7395
rect 38396 7364 40233 7392
rect 31628 7296 32352 7324
rect 32401 7327 32459 7333
rect 31628 7284 31634 7296
rect 32401 7293 32413 7327
rect 32447 7293 32459 7327
rect 32401 7287 32459 7293
rect 28994 7256 29000 7268
rect 27448 7228 29000 7256
rect 23308 7188 23336 7228
rect 28994 7216 29000 7228
rect 29052 7216 29058 7268
rect 32125 7259 32183 7265
rect 32125 7225 32137 7259
rect 32171 7225 32183 7259
rect 32416 7256 32444 7287
rect 32766 7284 32772 7336
rect 32824 7284 32830 7336
rect 32861 7327 32919 7333
rect 32861 7293 32873 7327
rect 32907 7293 32919 7327
rect 32861 7287 32919 7293
rect 33413 7327 33471 7333
rect 33413 7293 33425 7327
rect 33459 7324 33471 7327
rect 34057 7327 34115 7333
rect 34057 7324 34069 7327
rect 33459 7296 34069 7324
rect 33459 7293 33471 7296
rect 33413 7287 33471 7293
rect 34057 7293 34069 7296
rect 34103 7293 34115 7327
rect 34057 7287 34115 7293
rect 32125 7219 32183 7225
rect 32324 7228 32444 7256
rect 32876 7256 32904 7287
rect 34974 7284 34980 7336
rect 35032 7324 35038 7336
rect 37369 7327 37427 7333
rect 37369 7324 37381 7327
rect 35032 7296 37381 7324
rect 35032 7284 35038 7296
rect 37369 7293 37381 7296
rect 37415 7293 37427 7327
rect 38396 7324 38424 7364
rect 40221 7361 40233 7364
rect 40267 7361 40279 7395
rect 40221 7355 40279 7361
rect 41141 7395 41199 7401
rect 41141 7361 41153 7395
rect 41187 7361 41199 7395
rect 41386 7392 41414 7432
rect 42613 7395 42671 7401
rect 42613 7392 42625 7395
rect 41386 7364 42625 7392
rect 41141 7355 41199 7361
rect 42613 7361 42625 7364
rect 42659 7361 42671 7395
rect 42613 7355 42671 7361
rect 37369 7287 37427 7293
rect 37476 7296 38424 7324
rect 38841 7327 38899 7333
rect 33042 7256 33048 7268
rect 32876 7228 33048 7256
rect 21744 7160 23336 7188
rect 23382 7148 23388 7200
rect 23440 7188 23446 7200
rect 23566 7188 23572 7200
rect 23440 7160 23572 7188
rect 23440 7148 23446 7160
rect 23566 7148 23572 7160
rect 23624 7148 23630 7200
rect 26050 7148 26056 7200
rect 26108 7188 26114 7200
rect 30650 7188 30656 7200
rect 26108 7160 30656 7188
rect 26108 7148 26114 7160
rect 30650 7148 30656 7160
rect 30708 7148 30714 7200
rect 32140 7188 32168 7219
rect 32324 7188 32352 7228
rect 33042 7216 33048 7228
rect 33100 7216 33106 7268
rect 37090 7216 37096 7268
rect 37148 7256 37154 7268
rect 37476 7256 37504 7296
rect 38841 7293 38853 7327
rect 38887 7324 38899 7327
rect 39485 7327 39543 7333
rect 39485 7324 39497 7327
rect 38887 7296 39497 7324
rect 38887 7293 38899 7296
rect 38841 7287 38899 7293
rect 39485 7293 39497 7296
rect 39531 7293 39543 7327
rect 39485 7287 39543 7293
rect 41417 7327 41475 7333
rect 41417 7293 41429 7327
rect 41463 7324 41475 7327
rect 41598 7324 41604 7336
rect 41463 7296 41604 7324
rect 41463 7293 41475 7296
rect 41417 7287 41475 7293
rect 41598 7284 41604 7296
rect 41656 7284 41662 7336
rect 37148 7228 37504 7256
rect 37148 7216 37154 7228
rect 38102 7216 38108 7268
rect 38160 7256 38166 7268
rect 39669 7259 39727 7265
rect 39669 7256 39681 7259
rect 38160 7228 39681 7256
rect 38160 7216 38166 7228
rect 39669 7225 39681 7228
rect 39715 7225 39727 7259
rect 39669 7219 39727 7225
rect 32140 7160 32352 7188
rect 32398 7148 32404 7200
rect 32456 7188 32462 7200
rect 33137 7191 33195 7197
rect 33137 7188 33149 7191
rect 32456 7160 33149 7188
rect 32456 7148 32462 7160
rect 33137 7157 33149 7160
rect 33183 7157 33195 7191
rect 33137 7151 33195 7157
rect 35066 7148 35072 7200
rect 35124 7148 35130 7200
rect 35434 7148 35440 7200
rect 35492 7188 35498 7200
rect 35805 7191 35863 7197
rect 35805 7188 35817 7191
rect 35492 7160 35817 7188
rect 35492 7148 35498 7160
rect 35805 7157 35817 7160
rect 35851 7157 35863 7191
rect 35805 7151 35863 7157
rect 36538 7148 36544 7200
rect 36596 7188 36602 7200
rect 36633 7191 36691 7197
rect 36633 7188 36645 7191
rect 36596 7160 36645 7188
rect 36596 7148 36602 7160
rect 36633 7157 36645 7160
rect 36679 7157 36691 7191
rect 36633 7151 36691 7157
rect 37918 7148 37924 7200
rect 37976 7188 37982 7200
rect 38013 7191 38071 7197
rect 38013 7188 38025 7191
rect 37976 7160 38025 7188
rect 37976 7148 37982 7160
rect 38013 7157 38025 7160
rect 38059 7157 38071 7191
rect 38013 7151 38071 7157
rect 38930 7148 38936 7200
rect 38988 7148 38994 7200
rect 40586 7148 40592 7200
rect 40644 7148 40650 7200
rect 41969 7191 42027 7197
rect 41969 7157 41981 7191
rect 42015 7188 42027 7191
rect 42150 7188 42156 7200
rect 42015 7160 42156 7188
rect 42015 7157 42027 7160
rect 41969 7151 42027 7157
rect 42150 7148 42156 7160
rect 42208 7148 42214 7200
rect 2024 7098 77924 7120
rect 2024 7046 5134 7098
rect 5186 7046 5198 7098
rect 5250 7046 5262 7098
rect 5314 7046 5326 7098
rect 5378 7046 5390 7098
rect 5442 7046 35854 7098
rect 35906 7046 35918 7098
rect 35970 7046 35982 7098
rect 36034 7046 36046 7098
rect 36098 7046 36110 7098
rect 36162 7046 66574 7098
rect 66626 7046 66638 7098
rect 66690 7046 66702 7098
rect 66754 7046 66766 7098
rect 66818 7046 66830 7098
rect 66882 7046 77924 7098
rect 2024 7024 77924 7046
rect 10042 6944 10048 6996
rect 10100 6984 10106 6996
rect 13538 6984 13544 6996
rect 10100 6956 13544 6984
rect 10100 6944 10106 6956
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 16669 6987 16727 6993
rect 16669 6953 16681 6987
rect 16715 6984 16727 6987
rect 17862 6984 17868 6996
rect 16715 6956 17868 6984
rect 16715 6953 16727 6956
rect 16669 6947 16727 6953
rect 17862 6944 17868 6956
rect 17920 6944 17926 6996
rect 18966 6944 18972 6996
rect 19024 6944 19030 6996
rect 20898 6944 20904 6996
rect 20956 6984 20962 6996
rect 21925 6987 21983 6993
rect 21925 6984 21937 6987
rect 20956 6956 21937 6984
rect 20956 6944 20962 6956
rect 21925 6953 21937 6956
rect 21971 6953 21983 6987
rect 21925 6947 21983 6953
rect 22465 6987 22523 6993
rect 22465 6953 22477 6987
rect 22511 6984 22523 6987
rect 22922 6984 22928 6996
rect 22511 6956 22928 6984
rect 22511 6953 22523 6956
rect 22465 6947 22523 6953
rect 22922 6944 22928 6956
rect 22980 6984 22986 6996
rect 23750 6984 23756 6996
rect 22980 6956 23756 6984
rect 22980 6944 22986 6956
rect 23750 6944 23756 6956
rect 23808 6944 23814 6996
rect 24026 6944 24032 6996
rect 24084 6984 24090 6996
rect 25869 6987 25927 6993
rect 25869 6984 25881 6987
rect 24084 6956 25881 6984
rect 24084 6944 24090 6956
rect 25869 6953 25881 6956
rect 25915 6984 25927 6987
rect 26050 6984 26056 6996
rect 25915 6956 26056 6984
rect 25915 6953 25927 6956
rect 25869 6947 25927 6953
rect 26050 6944 26056 6956
rect 26108 6944 26114 6996
rect 26602 6944 26608 6996
rect 26660 6984 26666 6996
rect 26954 6987 27012 6993
rect 26954 6984 26966 6987
rect 26660 6956 26966 6984
rect 26660 6944 26666 6956
rect 26954 6953 26966 6956
rect 27000 6953 27012 6987
rect 26954 6947 27012 6953
rect 28994 6944 29000 6996
rect 29052 6984 29058 6996
rect 35066 6984 35072 6996
rect 29052 6956 35072 6984
rect 29052 6944 29058 6956
rect 35066 6944 35072 6956
rect 35124 6944 35130 6996
rect 37724 6987 37782 6993
rect 37724 6953 37736 6987
rect 37770 6984 37782 6987
rect 37918 6984 37924 6996
rect 37770 6956 37924 6984
rect 37770 6953 37782 6956
rect 37724 6947 37782 6953
rect 37918 6944 37924 6956
rect 37976 6944 37982 6996
rect 13630 6876 13636 6928
rect 13688 6916 13694 6928
rect 13688 6888 15056 6916
rect 13688 6876 13694 6888
rect 6362 6808 6368 6860
rect 6420 6848 6426 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 6420 6820 11989 6848
rect 6420 6808 6426 6820
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 13357 6851 13415 6857
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 14734 6848 14740 6860
rect 13403 6820 14740 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 14826 6808 14832 6860
rect 14884 6808 14890 6860
rect 15028 6848 15056 6888
rect 15838 6876 15844 6928
rect 15896 6916 15902 6928
rect 19058 6916 19064 6928
rect 15896 6888 19064 6916
rect 15896 6876 15902 6888
rect 19058 6876 19064 6888
rect 19116 6876 19122 6928
rect 22112 6888 22508 6916
rect 15286 6848 15292 6860
rect 15028 6820 15292 6848
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 11149 6783 11207 6789
rect 11149 6780 11161 6783
rect 6696 6752 11161 6780
rect 6696 6740 6702 6752
rect 11149 6749 11161 6752
rect 11195 6749 11207 6783
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 11149 6743 11207 6749
rect 11256 6752 12725 6780
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 11256 6712 11284 6752
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6780 14151 6783
rect 14642 6780 14648 6792
rect 14139 6752 14648 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 14642 6740 14648 6752
rect 14700 6740 14706 6792
rect 15028 6789 15056 6820
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 17405 6851 17463 6857
rect 17405 6817 17417 6851
rect 17451 6848 17463 6851
rect 19426 6848 19432 6860
rect 17451 6820 19432 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 20438 6848 20444 6860
rect 20180 6820 20444 6848
rect 15013 6783 15071 6789
rect 15013 6749 15025 6783
rect 15059 6749 15071 6783
rect 15013 6743 15071 6749
rect 15197 6783 15255 6789
rect 15197 6749 15209 6783
rect 15243 6780 15255 6783
rect 15470 6780 15476 6792
rect 15243 6752 15476 6780
rect 15243 6749 15255 6752
rect 15197 6743 15255 6749
rect 15470 6740 15476 6752
rect 15528 6780 15534 6792
rect 15746 6780 15752 6792
rect 15528 6752 15752 6780
rect 15528 6740 15534 6752
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 8720 6684 11284 6712
rect 8720 6672 8726 6684
rect 11514 6672 11520 6724
rect 11572 6712 11578 6724
rect 15856 6712 15884 6743
rect 16114 6740 16120 6792
rect 16172 6740 16178 6792
rect 16853 6783 16911 6789
rect 16853 6749 16865 6783
rect 16899 6749 16911 6783
rect 16853 6743 16911 6749
rect 11572 6684 15884 6712
rect 16868 6712 16896 6743
rect 17494 6740 17500 6792
rect 17552 6740 17558 6792
rect 18138 6740 18144 6792
rect 18196 6780 18202 6792
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 18196 6752 18245 6780
rect 18196 6740 18202 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 18782 6740 18788 6792
rect 18840 6740 18846 6792
rect 19518 6740 19524 6792
rect 19576 6740 19582 6792
rect 20180 6721 20208 6820
rect 20438 6808 20444 6820
rect 20496 6848 20502 6860
rect 22112 6848 22140 6888
rect 20496 6820 22140 6848
rect 22189 6851 22247 6857
rect 20496 6808 20502 6820
rect 22189 6817 22201 6851
rect 22235 6848 22247 6851
rect 22370 6848 22376 6860
rect 22235 6820 22376 6848
rect 22235 6817 22247 6820
rect 22189 6811 22247 6817
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 22480 6848 22508 6888
rect 23382 6876 23388 6928
rect 23440 6916 23446 6928
rect 25317 6919 25375 6925
rect 25317 6916 25329 6919
rect 23440 6888 25329 6916
rect 23440 6876 23446 6888
rect 25317 6885 25329 6888
rect 25363 6916 25375 6919
rect 25406 6916 25412 6928
rect 25363 6888 25412 6916
rect 25363 6885 25375 6888
rect 25317 6879 25375 6885
rect 25406 6876 25412 6888
rect 25464 6876 25470 6928
rect 25958 6876 25964 6928
rect 26016 6916 26022 6928
rect 26016 6888 26740 6916
rect 26016 6876 26022 6888
rect 23661 6851 23719 6857
rect 22480 6820 22692 6848
rect 22554 6740 22560 6792
rect 22612 6740 22618 6792
rect 20165 6715 20223 6721
rect 20165 6712 20177 6715
rect 16868 6684 20177 6712
rect 11572 6672 11578 6684
rect 20165 6681 20177 6684
rect 20211 6681 20223 6715
rect 20165 6675 20223 6681
rect 21358 6672 21364 6724
rect 21416 6672 21422 6724
rect 22449 6715 22507 6721
rect 22449 6681 22461 6715
rect 22495 6712 22507 6715
rect 22572 6712 22600 6740
rect 22664 6724 22692 6820
rect 23661 6817 23673 6851
rect 23707 6848 23719 6851
rect 23934 6848 23940 6860
rect 23707 6820 23940 6848
rect 23707 6817 23719 6820
rect 23661 6811 23719 6817
rect 23934 6808 23940 6820
rect 23992 6808 23998 6860
rect 24581 6851 24639 6857
rect 24581 6817 24593 6851
rect 24627 6848 24639 6851
rect 24854 6848 24860 6860
rect 24627 6820 24860 6848
rect 24627 6817 24639 6820
rect 24581 6811 24639 6817
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 24964 6820 26004 6848
rect 23477 6783 23535 6789
rect 23477 6749 23489 6783
rect 23523 6780 23535 6783
rect 24964 6780 24992 6820
rect 23523 6752 24992 6780
rect 23523 6749 23535 6752
rect 23477 6743 23535 6749
rect 25498 6740 25504 6792
rect 25556 6740 25562 6792
rect 25682 6740 25688 6792
rect 25740 6740 25746 6792
rect 25976 6789 26004 6820
rect 26510 6808 26516 6860
rect 26568 6808 26574 6860
rect 26712 6857 26740 6888
rect 30282 6876 30288 6928
rect 30340 6876 30346 6928
rect 30374 6876 30380 6928
rect 30432 6916 30438 6928
rect 31662 6916 31668 6928
rect 30432 6888 31668 6916
rect 30432 6876 30438 6888
rect 31662 6876 31668 6888
rect 31720 6916 31726 6928
rect 33870 6916 33876 6928
rect 31720 6888 33876 6916
rect 31720 6876 31726 6888
rect 33870 6876 33876 6888
rect 33928 6876 33934 6928
rect 34606 6876 34612 6928
rect 34664 6916 34670 6928
rect 35158 6916 35164 6928
rect 34664 6888 35164 6916
rect 34664 6876 34670 6888
rect 35158 6876 35164 6888
rect 35216 6916 35222 6928
rect 35710 6916 35716 6928
rect 35216 6888 35716 6916
rect 35216 6876 35222 6888
rect 35710 6876 35716 6888
rect 35768 6876 35774 6928
rect 26697 6851 26755 6857
rect 26697 6817 26709 6851
rect 26743 6817 26755 6851
rect 26697 6811 26755 6817
rect 28534 6808 28540 6860
rect 28592 6848 28598 6860
rect 28721 6851 28779 6857
rect 28721 6848 28733 6851
rect 28592 6820 28733 6848
rect 28592 6808 28598 6820
rect 28721 6817 28733 6820
rect 28767 6817 28779 6851
rect 28721 6811 28779 6817
rect 28905 6851 28963 6857
rect 28905 6817 28917 6851
rect 28951 6848 28963 6851
rect 29086 6848 29092 6860
rect 28951 6820 29092 6848
rect 28951 6817 28963 6820
rect 28905 6811 28963 6817
rect 29086 6808 29092 6820
rect 29144 6808 29150 6860
rect 29546 6808 29552 6860
rect 29604 6808 29610 6860
rect 29733 6851 29791 6857
rect 29733 6817 29745 6851
rect 29779 6848 29791 6851
rect 31389 6851 31447 6857
rect 31389 6848 31401 6851
rect 29779 6820 31401 6848
rect 29779 6817 29791 6820
rect 29733 6811 29791 6817
rect 31389 6817 31401 6820
rect 31435 6817 31447 6851
rect 31389 6811 31447 6817
rect 31754 6808 31760 6860
rect 31812 6848 31818 6860
rect 31941 6851 31999 6857
rect 31941 6848 31953 6851
rect 31812 6820 31953 6848
rect 31812 6808 31818 6820
rect 31941 6817 31953 6820
rect 31987 6817 31999 6851
rect 31941 6811 31999 6817
rect 32030 6808 32036 6860
rect 32088 6848 32094 6860
rect 32490 6848 32496 6860
rect 32088 6820 32496 6848
rect 32088 6808 32094 6820
rect 32490 6808 32496 6820
rect 32548 6808 32554 6860
rect 33134 6808 33140 6860
rect 33192 6848 33198 6860
rect 33229 6851 33287 6857
rect 33229 6848 33241 6851
rect 33192 6820 33241 6848
rect 33192 6808 33198 6820
rect 33229 6817 33241 6820
rect 33275 6817 33287 6851
rect 33229 6811 33287 6817
rect 33965 6851 34023 6857
rect 33965 6817 33977 6851
rect 34011 6848 34023 6851
rect 36354 6848 36360 6860
rect 34011 6820 36360 6848
rect 34011 6817 34023 6820
rect 33965 6811 34023 6817
rect 36354 6808 36360 6820
rect 36412 6808 36418 6860
rect 36538 6808 36544 6860
rect 36596 6808 36602 6860
rect 37277 6851 37335 6857
rect 37277 6817 37289 6851
rect 37323 6848 37335 6851
rect 37366 6848 37372 6860
rect 37323 6820 37372 6848
rect 37323 6817 37335 6820
rect 37277 6811 37335 6817
rect 37366 6808 37372 6820
rect 37424 6808 37430 6860
rect 37461 6851 37519 6857
rect 37461 6817 37473 6851
rect 37507 6848 37519 6851
rect 37826 6848 37832 6860
rect 37507 6820 37832 6848
rect 37507 6817 37519 6820
rect 37461 6811 37519 6817
rect 37826 6808 37832 6820
rect 37884 6808 37890 6860
rect 39574 6848 39580 6860
rect 39040 6820 39580 6848
rect 39040 6792 39068 6820
rect 39574 6808 39580 6820
rect 39632 6808 39638 6860
rect 39666 6808 39672 6860
rect 39724 6848 39730 6860
rect 42245 6851 42303 6857
rect 42245 6848 42257 6851
rect 39724 6820 42257 6848
rect 39724 6808 39730 6820
rect 42245 6817 42257 6820
rect 42291 6817 42303 6851
rect 42245 6811 42303 6817
rect 25961 6783 26019 6789
rect 25961 6749 25973 6783
rect 26007 6749 26019 6783
rect 25961 6743 26019 6749
rect 31297 6783 31355 6789
rect 31297 6749 31309 6783
rect 31343 6780 31355 6783
rect 31343 6752 31754 6780
rect 31343 6749 31355 6752
rect 31297 6743 31355 6749
rect 22495 6684 22600 6712
rect 22495 6681 22507 6684
rect 22449 6675 22507 6681
rect 22646 6672 22652 6724
rect 22704 6672 22710 6724
rect 24213 6715 24271 6721
rect 24213 6681 24225 6715
rect 24259 6712 24271 6715
rect 24762 6712 24768 6724
rect 24259 6684 24768 6712
rect 24259 6681 24271 6684
rect 24213 6675 24271 6681
rect 24762 6672 24768 6684
rect 24820 6672 24826 6724
rect 25133 6715 25191 6721
rect 25133 6681 25145 6715
rect 25179 6712 25191 6715
rect 30926 6712 30932 6724
rect 25179 6684 27384 6712
rect 28198 6684 30932 6712
rect 25179 6681 25191 6684
rect 25133 6675 25191 6681
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 10318 6644 10324 6656
rect 10091 6616 10324 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 11790 6604 11796 6656
rect 11848 6604 11854 6656
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 12621 6647 12679 6653
rect 12621 6644 12633 6647
rect 12492 6616 12633 6644
rect 12492 6604 12498 6616
rect 12621 6613 12633 6616
rect 12667 6613 12679 6647
rect 12621 6607 12679 6613
rect 13446 6604 13452 6656
rect 13504 6604 13510 6656
rect 14182 6604 14188 6656
rect 14240 6604 14246 6656
rect 14642 6604 14648 6656
rect 14700 6644 14706 6656
rect 15105 6647 15163 6653
rect 15105 6644 15117 6647
rect 14700 6616 15117 6644
rect 14700 6604 14706 6616
rect 15105 6613 15117 6616
rect 15151 6613 15163 6647
rect 15105 6607 15163 6613
rect 15289 6647 15347 6653
rect 15289 6613 15301 6647
rect 15335 6644 15347 6647
rect 15378 6644 15384 6656
rect 15335 6616 15384 6644
rect 15335 6613 15347 6616
rect 15289 6607 15347 6613
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 18141 6647 18199 6653
rect 18141 6644 18153 6647
rect 18104 6616 18153 6644
rect 18104 6604 18110 6616
rect 18141 6613 18153 6616
rect 18187 6613 18199 6647
rect 18141 6607 18199 6613
rect 21542 6604 21548 6656
rect 21600 6644 21606 6656
rect 22002 6644 22008 6656
rect 21600 6616 22008 6644
rect 21600 6604 21606 6616
rect 22002 6604 22008 6616
rect 22060 6604 22066 6656
rect 22278 6604 22284 6656
rect 22336 6604 22342 6656
rect 22554 6604 22560 6656
rect 22612 6644 22618 6656
rect 22833 6647 22891 6653
rect 22833 6644 22845 6647
rect 22612 6616 22845 6644
rect 22612 6604 22618 6616
rect 22833 6613 22845 6616
rect 22879 6613 22891 6647
rect 22833 6607 22891 6613
rect 25593 6647 25651 6653
rect 25593 6613 25605 6647
rect 25639 6644 25651 6647
rect 26602 6644 26608 6656
rect 25639 6616 26608 6644
rect 25639 6613 25651 6616
rect 25593 6607 25651 6613
rect 26602 6604 26608 6616
rect 26660 6604 26666 6656
rect 27356 6644 27384 6684
rect 30926 6672 30932 6684
rect 30984 6712 30990 6724
rect 30984 6684 31340 6712
rect 30984 6672 30990 6684
rect 31312 6656 31340 6684
rect 29362 6644 29368 6656
rect 27356 6616 29368 6644
rect 29362 6604 29368 6616
rect 29420 6604 29426 6656
rect 29546 6604 29552 6656
rect 29604 6644 29610 6656
rect 30374 6644 30380 6656
rect 29604 6616 30380 6644
rect 29604 6604 29610 6616
rect 30374 6604 30380 6616
rect 30432 6604 30438 6656
rect 30650 6604 30656 6656
rect 30708 6604 30714 6656
rect 31294 6604 31300 6656
rect 31352 6604 31358 6656
rect 31726 6644 31754 6752
rect 32582 6740 32588 6792
rect 32640 6740 32646 6792
rect 33318 6740 33324 6792
rect 33376 6740 33382 6792
rect 34238 6740 34244 6792
rect 34296 6780 34302 6792
rect 34609 6783 34667 6789
rect 34609 6780 34621 6783
rect 34296 6752 34621 6780
rect 34296 6740 34302 6752
rect 34609 6749 34621 6752
rect 34655 6780 34667 6783
rect 34882 6780 34888 6792
rect 34655 6752 34888 6780
rect 34655 6749 34667 6752
rect 34609 6743 34667 6749
rect 34882 6740 34888 6752
rect 34940 6780 34946 6792
rect 35250 6780 35256 6792
rect 34940 6752 35256 6780
rect 34940 6740 34946 6752
rect 35250 6740 35256 6752
rect 35308 6740 35314 6792
rect 35342 6740 35348 6792
rect 35400 6740 35406 6792
rect 35618 6740 35624 6792
rect 35676 6780 35682 6792
rect 35805 6783 35863 6789
rect 35805 6780 35817 6783
rect 35676 6752 35817 6780
rect 35676 6740 35682 6752
rect 35805 6749 35817 6752
rect 35851 6749 35863 6783
rect 35805 6743 35863 6749
rect 36725 6783 36783 6789
rect 36725 6749 36737 6783
rect 36771 6749 36783 6783
rect 39022 6780 39028 6792
rect 38870 6752 39028 6780
rect 36725 6743 36783 6749
rect 32030 6672 32036 6724
rect 32088 6712 32094 6724
rect 34057 6715 34115 6721
rect 34057 6712 34069 6715
rect 32088 6684 34069 6712
rect 32088 6672 32094 6684
rect 34057 6681 34069 6684
rect 34103 6681 34115 6715
rect 34057 6675 34115 6681
rect 35526 6672 35532 6724
rect 35584 6712 35590 6724
rect 35897 6715 35955 6721
rect 35897 6712 35909 6715
rect 35584 6684 35909 6712
rect 35584 6672 35590 6684
rect 35897 6681 35909 6684
rect 35943 6681 35955 6715
rect 35897 6675 35955 6681
rect 33226 6644 33232 6656
rect 31726 6616 33232 6644
rect 33226 6604 33232 6616
rect 33284 6604 33290 6656
rect 34790 6604 34796 6656
rect 34848 6604 34854 6656
rect 35066 6604 35072 6656
rect 35124 6644 35130 6656
rect 35713 6647 35771 6653
rect 35713 6644 35725 6647
rect 35124 6616 35725 6644
rect 35124 6604 35130 6616
rect 35713 6613 35725 6616
rect 35759 6613 35771 6647
rect 36740 6644 36768 6743
rect 39022 6740 39028 6752
rect 39080 6740 39086 6792
rect 40129 6783 40187 6789
rect 40129 6780 40141 6783
rect 39500 6752 40141 6780
rect 39500 6724 39528 6752
rect 40129 6749 40141 6752
rect 40175 6749 40187 6783
rect 40129 6743 40187 6749
rect 40218 6740 40224 6792
rect 40276 6780 40282 6792
rect 40773 6783 40831 6789
rect 40773 6780 40785 6783
rect 40276 6752 40785 6780
rect 40276 6740 40282 6752
rect 40773 6749 40785 6752
rect 40819 6749 40831 6783
rect 42061 6783 42119 6789
rect 42061 6780 42073 6783
rect 40773 6743 40831 6749
rect 41386 6752 42073 6780
rect 39482 6672 39488 6724
rect 39540 6672 39546 6724
rect 40402 6672 40408 6724
rect 40460 6712 40466 6724
rect 41386 6712 41414 6752
rect 42061 6749 42073 6752
rect 42107 6749 42119 6783
rect 42061 6743 42119 6749
rect 40460 6684 41414 6712
rect 40460 6672 40466 6684
rect 39022 6644 39028 6656
rect 36740 6616 39028 6644
rect 35713 6607 35771 6613
rect 39022 6604 39028 6616
rect 39080 6604 39086 6656
rect 39298 6604 39304 6656
rect 39356 6644 39362 6656
rect 39577 6647 39635 6653
rect 39577 6644 39589 6647
rect 39356 6616 39589 6644
rect 39356 6604 39362 6616
rect 39577 6613 39589 6616
rect 39623 6613 39635 6647
rect 39577 6607 39635 6613
rect 41414 6604 41420 6656
rect 41472 6604 41478 6656
rect 41506 6604 41512 6656
rect 41564 6604 41570 6656
rect 42889 6647 42947 6653
rect 42889 6613 42901 6647
rect 42935 6644 42947 6647
rect 46842 6644 46848 6656
rect 42935 6616 46848 6644
rect 42935 6613 42947 6616
rect 42889 6607 42947 6613
rect 46842 6604 46848 6616
rect 46900 6604 46906 6656
rect 2024 6554 77924 6576
rect 2024 6502 5794 6554
rect 5846 6502 5858 6554
rect 5910 6502 5922 6554
rect 5974 6502 5986 6554
rect 6038 6502 6050 6554
rect 6102 6502 36514 6554
rect 36566 6502 36578 6554
rect 36630 6502 36642 6554
rect 36694 6502 36706 6554
rect 36758 6502 36770 6554
rect 36822 6502 67234 6554
rect 67286 6502 67298 6554
rect 67350 6502 67362 6554
rect 67414 6502 67426 6554
rect 67478 6502 67490 6554
rect 67542 6502 77924 6554
rect 2024 6480 77924 6502
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 10704 6412 10885 6440
rect 8754 6332 8760 6384
rect 8812 6372 8818 6384
rect 10704 6372 10732 6412
rect 10873 6409 10885 6412
rect 10919 6409 10931 6443
rect 10873 6403 10931 6409
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 13446 6440 13452 6452
rect 11112 6412 13452 6440
rect 11112 6400 11118 6412
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 13725 6443 13783 6449
rect 13725 6409 13737 6443
rect 13771 6440 13783 6443
rect 16390 6440 16396 6452
rect 13771 6412 16396 6440
rect 13771 6409 13783 6412
rect 13725 6403 13783 6409
rect 16390 6400 16396 6412
rect 16448 6400 16454 6452
rect 17405 6443 17463 6449
rect 17405 6409 17417 6443
rect 17451 6440 17463 6443
rect 17678 6440 17684 6452
rect 17451 6412 17684 6440
rect 17451 6409 17463 6412
rect 17405 6403 17463 6409
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 18506 6400 18512 6452
rect 18564 6440 18570 6452
rect 18782 6440 18788 6452
rect 18564 6412 18788 6440
rect 18564 6400 18570 6412
rect 18782 6400 18788 6412
rect 18840 6400 18846 6452
rect 19150 6400 19156 6452
rect 19208 6440 19214 6452
rect 21358 6440 21364 6452
rect 19208 6412 21364 6440
rect 19208 6400 19214 6412
rect 21358 6400 21364 6412
rect 21416 6400 21422 6452
rect 22002 6400 22008 6452
rect 22060 6440 22066 6452
rect 23201 6443 23259 6449
rect 22060 6412 23060 6440
rect 22060 6400 22066 6412
rect 8812 6344 10732 6372
rect 10781 6375 10839 6381
rect 8812 6332 8818 6344
rect 10781 6341 10793 6375
rect 10827 6372 10839 6375
rect 10962 6372 10968 6384
rect 10827 6344 10968 6372
rect 10827 6341 10839 6344
rect 10781 6335 10839 6341
rect 10962 6332 10968 6344
rect 11020 6332 11026 6384
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 12253 6375 12311 6381
rect 11480 6344 12204 6372
rect 11480 6332 11486 6344
rect 9766 6264 9772 6316
rect 9824 6264 9830 6316
rect 11517 6307 11575 6313
rect 9876 6276 11284 6304
rect 8570 6196 8576 6248
rect 8628 6236 8634 6248
rect 9585 6239 9643 6245
rect 9585 6236 9597 6239
rect 8628 6208 9597 6236
rect 8628 6196 8634 6208
rect 9585 6205 9597 6208
rect 9631 6205 9643 6239
rect 9585 6199 9643 6205
rect 5626 6128 5632 6180
rect 5684 6168 5690 6180
rect 9876 6168 9904 6276
rect 10229 6239 10287 6245
rect 10229 6205 10241 6239
rect 10275 6236 10287 6239
rect 11146 6236 11152 6248
rect 10275 6208 11152 6236
rect 10275 6205 10287 6208
rect 10229 6199 10287 6205
rect 11146 6196 11152 6208
rect 11204 6196 11210 6248
rect 11256 6236 11284 6276
rect 11517 6273 11529 6307
rect 11563 6304 11575 6307
rect 12066 6304 12072 6316
rect 11563 6276 12072 6304
rect 11563 6273 11575 6276
rect 11517 6267 11575 6273
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 12176 6304 12204 6344
rect 12253 6341 12265 6375
rect 12299 6372 12311 6375
rect 14090 6372 14096 6384
rect 12299 6344 14096 6372
rect 12299 6341 12311 6344
rect 12253 6335 12311 6341
rect 14090 6332 14096 6344
rect 14148 6332 14154 6384
rect 15654 6372 15660 6384
rect 14384 6344 15660 6372
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 12176 6276 12449 6304
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 12805 6307 12863 6313
rect 12805 6273 12817 6307
rect 12851 6273 12863 6307
rect 12805 6267 12863 6273
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6304 13231 6307
rect 14384 6304 14412 6344
rect 15654 6332 15660 6344
rect 15712 6332 15718 6384
rect 17586 6332 17592 6384
rect 17644 6372 17650 6384
rect 17862 6372 17868 6384
rect 17644 6344 17868 6372
rect 17644 6332 17650 6344
rect 17862 6332 17868 6344
rect 17920 6332 17926 6384
rect 19242 6332 19248 6384
rect 19300 6372 19306 6384
rect 19300 6344 20576 6372
rect 19300 6332 19306 6344
rect 13219 6276 14412 6304
rect 13219 6273 13231 6276
rect 13173 6267 13231 6273
rect 11609 6239 11667 6245
rect 11609 6236 11621 6239
rect 11256 6208 11621 6236
rect 11609 6205 11621 6208
rect 11655 6205 11667 6239
rect 11609 6199 11667 6205
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 12820 6236 12848 6267
rect 14642 6264 14648 6316
rect 14700 6264 14706 6316
rect 14734 6264 14740 6316
rect 14792 6304 14798 6316
rect 15470 6304 15476 6316
rect 14792 6276 15476 6304
rect 14792 6264 14798 6276
rect 15470 6264 15476 6276
rect 15528 6264 15534 6316
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16206 6304 16212 6316
rect 15979 6276 16212 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 16666 6264 16672 6316
rect 16724 6264 16730 6316
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6304 16911 6307
rect 19610 6304 19616 6316
rect 16899 6276 19616 6304
rect 16899 6273 16911 6276
rect 16853 6267 16911 6273
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 19797 6307 19855 6313
rect 19797 6273 19809 6307
rect 19843 6304 19855 6307
rect 20070 6304 20076 6316
rect 19843 6276 20076 6304
rect 19843 6273 19855 6276
rect 19797 6267 19855 6273
rect 20070 6264 20076 6276
rect 20128 6264 20134 6316
rect 20548 6304 20576 6344
rect 21082 6332 21088 6384
rect 21140 6372 21146 6384
rect 21269 6375 21327 6381
rect 21269 6372 21281 6375
rect 21140 6344 21281 6372
rect 21140 6332 21146 6344
rect 21269 6341 21281 6344
rect 21315 6341 21327 6375
rect 21269 6335 21327 6341
rect 22189 6375 22247 6381
rect 22189 6341 22201 6375
rect 22235 6341 22247 6375
rect 22189 6335 22247 6341
rect 21358 6304 21364 6316
rect 20548 6276 21364 6304
rect 21358 6264 21364 6276
rect 21416 6304 21422 6316
rect 21729 6307 21787 6313
rect 21729 6304 21741 6307
rect 21416 6276 21741 6304
rect 21416 6264 21422 6276
rect 21729 6273 21741 6276
rect 21775 6273 21787 6307
rect 22204 6304 22232 6335
rect 22370 6332 22376 6384
rect 22428 6381 22434 6384
rect 23032 6381 23060 6412
rect 23201 6409 23213 6443
rect 23247 6440 23259 6443
rect 23290 6440 23296 6452
rect 23247 6412 23296 6440
rect 23247 6409 23259 6412
rect 23201 6403 23259 6409
rect 23290 6400 23296 6412
rect 23348 6400 23354 6452
rect 23385 6443 23443 6449
rect 23385 6409 23397 6443
rect 23431 6440 23443 6443
rect 24026 6440 24032 6452
rect 23431 6412 24032 6440
rect 23431 6409 23443 6412
rect 23385 6403 23443 6409
rect 24026 6400 24032 6412
rect 24084 6400 24090 6452
rect 24394 6400 24400 6452
rect 24452 6400 24458 6452
rect 26694 6400 26700 6452
rect 26752 6440 26758 6452
rect 26881 6443 26939 6449
rect 26881 6440 26893 6443
rect 26752 6412 26893 6440
rect 26752 6400 26758 6412
rect 26881 6409 26893 6412
rect 26927 6409 26939 6443
rect 26881 6403 26939 6409
rect 27249 6443 27307 6449
rect 27249 6409 27261 6443
rect 27295 6440 27307 6443
rect 27706 6440 27712 6452
rect 27295 6412 27712 6440
rect 27295 6409 27307 6412
rect 27249 6403 27307 6409
rect 27706 6400 27712 6412
rect 27764 6400 27770 6452
rect 30098 6440 30104 6452
rect 30024 6412 30104 6440
rect 22428 6375 22447 6381
rect 22435 6341 22447 6375
rect 22428 6335 22447 6341
rect 23017 6375 23075 6381
rect 23017 6341 23029 6375
rect 23063 6341 23075 6375
rect 26605 6375 26663 6381
rect 23017 6335 23075 6341
rect 23124 6344 23428 6372
rect 22428 6332 22434 6335
rect 23124 6304 23152 6344
rect 23400 6316 23428 6344
rect 26605 6341 26617 6375
rect 26651 6372 26663 6375
rect 26786 6372 26792 6384
rect 26651 6344 26792 6372
rect 26651 6341 26663 6344
rect 23584 6316 23796 6338
rect 26605 6335 26663 6341
rect 26786 6332 26792 6344
rect 26844 6332 26850 6384
rect 27341 6375 27399 6381
rect 27341 6341 27353 6375
rect 27387 6372 27399 6375
rect 27522 6372 27528 6384
rect 27387 6344 27528 6372
rect 27387 6341 27399 6344
rect 27341 6335 27399 6341
rect 27522 6332 27528 6344
rect 27580 6332 27586 6384
rect 27614 6332 27620 6384
rect 27672 6372 27678 6384
rect 29454 6372 29460 6384
rect 27672 6344 29460 6372
rect 27672 6332 27678 6344
rect 29454 6332 29460 6344
rect 29512 6332 29518 6384
rect 29730 6332 29736 6384
rect 29788 6372 29794 6384
rect 29788 6344 29868 6372
rect 29788 6332 29794 6344
rect 22204 6276 23152 6304
rect 21729 6267 21787 6273
rect 23290 6264 23296 6316
rect 23348 6264 23354 6316
rect 23382 6264 23388 6316
rect 23440 6264 23446 6316
rect 23584 6310 23756 6316
rect 13262 6236 13268 6248
rect 11848 6208 13268 6236
rect 11848 6196 11854 6208
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 13817 6239 13875 6245
rect 13817 6205 13829 6239
rect 13863 6236 13875 6239
rect 13906 6236 13912 6248
rect 13863 6208 13912 6236
rect 13863 6205 13875 6208
rect 13817 6199 13875 6205
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 14366 6196 14372 6248
rect 14424 6196 14430 6248
rect 15197 6239 15255 6245
rect 15197 6205 15209 6239
rect 15243 6236 15255 6239
rect 15562 6236 15568 6248
rect 15243 6208 15568 6236
rect 15243 6205 15255 6208
rect 15197 6199 15255 6205
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 17402 6196 17408 6248
rect 17460 6236 17466 6248
rect 17681 6239 17739 6245
rect 17681 6236 17693 6239
rect 17460 6208 17693 6236
rect 17460 6196 17466 6208
rect 17681 6205 17693 6208
rect 17727 6205 17739 6239
rect 17681 6199 17739 6205
rect 17862 6196 17868 6248
rect 17920 6236 17926 6248
rect 18233 6239 18291 6245
rect 18233 6236 18245 6239
rect 17920 6208 18245 6236
rect 17920 6196 17926 6208
rect 18233 6205 18245 6208
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 19061 6239 19119 6245
rect 19061 6205 19073 6239
rect 19107 6236 19119 6239
rect 19426 6236 19432 6248
rect 19107 6208 19432 6236
rect 19107 6205 19119 6208
rect 19061 6199 19119 6205
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 19886 6196 19892 6248
rect 19944 6196 19950 6248
rect 19978 6196 19984 6248
rect 20036 6236 20042 6248
rect 20625 6239 20683 6245
rect 20625 6236 20637 6239
rect 20036 6208 20637 6236
rect 20036 6196 20042 6208
rect 20625 6205 20637 6208
rect 20671 6205 20683 6239
rect 20625 6199 20683 6205
rect 21634 6196 21640 6248
rect 21692 6236 21698 6248
rect 21821 6239 21879 6245
rect 21821 6236 21833 6239
rect 21692 6208 21833 6236
rect 21692 6196 21698 6208
rect 21821 6205 21833 6208
rect 21867 6205 21879 6239
rect 21821 6199 21879 6205
rect 21913 6239 21971 6245
rect 21913 6205 21925 6239
rect 21959 6205 21971 6239
rect 21913 6199 21971 6205
rect 5684 6140 9904 6168
rect 9953 6171 10011 6177
rect 5684 6128 5690 6140
rect 9953 6137 9965 6171
rect 9999 6168 10011 6171
rect 9999 6140 18920 6168
rect 9999 6137 10011 6140
rect 9953 6131 10011 6137
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 9033 6103 9091 6109
rect 9033 6100 9045 6103
rect 6972 6072 9045 6100
rect 6972 6060 6978 6072
rect 9033 6069 9045 6072
rect 9079 6069 9091 6103
rect 9033 6063 9091 6069
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 13630 6100 13636 6112
rect 9640 6072 13636 6100
rect 9640 6060 9646 6072
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 14090 6060 14096 6112
rect 14148 6100 14154 6112
rect 15289 6103 15347 6109
rect 15289 6100 15301 6103
rect 14148 6072 15301 6100
rect 14148 6060 14154 6072
rect 15289 6069 15301 6072
rect 15335 6069 15347 6103
rect 15289 6063 15347 6069
rect 16022 6060 16028 6112
rect 16080 6060 16086 6112
rect 16574 6060 16580 6112
rect 16632 6100 16638 6112
rect 18417 6103 18475 6109
rect 18417 6100 18429 6103
rect 16632 6072 18429 6100
rect 16632 6060 16638 6072
rect 18417 6069 18429 6072
rect 18463 6069 18475 6103
rect 18892 6100 18920 6140
rect 19150 6128 19156 6180
rect 19208 6128 19214 6180
rect 20346 6128 20352 6180
rect 20404 6168 20410 6180
rect 20533 6171 20591 6177
rect 20533 6168 20545 6171
rect 20404 6140 20545 6168
rect 20404 6128 20410 6140
rect 20533 6137 20545 6140
rect 20579 6137 20591 6171
rect 20533 6131 20591 6137
rect 21726 6128 21732 6180
rect 21784 6168 21790 6180
rect 21928 6168 21956 6199
rect 22738 6196 22744 6248
rect 22796 6236 22802 6248
rect 23308 6236 23336 6264
rect 23584 6236 23612 6310
rect 23750 6264 23756 6310
rect 23808 6264 23814 6316
rect 23842 6264 23848 6316
rect 23900 6264 23906 6316
rect 25038 6264 25044 6316
rect 25096 6304 25102 6316
rect 26053 6307 26111 6313
rect 25096 6276 25452 6304
rect 25096 6264 25102 6276
rect 22796 6208 23336 6236
rect 23492 6208 23612 6236
rect 22796 6196 22802 6208
rect 22557 6171 22615 6177
rect 21784 6140 22508 6168
rect 21784 6128 21790 6140
rect 19242 6100 19248 6112
rect 18892 6072 19248 6100
rect 18417 6063 18475 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 21361 6103 21419 6109
rect 21361 6069 21373 6103
rect 21407 6100 21419 6103
rect 21818 6100 21824 6112
rect 21407 6072 21824 6100
rect 21407 6069 21419 6072
rect 21361 6063 21419 6069
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 22186 6060 22192 6112
rect 22244 6100 22250 6112
rect 22333 6103 22391 6109
rect 22333 6100 22345 6103
rect 22244 6072 22345 6100
rect 22244 6060 22250 6072
rect 22333 6069 22345 6072
rect 22379 6069 22391 6103
rect 22480 6100 22508 6140
rect 22557 6137 22569 6171
rect 22603 6168 22615 6171
rect 23492 6168 23520 6208
rect 23934 6196 23940 6248
rect 23992 6236 23998 6248
rect 24489 6239 24547 6245
rect 24489 6236 24501 6239
rect 23992 6208 24501 6236
rect 23992 6196 23998 6208
rect 24489 6205 24501 6208
rect 24535 6205 24547 6239
rect 24489 6199 24547 6205
rect 25314 6196 25320 6248
rect 25372 6196 25378 6248
rect 25424 6236 25452 6276
rect 26053 6273 26065 6307
rect 26099 6304 26111 6307
rect 26142 6304 26148 6316
rect 26099 6276 26148 6304
rect 26099 6273 26111 6276
rect 26053 6267 26111 6273
rect 26142 6264 26148 6276
rect 26200 6264 26206 6316
rect 27893 6307 27951 6313
rect 27893 6273 27905 6307
rect 27939 6304 27951 6307
rect 28994 6304 29000 6316
rect 27939 6276 29000 6304
rect 27939 6273 27951 6276
rect 27893 6267 27951 6273
rect 28994 6264 29000 6276
rect 29052 6264 29058 6316
rect 29840 6313 29868 6344
rect 30024 6313 30052 6412
rect 30098 6400 30104 6412
rect 30156 6400 30162 6452
rect 30374 6440 30380 6452
rect 30208 6412 30380 6440
rect 30208 6372 30236 6412
rect 30374 6400 30380 6412
rect 30432 6400 30438 6452
rect 31294 6400 31300 6452
rect 31352 6440 31358 6452
rect 35621 6443 35679 6449
rect 31352 6412 32720 6440
rect 31352 6400 31358 6412
rect 30116 6344 30236 6372
rect 30116 6313 30144 6344
rect 30282 6332 30288 6384
rect 30340 6372 30346 6384
rect 30340 6344 31432 6372
rect 30340 6332 30346 6344
rect 29825 6307 29883 6313
rect 29825 6273 29837 6307
rect 29871 6273 29883 6307
rect 29825 6267 29883 6273
rect 30009 6307 30067 6313
rect 30009 6273 30021 6307
rect 30055 6273 30067 6307
rect 30009 6267 30067 6273
rect 30101 6307 30159 6313
rect 30101 6273 30113 6307
rect 30147 6273 30159 6307
rect 30101 6267 30159 6273
rect 30208 6276 30696 6304
rect 26786 6236 26792 6248
rect 25424 6208 26792 6236
rect 26786 6196 26792 6208
rect 26844 6236 26850 6248
rect 27433 6239 27491 6245
rect 27433 6236 27445 6239
rect 26844 6208 27445 6236
rect 26844 6196 26850 6208
rect 27433 6205 27445 6208
rect 27479 6236 27491 6239
rect 28902 6236 28908 6248
rect 27479 6208 28908 6236
rect 27479 6205 27491 6208
rect 27433 6199 27491 6205
rect 28902 6196 28908 6208
rect 28960 6196 28966 6248
rect 29638 6196 29644 6248
rect 29696 6196 29702 6248
rect 29914 6196 29920 6248
rect 29972 6196 29978 6248
rect 22603 6140 23520 6168
rect 23569 6171 23627 6177
rect 22603 6137 22615 6140
rect 22557 6131 22615 6137
rect 23569 6137 23581 6171
rect 23615 6168 23627 6171
rect 29546 6168 29552 6180
rect 23615 6140 29552 6168
rect 23615 6137 23627 6140
rect 23569 6131 23627 6137
rect 29546 6128 29552 6140
rect 29604 6128 29610 6180
rect 25038 6100 25044 6112
rect 22480 6072 25044 6100
rect 22333 6063 22391 6069
rect 25038 6060 25044 6072
rect 25096 6060 25102 6112
rect 25130 6060 25136 6112
rect 25188 6060 25194 6112
rect 25869 6103 25927 6109
rect 25869 6069 25881 6103
rect 25915 6100 25927 6103
rect 28534 6100 28540 6112
rect 25915 6072 28540 6100
rect 25915 6069 25927 6072
rect 25869 6063 25927 6069
rect 28534 6060 28540 6072
rect 28592 6060 28598 6112
rect 29730 6060 29736 6112
rect 29788 6100 29794 6112
rect 30208 6100 30236 6276
rect 30285 6239 30343 6245
rect 30285 6205 30297 6239
rect 30331 6236 30343 6239
rect 30668 6236 30696 6276
rect 30926 6264 30932 6316
rect 30984 6264 30990 6316
rect 31404 6304 31432 6344
rect 31754 6332 31760 6384
rect 31812 6372 31818 6384
rect 32692 6372 32720 6412
rect 35621 6409 35633 6443
rect 35667 6440 35679 6443
rect 38838 6440 38844 6452
rect 35667 6412 38844 6440
rect 35667 6409 35679 6412
rect 35621 6403 35679 6409
rect 38838 6400 38844 6412
rect 38896 6400 38902 6452
rect 31812 6344 31984 6372
rect 32692 6344 33810 6372
rect 31812 6332 31818 6344
rect 31849 6307 31907 6313
rect 31849 6304 31861 6307
rect 31404 6276 31861 6304
rect 31849 6273 31861 6276
rect 31895 6273 31907 6307
rect 31956 6304 31984 6344
rect 34882 6332 34888 6384
rect 34940 6372 34946 6384
rect 35069 6375 35127 6381
rect 35069 6372 35081 6375
rect 34940 6344 35081 6372
rect 34940 6332 34946 6344
rect 35069 6341 35081 6344
rect 35115 6341 35127 6375
rect 35069 6335 35127 6341
rect 38013 6375 38071 6381
rect 38013 6341 38025 6375
rect 38059 6372 38071 6375
rect 38473 6375 38531 6381
rect 38473 6372 38485 6375
rect 38059 6344 38485 6372
rect 38059 6341 38071 6344
rect 38013 6335 38071 6341
rect 38473 6341 38485 6344
rect 38519 6341 38531 6375
rect 38473 6335 38531 6341
rect 40218 6332 40224 6384
rect 40276 6332 40282 6384
rect 43346 6372 43352 6384
rect 42996 6344 43352 6372
rect 32585 6307 32643 6313
rect 31956 6294 32536 6304
rect 32585 6294 32597 6307
rect 31956 6276 32597 6294
rect 31849 6267 31907 6273
rect 32508 6273 32597 6276
rect 32631 6273 32643 6307
rect 32508 6267 32643 6273
rect 32508 6266 32628 6267
rect 35158 6264 35164 6316
rect 35216 6264 35222 6316
rect 35250 6264 35256 6316
rect 35308 6264 35314 6316
rect 35437 6307 35495 6313
rect 35437 6273 35449 6307
rect 35483 6273 35495 6307
rect 35437 6267 35495 6273
rect 31113 6239 31171 6245
rect 31113 6236 31125 6239
rect 30331 6208 30604 6236
rect 30668 6208 31125 6236
rect 30331 6205 30343 6208
rect 30285 6199 30343 6205
rect 29788 6072 30236 6100
rect 29788 6060 29794 6072
rect 30374 6060 30380 6112
rect 30432 6060 30438 6112
rect 30576 6100 30604 6208
rect 31113 6205 31125 6208
rect 31159 6205 31171 6239
rect 31113 6199 31171 6205
rect 31754 6196 31760 6248
rect 31812 6196 31818 6248
rect 32122 6196 32128 6248
rect 32180 6236 32186 6248
rect 32677 6239 32735 6245
rect 32677 6236 32689 6239
rect 32180 6208 32689 6236
rect 32180 6196 32186 6208
rect 32677 6205 32689 6208
rect 32723 6205 32735 6239
rect 32677 6199 32735 6205
rect 32950 6196 32956 6248
rect 33008 6236 33014 6248
rect 33045 6239 33103 6245
rect 33045 6236 33057 6239
rect 33008 6208 33057 6236
rect 33008 6196 33014 6208
rect 33045 6205 33057 6208
rect 33091 6205 33103 6239
rect 33045 6199 33103 6205
rect 33321 6239 33379 6245
rect 33321 6205 33333 6239
rect 33367 6236 33379 6239
rect 33410 6236 33416 6248
rect 33367 6208 33416 6236
rect 33367 6205 33379 6208
rect 33321 6199 33379 6205
rect 33410 6196 33416 6208
rect 33468 6196 33474 6248
rect 34882 6196 34888 6248
rect 34940 6236 34946 6248
rect 35452 6236 35480 6267
rect 35710 6264 35716 6316
rect 35768 6304 35774 6316
rect 36265 6307 36323 6313
rect 36265 6304 36277 6307
rect 35768 6276 36277 6304
rect 35768 6264 35774 6276
rect 36265 6273 36277 6276
rect 36311 6273 36323 6307
rect 36265 6267 36323 6273
rect 36998 6264 37004 6316
rect 37056 6304 37062 6316
rect 37369 6307 37427 6313
rect 37369 6304 37381 6307
rect 37056 6276 37381 6304
rect 37056 6264 37062 6276
rect 37369 6273 37381 6276
rect 37415 6273 37427 6307
rect 37369 6267 37427 6273
rect 39574 6264 39580 6316
rect 39632 6264 39638 6316
rect 41414 6264 41420 6316
rect 41472 6304 41478 6316
rect 41785 6307 41843 6313
rect 41785 6304 41797 6307
rect 41472 6276 41797 6304
rect 41472 6264 41478 6276
rect 41785 6273 41797 6276
rect 41831 6273 41843 6307
rect 41785 6267 41843 6273
rect 42702 6264 42708 6316
rect 42760 6264 42766 6316
rect 42794 6264 42800 6316
rect 42852 6264 42858 6316
rect 42996 6313 43024 6344
rect 43346 6332 43352 6344
rect 43404 6332 43410 6384
rect 42981 6307 43039 6313
rect 42981 6273 42993 6307
rect 43027 6273 43039 6307
rect 42981 6267 43039 6273
rect 43254 6264 43260 6316
rect 43312 6304 43318 6316
rect 44085 6307 44143 6313
rect 44085 6304 44097 6307
rect 43312 6276 44097 6304
rect 43312 6264 43318 6276
rect 44085 6273 44097 6276
rect 44131 6273 44143 6307
rect 44085 6267 44143 6273
rect 34940 6208 35480 6236
rect 34940 6196 34946 6208
rect 35618 6196 35624 6248
rect 35676 6236 35682 6248
rect 37277 6239 37335 6245
rect 35676 6208 37228 6236
rect 35676 6196 35682 6208
rect 32493 6171 32551 6177
rect 32493 6137 32505 6171
rect 32539 6168 32551 6171
rect 32582 6168 32588 6180
rect 32539 6140 32588 6168
rect 32539 6137 32551 6140
rect 32493 6131 32551 6137
rect 32582 6128 32588 6140
rect 32640 6128 32646 6180
rect 34330 6128 34336 6180
rect 34388 6168 34394 6180
rect 35713 6171 35771 6177
rect 35713 6168 35725 6171
rect 34388 6140 35725 6168
rect 34388 6128 34394 6140
rect 35713 6137 35725 6140
rect 35759 6137 35771 6171
rect 35713 6131 35771 6137
rect 33134 6100 33140 6112
rect 30576 6072 33140 6100
rect 33134 6060 33140 6072
rect 33192 6060 33198 6112
rect 35250 6060 35256 6112
rect 35308 6100 35314 6112
rect 35618 6100 35624 6112
rect 35308 6072 35624 6100
rect 35308 6060 35314 6072
rect 35618 6060 35624 6072
rect 35676 6100 35682 6112
rect 36446 6100 36452 6112
rect 35676 6072 36452 6100
rect 35676 6060 35682 6072
rect 36446 6060 36452 6072
rect 36504 6060 36510 6112
rect 36633 6103 36691 6109
rect 36633 6069 36645 6103
rect 36679 6100 36691 6103
rect 36906 6100 36912 6112
rect 36679 6072 36912 6100
rect 36679 6069 36691 6072
rect 36633 6063 36691 6069
rect 36906 6060 36912 6072
rect 36964 6060 36970 6112
rect 37200 6100 37228 6208
rect 37277 6205 37289 6239
rect 37323 6205 37335 6239
rect 37277 6199 37335 6205
rect 37292 6168 37320 6199
rect 37918 6196 37924 6248
rect 37976 6236 37982 6248
rect 38197 6239 38255 6245
rect 38197 6236 38209 6239
rect 37976 6208 38209 6236
rect 37976 6196 37982 6208
rect 38197 6205 38209 6208
rect 38243 6205 38255 6239
rect 38930 6236 38936 6248
rect 38197 6199 38255 6205
rect 38304 6208 38936 6236
rect 38304 6168 38332 6208
rect 38930 6196 38936 6208
rect 38988 6196 38994 6248
rect 40589 6239 40647 6245
rect 40589 6205 40601 6239
rect 40635 6236 40647 6239
rect 41233 6239 41291 6245
rect 41233 6236 41245 6239
rect 40635 6208 41245 6236
rect 40635 6205 40647 6208
rect 40589 6199 40647 6205
rect 41233 6205 41245 6208
rect 41279 6205 41291 6239
rect 41233 6199 41291 6205
rect 42613 6239 42671 6245
rect 42613 6205 42625 6239
rect 42659 6236 42671 6239
rect 43165 6239 43223 6245
rect 43165 6236 43177 6239
rect 42659 6208 43177 6236
rect 42659 6205 42671 6208
rect 42613 6199 42671 6205
rect 43165 6205 43177 6208
rect 43211 6205 43223 6239
rect 43165 6199 43223 6205
rect 43349 6239 43407 6245
rect 43349 6205 43361 6239
rect 43395 6205 43407 6239
rect 43349 6199 43407 6205
rect 37292 6140 38332 6168
rect 39482 6100 39488 6112
rect 37200 6072 39488 6100
rect 39482 6060 39488 6072
rect 39540 6060 39546 6112
rect 41138 6060 41144 6112
rect 41196 6060 41202 6112
rect 41966 6060 41972 6112
rect 42024 6060 42030 6112
rect 42610 6060 42616 6112
rect 42668 6100 42674 6112
rect 43364 6100 43392 6199
rect 43993 6171 44051 6177
rect 43993 6137 44005 6171
rect 44039 6168 44051 6171
rect 45462 6168 45468 6180
rect 44039 6140 45468 6168
rect 44039 6137 44051 6140
rect 43993 6131 44051 6137
rect 45462 6128 45468 6140
rect 45520 6128 45526 6180
rect 42668 6072 43392 6100
rect 44729 6103 44787 6109
rect 42668 6060 42674 6072
rect 44729 6069 44741 6103
rect 44775 6100 44787 6103
rect 48866 6100 48872 6112
rect 44775 6072 48872 6100
rect 44775 6069 44787 6072
rect 44729 6063 44787 6069
rect 48866 6060 48872 6072
rect 48924 6060 48930 6112
rect 2024 6010 77924 6032
rect 2024 5958 5134 6010
rect 5186 5958 5198 6010
rect 5250 5958 5262 6010
rect 5314 5958 5326 6010
rect 5378 5958 5390 6010
rect 5442 5958 35854 6010
rect 35906 5958 35918 6010
rect 35970 5958 35982 6010
rect 36034 5958 36046 6010
rect 36098 5958 36110 6010
rect 36162 5958 66574 6010
rect 66626 5958 66638 6010
rect 66690 5958 66702 6010
rect 66754 5958 66766 6010
rect 66818 5958 66830 6010
rect 66882 5958 77924 6010
rect 2024 5936 77924 5958
rect 8570 5856 8576 5908
rect 8628 5856 8634 5908
rect 12713 5899 12771 5905
rect 12713 5896 12725 5899
rect 11256 5868 12725 5896
rect 5718 5788 5724 5840
rect 5776 5828 5782 5840
rect 11054 5828 11060 5840
rect 5776 5800 11060 5828
rect 5776 5788 5782 5800
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 7800 5732 10548 5760
rect 7800 5720 7806 5732
rect 8018 5652 8024 5704
rect 8076 5652 8082 5704
rect 9030 5652 9036 5704
rect 9088 5652 9094 5704
rect 9582 5652 9588 5704
rect 9640 5692 9646 5704
rect 10336 5701 10364 5732
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 9640 5664 10149 5692
rect 9640 5652 9646 5664
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5661 10379 5695
rect 10321 5655 10379 5661
rect 10410 5652 10416 5704
rect 10468 5652 10474 5704
rect 10520 5692 10548 5732
rect 10594 5720 10600 5772
rect 10652 5720 10658 5772
rect 11256 5769 11284 5868
rect 12713 5865 12725 5868
rect 12759 5865 12771 5899
rect 12713 5859 12771 5865
rect 14829 5899 14887 5905
rect 14829 5865 14841 5899
rect 14875 5896 14887 5899
rect 17494 5896 17500 5908
rect 14875 5868 17500 5896
rect 14875 5865 14887 5868
rect 14829 5859 14887 5865
rect 17494 5856 17500 5868
rect 17552 5856 17558 5908
rect 18509 5899 18567 5905
rect 18509 5865 18521 5899
rect 18555 5896 18567 5899
rect 18555 5868 20116 5896
rect 18555 5865 18567 5868
rect 18509 5859 18567 5865
rect 15565 5831 15623 5837
rect 11808 5800 14688 5828
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5729 11299 5763
rect 11241 5723 11299 5729
rect 11808 5692 11836 5800
rect 11882 5720 11888 5772
rect 11940 5720 11946 5772
rect 14550 5760 14556 5772
rect 13372 5732 14556 5760
rect 10520 5664 11836 5692
rect 11974 5652 11980 5704
rect 12032 5652 12038 5704
rect 13262 5652 13268 5704
rect 13320 5652 13326 5704
rect 8570 5584 8576 5636
rect 8628 5624 8634 5636
rect 9600 5624 9628 5652
rect 8628 5596 9628 5624
rect 9677 5627 9735 5633
rect 8628 5584 8634 5596
rect 9677 5593 9689 5627
rect 9723 5624 9735 5627
rect 10226 5624 10232 5636
rect 9723 5596 10232 5624
rect 9723 5593 9735 5596
rect 9677 5587 9735 5593
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 11149 5627 11207 5633
rect 11149 5593 11161 5627
rect 11195 5624 11207 5627
rect 13372 5624 13400 5732
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 14660 5760 14688 5800
rect 15565 5797 15577 5831
rect 15611 5828 15623 5831
rect 16301 5831 16359 5837
rect 15611 5800 15700 5828
rect 15611 5797 15623 5800
rect 15565 5791 15623 5797
rect 14826 5760 14832 5772
rect 14660 5732 14832 5760
rect 14826 5720 14832 5732
rect 14884 5760 14890 5772
rect 15672 5769 15700 5800
rect 16301 5797 16313 5831
rect 16347 5828 16359 5831
rect 19518 5828 19524 5840
rect 16347 5800 19524 5828
rect 16347 5797 16359 5800
rect 16301 5791 16359 5797
rect 19518 5788 19524 5800
rect 19576 5788 19582 5840
rect 20088 5828 20116 5868
rect 20162 5856 20168 5908
rect 20220 5856 20226 5908
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20349 5899 20407 5905
rect 20349 5896 20361 5899
rect 20312 5868 20361 5896
rect 20312 5856 20318 5868
rect 20349 5865 20361 5868
rect 20395 5896 20407 5899
rect 20806 5896 20812 5908
rect 20395 5868 20812 5896
rect 20395 5865 20407 5868
rect 20349 5859 20407 5865
rect 20806 5856 20812 5868
rect 20864 5856 20870 5908
rect 21450 5856 21456 5908
rect 21508 5856 21514 5908
rect 22002 5856 22008 5908
rect 22060 5896 22066 5908
rect 23934 5896 23940 5908
rect 22060 5868 23940 5896
rect 22060 5856 22066 5868
rect 23934 5856 23940 5868
rect 23992 5856 23998 5908
rect 24302 5856 24308 5908
rect 24360 5896 24366 5908
rect 24397 5899 24455 5905
rect 24397 5896 24409 5899
rect 24360 5868 24409 5896
rect 24360 5856 24366 5868
rect 24397 5865 24409 5868
rect 24443 5865 24455 5899
rect 26326 5896 26332 5908
rect 24397 5859 24455 5865
rect 25056 5868 26332 5896
rect 20530 5828 20536 5840
rect 20088 5800 20536 5828
rect 20530 5788 20536 5800
rect 20588 5788 20594 5840
rect 20717 5831 20775 5837
rect 20717 5797 20729 5831
rect 20763 5828 20775 5831
rect 22278 5828 22284 5840
rect 20763 5800 22284 5828
rect 20763 5797 20775 5800
rect 20717 5791 20775 5797
rect 22278 5788 22284 5800
rect 22336 5828 22342 5840
rect 23750 5828 23756 5840
rect 22336 5800 23756 5828
rect 22336 5788 22342 5800
rect 23750 5788 23756 5800
rect 23808 5788 23814 5840
rect 24670 5828 24676 5840
rect 24504 5800 24676 5828
rect 15657 5763 15715 5769
rect 14884 5732 15240 5760
rect 14884 5720 14890 5732
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5692 14335 5695
rect 14642 5692 14648 5704
rect 14323 5664 14648 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 11195 5596 13400 5624
rect 11195 5593 11207 5596
rect 11149 5587 11207 5593
rect 13446 5584 13452 5636
rect 13504 5584 13510 5636
rect 14108 5624 14136 5655
rect 14642 5652 14648 5664
rect 14700 5652 14706 5704
rect 15102 5652 15108 5704
rect 15160 5652 15166 5704
rect 15212 5701 15240 5732
rect 15657 5729 15669 5763
rect 15703 5729 15715 5763
rect 16945 5763 17003 5769
rect 16945 5760 16957 5763
rect 15657 5723 15715 5729
rect 16316 5732 16957 5760
rect 16316 5704 16344 5732
rect 16945 5729 16957 5732
rect 16991 5729 17003 5763
rect 16945 5723 17003 5729
rect 17604 5732 18000 5760
rect 15197 5695 15255 5701
rect 15197 5661 15209 5695
rect 15243 5661 15255 5695
rect 15197 5655 15255 5661
rect 15286 5652 15292 5704
rect 15344 5692 15350 5704
rect 15381 5695 15439 5701
rect 15381 5692 15393 5695
rect 15344 5664 15393 5692
rect 15344 5652 15350 5664
rect 15381 5661 15393 5664
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 15672 5664 16252 5692
rect 14918 5624 14924 5636
rect 14108 5596 14924 5624
rect 14918 5584 14924 5596
rect 14976 5584 14982 5636
rect 15672 5624 15700 5664
rect 15580 5596 15700 5624
rect 16224 5624 16252 5664
rect 16298 5652 16304 5704
rect 16356 5652 16362 5704
rect 17604 5692 17632 5732
rect 16408 5664 17632 5692
rect 16408 5624 16436 5664
rect 17678 5652 17684 5704
rect 17736 5652 17742 5704
rect 17862 5652 17868 5704
rect 17920 5652 17926 5704
rect 17972 5692 18000 5732
rect 18874 5720 18880 5772
rect 18932 5760 18938 5772
rect 19153 5763 19211 5769
rect 19153 5760 19165 5763
rect 18932 5732 19165 5760
rect 18932 5720 18938 5732
rect 19153 5729 19165 5732
rect 19199 5729 19211 5763
rect 19153 5723 19211 5729
rect 19429 5763 19487 5769
rect 19429 5729 19441 5763
rect 19475 5760 19487 5763
rect 22554 5760 22560 5772
rect 19475 5732 22560 5760
rect 19475 5729 19487 5732
rect 19429 5723 19487 5729
rect 22554 5720 22560 5732
rect 22612 5720 22618 5772
rect 22925 5763 22983 5769
rect 22925 5729 22937 5763
rect 22971 5760 22983 5763
rect 23382 5760 23388 5772
rect 22971 5732 23388 5760
rect 22971 5729 22983 5732
rect 22925 5723 22983 5729
rect 23382 5720 23388 5732
rect 23440 5720 23446 5772
rect 23661 5763 23719 5769
rect 23661 5729 23673 5763
rect 23707 5760 23719 5763
rect 24302 5760 24308 5772
rect 23707 5732 24308 5760
rect 23707 5729 23719 5732
rect 23661 5723 23719 5729
rect 24302 5720 24308 5732
rect 24360 5720 24366 5772
rect 24504 5769 24532 5800
rect 24670 5788 24676 5800
rect 24728 5788 24734 5840
rect 24489 5763 24547 5769
rect 24489 5729 24501 5763
rect 24535 5729 24547 5763
rect 24489 5723 24547 5729
rect 20162 5692 20168 5704
rect 17972 5664 20168 5692
rect 20162 5652 20168 5664
rect 20220 5652 20226 5704
rect 20901 5695 20959 5701
rect 20901 5661 20913 5695
rect 20947 5692 20959 5695
rect 21174 5692 21180 5704
rect 20947 5664 21180 5692
rect 20947 5661 20959 5664
rect 20901 5655 20959 5661
rect 21174 5652 21180 5664
rect 21232 5652 21238 5704
rect 22186 5652 22192 5704
rect 22244 5652 22250 5704
rect 22373 5695 22431 5701
rect 22373 5661 22385 5695
rect 22419 5692 22431 5695
rect 23845 5695 23903 5701
rect 22419 5664 23796 5692
rect 22419 5661 22431 5664
rect 22373 5655 22431 5661
rect 16224 5596 16436 5624
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 6730 5556 6736 5568
rect 3936 5528 6736 5556
rect 3936 5516 3942 5528
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 9950 5516 9956 5568
rect 10008 5516 10014 5568
rect 12621 5559 12679 5565
rect 12621 5525 12633 5559
rect 12667 5556 12679 5559
rect 15580 5556 15608 5596
rect 16666 5584 16672 5636
rect 16724 5624 16730 5636
rect 23017 5627 23075 5633
rect 23017 5624 23029 5627
rect 16724 5596 23029 5624
rect 16724 5584 16730 5596
rect 23017 5593 23029 5596
rect 23063 5593 23075 5627
rect 23768 5624 23796 5664
rect 23845 5661 23857 5695
rect 23891 5692 23903 5695
rect 24210 5692 24216 5704
rect 23891 5664 24216 5692
rect 23891 5661 23903 5664
rect 23845 5655 23903 5661
rect 24210 5652 24216 5664
rect 24268 5652 24274 5704
rect 25056 5692 25084 5868
rect 26326 5856 26332 5868
rect 26384 5856 26390 5908
rect 26605 5899 26663 5905
rect 26605 5865 26617 5899
rect 26651 5896 26663 5899
rect 27062 5896 27068 5908
rect 26651 5868 27068 5896
rect 26651 5865 26663 5868
rect 26605 5859 26663 5865
rect 27062 5856 27068 5868
rect 27120 5856 27126 5908
rect 27430 5856 27436 5908
rect 27488 5896 27494 5908
rect 27488 5868 30236 5896
rect 27488 5856 27494 5868
rect 25130 5788 25136 5840
rect 25188 5828 25194 5840
rect 25188 5800 30051 5828
rect 25188 5788 25194 5800
rect 25314 5720 25320 5772
rect 25372 5720 25378 5772
rect 25498 5720 25504 5772
rect 25556 5720 25562 5772
rect 25777 5763 25835 5769
rect 25777 5729 25789 5763
rect 25823 5760 25835 5763
rect 25866 5760 25872 5772
rect 25823 5732 25872 5760
rect 25823 5729 25835 5732
rect 25777 5723 25835 5729
rect 25866 5720 25872 5732
rect 25924 5720 25930 5772
rect 25961 5763 26019 5769
rect 25961 5729 25973 5763
rect 26007 5729 26019 5763
rect 25961 5723 26019 5729
rect 24320 5664 25084 5692
rect 25593 5695 25651 5701
rect 24320 5624 24348 5664
rect 25593 5661 25605 5695
rect 25639 5661 25651 5695
rect 25593 5655 25651 5661
rect 23768 5596 24348 5624
rect 23017 5587 23075 5593
rect 25038 5584 25044 5636
rect 25096 5624 25102 5636
rect 25608 5624 25636 5655
rect 25682 5652 25688 5704
rect 25740 5652 25746 5704
rect 25976 5692 26004 5723
rect 27338 5720 27344 5772
rect 27396 5720 27402 5772
rect 28813 5763 28871 5769
rect 28813 5729 28825 5763
rect 28859 5760 28871 5763
rect 29454 5760 29460 5772
rect 28859 5732 29460 5760
rect 28859 5729 28871 5732
rect 28813 5723 28871 5729
rect 29454 5720 29460 5732
rect 29512 5720 29518 5772
rect 29546 5720 29552 5772
rect 29604 5720 29610 5772
rect 29641 5763 29699 5769
rect 29641 5729 29653 5763
rect 29687 5760 29699 5763
rect 29914 5760 29920 5772
rect 29687 5732 29920 5760
rect 29687 5729 29699 5732
rect 29641 5723 29699 5729
rect 29914 5720 29920 5732
rect 29972 5720 29978 5772
rect 26142 5692 26148 5704
rect 25976 5664 26148 5692
rect 26142 5652 26148 5664
rect 26200 5652 26206 5704
rect 28077 5695 28135 5701
rect 28077 5661 28089 5695
rect 28123 5692 28135 5695
rect 28123 5664 28672 5692
rect 28123 5661 28135 5664
rect 28077 5655 28135 5661
rect 25096 5596 25636 5624
rect 25096 5584 25102 5596
rect 25866 5584 25872 5636
rect 25924 5624 25930 5636
rect 28169 5627 28227 5633
rect 28169 5624 28181 5627
rect 25924 5596 28181 5624
rect 25924 5584 25930 5596
rect 28169 5593 28181 5596
rect 28215 5593 28227 5627
rect 28644 5624 28672 5664
rect 28902 5652 28908 5704
rect 28960 5702 28966 5704
rect 28960 5692 29316 5702
rect 30023 5692 30051 5800
rect 30208 5760 30236 5868
rect 30466 5856 30472 5908
rect 30524 5856 30530 5908
rect 31297 5899 31355 5905
rect 31297 5865 31309 5899
rect 31343 5896 31355 5899
rect 31938 5896 31944 5908
rect 31343 5868 31944 5896
rect 31343 5865 31355 5868
rect 31297 5859 31355 5865
rect 31938 5856 31944 5868
rect 31996 5856 32002 5908
rect 32493 5899 32551 5905
rect 32493 5865 32505 5899
rect 32539 5896 32551 5899
rect 32539 5868 32904 5896
rect 32539 5865 32551 5868
rect 32493 5859 32551 5865
rect 30285 5831 30343 5837
rect 30285 5797 30297 5831
rect 30331 5828 30343 5831
rect 32876 5828 32904 5868
rect 32950 5856 32956 5908
rect 33008 5896 33014 5908
rect 33778 5896 33784 5908
rect 33008 5868 33784 5896
rect 33008 5856 33014 5868
rect 33778 5856 33784 5868
rect 33836 5896 33842 5908
rect 33873 5899 33931 5905
rect 33873 5896 33885 5899
rect 33836 5868 33885 5896
rect 33836 5856 33842 5868
rect 33873 5865 33885 5868
rect 33919 5865 33931 5899
rect 35342 5896 35348 5908
rect 33873 5859 33931 5865
rect 33980 5868 35348 5896
rect 33980 5828 34008 5868
rect 35342 5856 35348 5868
rect 35400 5856 35406 5908
rect 36814 5856 36820 5908
rect 36872 5896 36878 5908
rect 37274 5896 37280 5908
rect 36872 5868 37280 5896
rect 36872 5856 36878 5868
rect 37274 5856 37280 5868
rect 37332 5856 37338 5908
rect 38654 5856 38660 5908
rect 38712 5896 38718 5908
rect 42981 5899 43039 5905
rect 42981 5896 42993 5899
rect 38712 5868 42993 5896
rect 38712 5856 38718 5868
rect 42981 5865 42993 5868
rect 43027 5865 43039 5899
rect 42981 5859 43039 5865
rect 30331 5800 32720 5828
rect 32876 5800 34008 5828
rect 30331 5797 30343 5800
rect 30285 5791 30343 5797
rect 30926 5760 30932 5772
rect 30208 5732 30932 5760
rect 30926 5720 30932 5732
rect 30984 5720 30990 5772
rect 31113 5763 31171 5769
rect 31113 5729 31125 5763
rect 31159 5729 31171 5763
rect 31113 5723 31171 5729
rect 31941 5763 31999 5769
rect 31941 5729 31953 5763
rect 31987 5760 31999 5763
rect 32030 5760 32036 5772
rect 31987 5732 32036 5760
rect 31987 5729 31999 5732
rect 31941 5723 31999 5729
rect 30837 5695 30895 5701
rect 30837 5692 30849 5695
rect 28960 5674 29684 5692
rect 28960 5664 28994 5674
rect 29288 5664 29684 5674
rect 30023 5664 30849 5692
rect 28960 5652 28966 5664
rect 29086 5624 29092 5636
rect 28644 5596 29092 5624
rect 28169 5587 28227 5593
rect 29086 5584 29092 5596
rect 29144 5584 29150 5636
rect 12667 5528 15608 5556
rect 12667 5525 12679 5528
rect 12621 5519 12679 5525
rect 16390 5516 16396 5568
rect 16448 5516 16454 5568
rect 17126 5516 17132 5568
rect 17184 5516 17190 5568
rect 18598 5516 18604 5568
rect 18656 5556 18662 5568
rect 18966 5556 18972 5568
rect 18656 5528 18972 5556
rect 18656 5516 18662 5528
rect 18966 5516 18972 5528
rect 19024 5516 19030 5568
rect 19150 5516 19156 5568
rect 19208 5556 19214 5568
rect 19886 5556 19892 5568
rect 19208 5528 19892 5556
rect 19208 5516 19214 5528
rect 19886 5516 19892 5528
rect 19944 5516 19950 5568
rect 19981 5559 20039 5565
rect 19981 5525 19993 5559
rect 20027 5556 20039 5559
rect 20070 5556 20076 5568
rect 20027 5528 20076 5556
rect 20027 5525 20039 5528
rect 19981 5519 20039 5525
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 20349 5559 20407 5565
rect 20349 5525 20361 5559
rect 20395 5556 20407 5559
rect 20806 5556 20812 5568
rect 20395 5528 20812 5556
rect 20395 5525 20407 5528
rect 20349 5519 20407 5525
rect 20806 5516 20812 5528
rect 20864 5516 20870 5568
rect 21545 5559 21603 5565
rect 21545 5525 21557 5559
rect 21591 5556 21603 5559
rect 21634 5556 21640 5568
rect 21591 5528 21640 5556
rect 21591 5525 21603 5528
rect 21545 5519 21603 5525
rect 21634 5516 21640 5528
rect 21692 5516 21698 5568
rect 22186 5516 22192 5568
rect 22244 5556 22250 5568
rect 24946 5556 24952 5568
rect 22244 5528 24952 5556
rect 22244 5516 22250 5528
rect 24946 5516 24952 5528
rect 25004 5516 25010 5568
rect 25133 5559 25191 5565
rect 25133 5525 25145 5559
rect 25179 5556 25191 5559
rect 25590 5556 25596 5568
rect 25179 5528 25596 5556
rect 25179 5525 25191 5528
rect 25133 5519 25191 5525
rect 25590 5516 25596 5528
rect 25648 5516 25654 5568
rect 26694 5516 26700 5568
rect 26752 5516 26758 5568
rect 27430 5516 27436 5568
rect 27488 5516 27494 5568
rect 28074 5516 28080 5568
rect 28132 5556 28138 5568
rect 28905 5559 28963 5565
rect 28905 5556 28917 5559
rect 28132 5528 28917 5556
rect 28132 5516 28138 5528
rect 28905 5525 28917 5528
rect 28951 5525 28963 5559
rect 29656 5556 29684 5664
rect 30837 5661 30849 5664
rect 30883 5661 30895 5695
rect 30837 5655 30895 5661
rect 31128 5556 31156 5723
rect 32030 5720 32036 5732
rect 32088 5720 32094 5772
rect 31481 5695 31539 5701
rect 31481 5661 31493 5695
rect 31527 5692 31539 5695
rect 31570 5692 31576 5704
rect 31527 5664 31576 5692
rect 31527 5661 31539 5664
rect 31481 5655 31539 5661
rect 31570 5652 31576 5664
rect 31628 5652 31634 5704
rect 31757 5695 31815 5701
rect 31757 5661 31769 5695
rect 31803 5692 31815 5695
rect 32214 5692 32220 5704
rect 31803 5664 32220 5692
rect 31803 5661 31815 5664
rect 31757 5655 31815 5661
rect 32214 5652 32220 5664
rect 32272 5652 32278 5704
rect 32582 5652 32588 5704
rect 32640 5652 32646 5704
rect 32692 5692 32720 5800
rect 34422 5788 34428 5840
rect 34480 5788 34486 5840
rect 34793 5831 34851 5837
rect 34793 5797 34805 5831
rect 34839 5828 34851 5831
rect 34974 5828 34980 5840
rect 34839 5800 34980 5828
rect 34839 5797 34851 5800
rect 34793 5791 34851 5797
rect 34974 5788 34980 5800
rect 35032 5788 35038 5840
rect 36446 5788 36452 5840
rect 36504 5828 36510 5840
rect 36504 5800 37044 5828
rect 36504 5788 36510 5800
rect 33520 5732 35204 5760
rect 33410 5692 33416 5704
rect 32692 5664 33416 5692
rect 33410 5652 33416 5664
rect 33468 5652 33474 5704
rect 31662 5584 31668 5636
rect 31720 5624 31726 5636
rect 32490 5624 32496 5636
rect 31720 5596 32496 5624
rect 31720 5584 31726 5596
rect 32490 5584 32496 5596
rect 32548 5584 32554 5636
rect 32858 5584 32864 5636
rect 32916 5624 32922 5636
rect 33520 5624 33548 5732
rect 34238 5652 34244 5704
rect 34296 5692 34302 5704
rect 34425 5695 34483 5701
rect 34425 5692 34437 5695
rect 34296 5664 34437 5692
rect 34296 5652 34302 5664
rect 34425 5661 34437 5664
rect 34471 5661 34483 5695
rect 34425 5655 34483 5661
rect 34514 5652 34520 5704
rect 34572 5652 34578 5704
rect 35066 5652 35072 5704
rect 35124 5652 35130 5704
rect 35176 5701 35204 5732
rect 35894 5720 35900 5772
rect 35952 5760 35958 5772
rect 35952 5732 36400 5760
rect 35952 5720 35958 5732
rect 35161 5695 35219 5701
rect 35161 5661 35173 5695
rect 35207 5661 35219 5695
rect 35161 5655 35219 5661
rect 35250 5652 35256 5704
rect 35308 5652 35314 5704
rect 35434 5652 35440 5704
rect 35492 5652 35498 5704
rect 35713 5695 35771 5701
rect 35713 5661 35725 5695
rect 35759 5692 35771 5695
rect 36262 5692 36268 5704
rect 35759 5664 36268 5692
rect 35759 5661 35771 5664
rect 35713 5655 35771 5661
rect 36262 5652 36268 5664
rect 36320 5652 36326 5704
rect 36372 5692 36400 5732
rect 36906 5720 36912 5772
rect 36964 5720 36970 5772
rect 37016 5760 37044 5800
rect 38838 5788 38844 5840
rect 38896 5828 38902 5840
rect 39666 5828 39672 5840
rect 38896 5800 39672 5828
rect 38896 5788 38902 5800
rect 39666 5788 39672 5800
rect 39724 5788 39730 5840
rect 42794 5828 42800 5840
rect 39776 5800 42800 5828
rect 37016 5732 39068 5760
rect 38933 5695 38991 5701
rect 38933 5692 38945 5695
rect 36372 5664 38945 5692
rect 38933 5661 38945 5664
rect 38979 5661 38991 5695
rect 39040 5692 39068 5732
rect 39298 5720 39304 5772
rect 39356 5720 39362 5772
rect 39776 5692 39804 5800
rect 42794 5788 42800 5800
rect 42852 5788 42858 5840
rect 41138 5720 41144 5772
rect 41196 5760 41202 5772
rect 42061 5763 42119 5769
rect 42061 5760 42073 5763
rect 41196 5732 42073 5760
rect 41196 5720 41202 5732
rect 42061 5729 42073 5732
rect 42107 5729 42119 5763
rect 42061 5723 42119 5729
rect 42978 5720 42984 5772
rect 43036 5760 43042 5772
rect 44453 5763 44511 5769
rect 44453 5760 44465 5763
rect 43036 5732 44465 5760
rect 43036 5720 43042 5732
rect 44453 5729 44465 5732
rect 44499 5729 44511 5763
rect 44453 5723 44511 5729
rect 45186 5720 45192 5772
rect 45244 5760 45250 5772
rect 45925 5763 45983 5769
rect 45925 5760 45937 5763
rect 45244 5732 45937 5760
rect 45244 5720 45250 5732
rect 45925 5729 45937 5732
rect 45971 5729 45983 5763
rect 45925 5723 45983 5729
rect 39040 5664 39804 5692
rect 39853 5695 39911 5701
rect 38933 5655 38991 5661
rect 39853 5661 39865 5695
rect 39899 5692 39911 5695
rect 40497 5695 40555 5701
rect 40497 5692 40509 5695
rect 39899 5664 40509 5692
rect 39899 5661 39911 5664
rect 39853 5655 39911 5661
rect 40497 5661 40509 5664
rect 40543 5661 40555 5695
rect 40497 5655 40555 5661
rect 41417 5695 41475 5701
rect 41417 5661 41429 5695
rect 41463 5692 41475 5695
rect 41509 5695 41567 5701
rect 41509 5692 41521 5695
rect 41463 5664 41521 5692
rect 41463 5661 41475 5664
rect 41417 5655 41475 5661
rect 41509 5661 41521 5664
rect 41555 5661 41567 5695
rect 41509 5655 41567 5661
rect 42886 5652 42892 5704
rect 42944 5652 42950 5704
rect 43625 5695 43683 5701
rect 43625 5661 43637 5695
rect 43671 5661 43683 5695
rect 43625 5655 43683 5661
rect 32916 5596 33548 5624
rect 32916 5584 32922 5596
rect 34606 5584 34612 5636
rect 34664 5624 34670 5636
rect 34701 5627 34759 5633
rect 34701 5624 34713 5627
rect 34664 5596 34713 5624
rect 34664 5584 34670 5596
rect 34701 5593 34713 5596
rect 34747 5593 34759 5627
rect 34701 5587 34759 5593
rect 35802 5584 35808 5636
rect 35860 5624 35866 5636
rect 36357 5627 36415 5633
rect 36357 5624 36369 5627
rect 35860 5596 36369 5624
rect 35860 5584 35866 5596
rect 36357 5593 36369 5596
rect 36403 5593 36415 5627
rect 36357 5587 36415 5593
rect 36446 5584 36452 5636
rect 36504 5624 36510 5636
rect 37093 5627 37151 5633
rect 37093 5624 37105 5627
rect 36504 5596 37105 5624
rect 36504 5584 36510 5596
rect 37093 5593 37105 5596
rect 37139 5593 37151 5627
rect 37093 5587 37151 5593
rect 37274 5584 37280 5636
rect 37332 5624 37338 5636
rect 42245 5627 42303 5633
rect 42245 5624 42257 5627
rect 37332 5596 42257 5624
rect 37332 5584 37338 5596
rect 42245 5593 42257 5596
rect 42291 5593 42303 5627
rect 43640 5624 43668 5655
rect 44358 5652 44364 5704
rect 44416 5652 44422 5704
rect 45097 5695 45155 5701
rect 45097 5661 45109 5695
rect 45143 5692 45155 5695
rect 45830 5692 45836 5704
rect 45143 5664 45836 5692
rect 45143 5661 45155 5664
rect 45097 5655 45155 5661
rect 45830 5652 45836 5664
rect 45888 5652 45894 5704
rect 45646 5624 45652 5636
rect 43640 5596 45652 5624
rect 42245 5587 42303 5593
rect 45646 5584 45652 5596
rect 45704 5584 45710 5636
rect 36170 5556 36176 5568
rect 29656 5528 36176 5556
rect 28905 5519 28963 5525
rect 36170 5516 36176 5528
rect 36228 5516 36234 5568
rect 36265 5559 36323 5565
rect 36265 5525 36277 5559
rect 36311 5556 36323 5559
rect 37826 5556 37832 5568
rect 36311 5528 37832 5556
rect 36311 5525 36323 5528
rect 36265 5519 36323 5525
rect 37826 5516 37832 5528
rect 37884 5516 37890 5568
rect 37918 5516 37924 5568
rect 37976 5556 37982 5568
rect 38381 5559 38439 5565
rect 38381 5556 38393 5559
rect 37976 5528 38393 5556
rect 37976 5516 37982 5528
rect 38381 5525 38393 5528
rect 38427 5525 38439 5559
rect 38381 5519 38439 5525
rect 38930 5516 38936 5568
rect 38988 5556 38994 5568
rect 39025 5559 39083 5565
rect 39025 5556 39037 5559
rect 38988 5528 39037 5556
rect 38988 5516 38994 5528
rect 39025 5525 39037 5528
rect 39071 5525 39083 5559
rect 39025 5519 39083 5525
rect 39942 5516 39948 5568
rect 40000 5516 40006 5568
rect 40770 5516 40776 5568
rect 40828 5516 40834 5568
rect 43714 5516 43720 5568
rect 43772 5516 43778 5568
rect 46569 5559 46627 5565
rect 46569 5525 46581 5559
rect 46615 5556 46627 5559
rect 47026 5556 47032 5568
rect 46615 5528 47032 5556
rect 46615 5525 46627 5528
rect 46569 5519 46627 5525
rect 47026 5516 47032 5528
rect 47084 5516 47090 5568
rect 2024 5466 77924 5488
rect 2024 5414 5794 5466
rect 5846 5414 5858 5466
rect 5910 5414 5922 5466
rect 5974 5414 5986 5466
rect 6038 5414 6050 5466
rect 6102 5414 36514 5466
rect 36566 5414 36578 5466
rect 36630 5414 36642 5466
rect 36694 5414 36706 5466
rect 36758 5414 36770 5466
rect 36822 5414 67234 5466
rect 67286 5414 67298 5466
rect 67350 5414 67362 5466
rect 67414 5414 67426 5466
rect 67478 5414 67490 5466
rect 67542 5414 77924 5466
rect 2024 5392 77924 5414
rect 8389 5355 8447 5361
rect 8389 5321 8401 5355
rect 8435 5352 8447 5355
rect 9030 5352 9036 5364
rect 8435 5324 9036 5352
rect 8435 5321 8447 5324
rect 8389 5315 8447 5321
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9122 5312 9128 5364
rect 9180 5312 9186 5364
rect 11514 5312 11520 5364
rect 11572 5312 11578 5364
rect 12250 5312 12256 5364
rect 12308 5312 12314 5364
rect 12621 5355 12679 5361
rect 12621 5321 12633 5355
rect 12667 5352 12679 5355
rect 13354 5352 13360 5364
rect 12667 5324 13360 5352
rect 12667 5321 12679 5324
rect 12621 5315 12679 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 15197 5355 15255 5361
rect 15197 5321 15209 5355
rect 15243 5352 15255 5355
rect 15562 5352 15568 5364
rect 15243 5324 15568 5352
rect 15243 5321 15255 5324
rect 15197 5315 15255 5321
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 16117 5355 16175 5361
rect 16117 5321 16129 5355
rect 16163 5352 16175 5355
rect 16206 5352 16212 5364
rect 16163 5324 16212 5352
rect 16163 5321 16175 5324
rect 16117 5315 16175 5321
rect 16206 5312 16212 5324
rect 16264 5352 16270 5364
rect 16942 5352 16948 5364
rect 16264 5324 16948 5352
rect 16264 5312 16270 5324
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 17218 5312 17224 5364
rect 17276 5352 17282 5364
rect 17678 5352 17684 5364
rect 17276 5324 17684 5352
rect 17276 5312 17282 5324
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18230 5352 18236 5364
rect 18012 5324 18236 5352
rect 18012 5312 18018 5324
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 20254 5352 20260 5364
rect 18984 5324 20260 5352
rect 7098 5244 7104 5296
rect 7156 5284 7162 5296
rect 9953 5287 10011 5293
rect 9953 5284 9965 5287
rect 7156 5256 9965 5284
rect 7156 5244 7162 5256
rect 9953 5253 9965 5256
rect 9999 5253 10011 5287
rect 9953 5247 10011 5253
rect 13541 5287 13599 5293
rect 13541 5253 13553 5287
rect 13587 5284 13599 5287
rect 16482 5284 16488 5296
rect 13587 5256 16488 5284
rect 13587 5253 13599 5256
rect 13541 5247 13599 5253
rect 16482 5244 16488 5256
rect 16540 5244 16546 5296
rect 16666 5244 16672 5296
rect 16724 5244 16730 5296
rect 18322 5244 18328 5296
rect 18380 5284 18386 5296
rect 18506 5284 18512 5296
rect 18380 5256 18512 5284
rect 18380 5244 18386 5256
rect 18506 5244 18512 5256
rect 18564 5244 18570 5296
rect 7466 5176 7472 5228
rect 7524 5176 7530 5228
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5216 8631 5219
rect 8662 5216 8668 5228
rect 8619 5188 8668 5216
rect 8619 5185 8631 5188
rect 8573 5179 8631 5185
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5216 9827 5219
rect 10042 5216 10048 5228
rect 9815 5188 10048 5216
rect 9815 5185 9827 5188
rect 9769 5179 9827 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 11698 5176 11704 5228
rect 11756 5176 11762 5228
rect 12434 5176 12440 5228
rect 12492 5176 12498 5228
rect 13725 5219 13783 5225
rect 13725 5185 13737 5219
rect 13771 5216 13783 5219
rect 16022 5216 16028 5228
rect 13771 5188 16028 5216
rect 13771 5185 13783 5188
rect 13725 5179 13783 5185
rect 16022 5176 16028 5188
rect 16080 5176 16086 5228
rect 16393 5219 16451 5225
rect 16393 5185 16405 5219
rect 16439 5216 16451 5219
rect 17681 5219 17739 5225
rect 16439 5188 16528 5216
rect 16439 5185 16451 5188
rect 16393 5179 16451 5185
rect 16500 5160 16528 5188
rect 17681 5185 17693 5219
rect 17727 5216 17739 5219
rect 18984 5216 19012 5324
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 20714 5312 20720 5364
rect 20772 5352 20778 5364
rect 20809 5355 20867 5361
rect 20809 5352 20821 5355
rect 20772 5324 20821 5352
rect 20772 5312 20778 5324
rect 20809 5321 20821 5324
rect 20855 5321 20867 5355
rect 20809 5315 20867 5321
rect 21269 5355 21327 5361
rect 21269 5321 21281 5355
rect 21315 5352 21327 5355
rect 21358 5352 21364 5364
rect 21315 5324 21364 5352
rect 21315 5321 21327 5324
rect 21269 5315 21327 5321
rect 21358 5312 21364 5324
rect 21416 5312 21422 5364
rect 21821 5355 21879 5361
rect 21821 5321 21833 5355
rect 21867 5352 21879 5355
rect 21910 5352 21916 5364
rect 21867 5324 21916 5352
rect 21867 5321 21879 5324
rect 21821 5315 21879 5321
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 22557 5355 22615 5361
rect 22557 5321 22569 5355
rect 22603 5352 22615 5355
rect 23014 5352 23020 5364
rect 22603 5324 23020 5352
rect 22603 5321 22615 5324
rect 22557 5315 22615 5321
rect 23014 5312 23020 5324
rect 23072 5312 23078 5364
rect 23474 5312 23480 5364
rect 23532 5352 23538 5364
rect 24029 5355 24087 5361
rect 24029 5352 24041 5355
rect 23532 5324 24041 5352
rect 23532 5312 23538 5324
rect 24029 5321 24041 5324
rect 24075 5352 24087 5355
rect 24210 5352 24216 5364
rect 24075 5324 24216 5352
rect 24075 5321 24087 5324
rect 24029 5315 24087 5321
rect 24210 5312 24216 5324
rect 24268 5312 24274 5364
rect 25498 5312 25504 5364
rect 25556 5312 25562 5364
rect 26142 5312 26148 5364
rect 26200 5352 26206 5364
rect 26418 5352 26424 5364
rect 26200 5324 26424 5352
rect 26200 5312 26206 5324
rect 26418 5312 26424 5324
rect 26476 5312 26482 5364
rect 29549 5355 29607 5361
rect 29549 5321 29561 5355
rect 29595 5352 29607 5355
rect 29730 5352 29736 5364
rect 29595 5324 29736 5352
rect 29595 5321 29607 5324
rect 29549 5315 29607 5321
rect 29730 5312 29736 5324
rect 29788 5312 29794 5364
rect 30282 5312 30288 5364
rect 30340 5312 30346 5364
rect 32769 5355 32827 5361
rect 32769 5321 32781 5355
rect 32815 5352 32827 5355
rect 33318 5352 33324 5364
rect 32815 5324 33324 5352
rect 32815 5321 32827 5324
rect 32769 5315 32827 5321
rect 33318 5312 33324 5324
rect 33376 5312 33382 5364
rect 33594 5312 33600 5364
rect 33652 5312 33658 5364
rect 35158 5312 35164 5364
rect 35216 5312 35222 5364
rect 36170 5312 36176 5364
rect 36228 5352 36234 5364
rect 36446 5352 36452 5364
rect 36228 5324 36452 5352
rect 36228 5312 36234 5324
rect 36446 5312 36452 5324
rect 36504 5312 36510 5364
rect 36541 5355 36599 5361
rect 36541 5321 36553 5355
rect 36587 5352 36599 5355
rect 36998 5352 37004 5364
rect 36587 5324 37004 5352
rect 36587 5321 36599 5324
rect 36541 5315 36599 5321
rect 36998 5312 37004 5324
rect 37056 5312 37062 5364
rect 38930 5352 38936 5364
rect 37384 5324 38936 5352
rect 19242 5244 19248 5296
rect 19300 5244 19306 5296
rect 20530 5244 20536 5296
rect 20588 5284 20594 5296
rect 20588 5256 21956 5284
rect 20588 5244 20594 5256
rect 20806 5216 20812 5228
rect 17727 5188 19012 5216
rect 20378 5188 20812 5216
rect 17727 5185 17739 5188
rect 17681 5179 17739 5185
rect 20806 5176 20812 5188
rect 20864 5216 20870 5228
rect 21082 5216 21088 5228
rect 20864 5188 21088 5216
rect 20864 5176 20870 5188
rect 21082 5176 21088 5188
rect 21140 5176 21146 5228
rect 21177 5219 21235 5225
rect 21177 5185 21189 5219
rect 21223 5216 21235 5219
rect 21542 5216 21548 5228
rect 21223 5188 21548 5216
rect 21223 5185 21235 5188
rect 21177 5179 21235 5185
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5148 7895 5151
rect 9674 5148 9680 5160
rect 7883 5120 9680 5148
rect 7883 5117 7895 5120
rect 7837 5111 7895 5117
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 9858 5108 9864 5160
rect 9916 5148 9922 5160
rect 10505 5151 10563 5157
rect 10505 5148 10517 5151
rect 9916 5120 10517 5148
rect 9916 5108 9922 5120
rect 10505 5117 10517 5120
rect 10551 5117 10563 5151
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10505 5111 10563 5117
rect 10704 5120 10885 5148
rect 8386 5040 8392 5092
rect 8444 5080 8450 5092
rect 9217 5083 9275 5089
rect 9217 5080 9229 5083
rect 8444 5052 9229 5080
rect 8444 5040 8450 5052
rect 9217 5049 9229 5052
rect 9263 5049 9275 5083
rect 9217 5043 9275 5049
rect 10704 5024 10732 5120
rect 10873 5117 10885 5120
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 12989 5151 13047 5157
rect 12989 5117 13001 5151
rect 13035 5148 13047 5151
rect 13998 5148 14004 5160
rect 13035 5120 14004 5148
rect 13035 5117 13047 5120
rect 12989 5111 13047 5117
rect 13998 5108 14004 5120
rect 14056 5108 14062 5160
rect 14461 5151 14519 5157
rect 14461 5117 14473 5151
rect 14507 5148 14519 5151
rect 14642 5148 14648 5160
rect 14507 5120 14648 5148
rect 14507 5117 14519 5120
rect 14461 5111 14519 5117
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5148 15991 5151
rect 16206 5148 16212 5160
rect 15979 5120 16212 5148
rect 15979 5117 15991 5120
rect 15933 5111 15991 5117
rect 16206 5108 16212 5120
rect 16264 5108 16270 5160
rect 16482 5108 16488 5160
rect 16540 5108 16546 5160
rect 16577 5151 16635 5157
rect 16577 5117 16589 5151
rect 16623 5148 16635 5151
rect 16623 5120 16712 5148
rect 16623 5117 16635 5120
rect 16577 5111 16635 5117
rect 16684 5092 16712 5120
rect 16758 5108 16764 5160
rect 16816 5108 16822 5160
rect 17770 5108 17776 5160
rect 17828 5108 17834 5160
rect 17862 5108 17868 5160
rect 17920 5108 17926 5160
rect 17957 5151 18015 5157
rect 17957 5117 17969 5151
rect 18003 5148 18015 5151
rect 18230 5148 18236 5160
rect 18003 5120 18236 5148
rect 18003 5117 18015 5120
rect 17957 5111 18015 5117
rect 18230 5108 18236 5120
rect 18288 5108 18294 5160
rect 18325 5151 18383 5157
rect 18325 5117 18337 5151
rect 18371 5148 18383 5151
rect 18506 5148 18512 5160
rect 18371 5120 18512 5148
rect 18371 5117 18383 5120
rect 18325 5111 18383 5117
rect 18506 5108 18512 5120
rect 18564 5108 18570 5160
rect 18598 5108 18604 5160
rect 18656 5148 18662 5160
rect 18969 5151 19027 5157
rect 18969 5148 18981 5151
rect 18656 5120 18981 5148
rect 18656 5108 18662 5120
rect 18969 5117 18981 5120
rect 19015 5117 19027 5151
rect 18969 5111 19027 5117
rect 20717 5151 20775 5157
rect 20717 5117 20729 5151
rect 20763 5148 20775 5151
rect 21192 5148 21220 5179
rect 21542 5176 21548 5188
rect 21600 5176 21606 5228
rect 21634 5176 21640 5228
rect 21692 5176 21698 5228
rect 21928 5225 21956 5256
rect 22738 5244 22744 5296
rect 22796 5284 22802 5296
rect 29638 5284 29644 5296
rect 22796 5256 28028 5284
rect 22796 5244 22802 5256
rect 21913 5219 21971 5225
rect 21913 5185 21925 5219
rect 21959 5185 21971 5219
rect 21913 5179 21971 5185
rect 23842 5176 23848 5228
rect 23900 5216 23906 5228
rect 24765 5219 24823 5225
rect 24765 5216 24777 5219
rect 23900 5188 24777 5216
rect 23900 5176 23906 5188
rect 24765 5185 24777 5188
rect 24811 5216 24823 5219
rect 24854 5216 24860 5228
rect 24811 5188 24860 5216
rect 24811 5185 24823 5188
rect 24765 5179 24823 5185
rect 24854 5176 24860 5188
rect 24912 5176 24918 5228
rect 24949 5219 25007 5225
rect 24949 5185 24961 5219
rect 24995 5216 25007 5219
rect 25866 5216 25872 5228
rect 24995 5188 25872 5216
rect 24995 5185 25007 5188
rect 24949 5179 25007 5185
rect 25866 5176 25872 5188
rect 25924 5176 25930 5228
rect 26421 5219 26479 5225
rect 26421 5185 26433 5219
rect 26467 5216 26479 5219
rect 26467 5188 27844 5216
rect 26467 5185 26479 5188
rect 26421 5179 26479 5185
rect 20763 5120 21220 5148
rect 20763 5117 20775 5120
rect 20717 5111 20775 5117
rect 21358 5108 21364 5160
rect 21416 5108 21422 5160
rect 25685 5151 25743 5157
rect 25685 5117 25697 5151
rect 25731 5117 25743 5151
rect 25685 5111 25743 5117
rect 27157 5151 27215 5157
rect 27157 5117 27169 5151
rect 27203 5148 27215 5151
rect 27338 5148 27344 5160
rect 27203 5120 27344 5148
rect 27203 5117 27215 5120
rect 27157 5111 27215 5117
rect 11054 5040 11060 5092
rect 11112 5080 11118 5092
rect 12710 5080 12716 5092
rect 11112 5052 12716 5080
rect 11112 5040 11118 5052
rect 12710 5040 12716 5052
rect 12768 5040 12774 5092
rect 12802 5040 12808 5092
rect 12860 5080 12866 5092
rect 15289 5083 15347 5089
rect 15289 5080 15301 5083
rect 12860 5052 15301 5080
rect 12860 5040 12866 5052
rect 15289 5049 15301 5052
rect 15335 5049 15347 5083
rect 15289 5043 15347 5049
rect 16666 5040 16672 5092
rect 16724 5040 16730 5092
rect 23382 5080 23388 5092
rect 17328 5052 19012 5080
rect 7653 5015 7711 5021
rect 7653 4981 7665 5015
rect 7699 5012 7711 5015
rect 8294 5012 8300 5024
rect 7699 4984 8300 5012
rect 7699 4981 7711 4984
rect 7653 4975 7711 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 10686 4972 10692 5024
rect 10744 4972 10750 5024
rect 10870 4972 10876 5024
rect 10928 5012 10934 5024
rect 13446 5012 13452 5024
rect 10928 4984 13452 5012
rect 10928 4972 10934 4984
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 14274 4972 14280 5024
rect 14332 4972 14338 5024
rect 16206 4972 16212 5024
rect 16264 4972 16270 5024
rect 16577 5015 16635 5021
rect 16577 4981 16589 5015
rect 16623 5012 16635 5015
rect 17328 5012 17356 5052
rect 16623 4984 17356 5012
rect 17405 5015 17463 5021
rect 16623 4981 16635 4984
rect 16577 4975 16635 4981
rect 17405 4981 17417 5015
rect 17451 5012 17463 5015
rect 17770 5012 17776 5024
rect 17451 4984 17776 5012
rect 17451 4981 17463 4984
rect 17405 4975 17463 4981
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18046 4972 18052 5024
rect 18104 5012 18110 5024
rect 18141 5015 18199 5021
rect 18141 5012 18153 5015
rect 18104 4984 18153 5012
rect 18104 4972 18110 4984
rect 18141 4981 18153 4984
rect 18187 4981 18199 5015
rect 18141 4975 18199 4981
rect 18322 4972 18328 5024
rect 18380 5012 18386 5024
rect 18690 5012 18696 5024
rect 18380 4984 18696 5012
rect 18380 4972 18386 4984
rect 18690 4972 18696 4984
rect 18748 4972 18754 5024
rect 18874 4972 18880 5024
rect 18932 4972 18938 5024
rect 18984 5012 19012 5052
rect 20272 5052 23388 5080
rect 20272 5012 20300 5052
rect 23382 5040 23388 5052
rect 23440 5040 23446 5092
rect 23566 5040 23572 5092
rect 23624 5080 23630 5092
rect 24394 5080 24400 5092
rect 23624 5052 24400 5080
rect 23624 5040 23630 5052
rect 24394 5040 24400 5052
rect 24452 5040 24458 5092
rect 18984 4984 20300 5012
rect 23106 4972 23112 5024
rect 23164 5012 23170 5024
rect 24581 5015 24639 5021
rect 24581 5012 24593 5015
rect 23164 4984 24593 5012
rect 23164 4972 23170 4984
rect 24581 4981 24593 4984
rect 24627 4981 24639 5015
rect 25700 5012 25728 5111
rect 27338 5108 27344 5120
rect 27396 5108 27402 5160
rect 27816 5148 27844 5188
rect 27890 5176 27896 5228
rect 27948 5176 27954 5228
rect 28000 5216 28028 5256
rect 28460 5256 29644 5284
rect 28460 5216 28488 5256
rect 29638 5244 29644 5256
rect 29696 5244 29702 5296
rect 30837 5287 30895 5293
rect 30837 5284 30849 5287
rect 29748 5256 30849 5284
rect 28000 5188 28488 5216
rect 28534 5176 28540 5228
rect 28592 5216 28598 5228
rect 29748 5216 29776 5256
rect 30837 5253 30849 5256
rect 30883 5253 30895 5287
rect 30837 5247 30895 5253
rect 31294 5244 31300 5296
rect 31352 5244 31358 5296
rect 32398 5244 32404 5296
rect 32456 5284 32462 5296
rect 32456 5256 33088 5284
rect 32456 5244 32462 5256
rect 28592 5188 29776 5216
rect 28592 5176 28598 5188
rect 32122 5176 32128 5228
rect 32180 5216 32186 5228
rect 33060 5225 33088 5256
rect 33134 5244 33140 5296
rect 33192 5284 33198 5296
rect 33229 5287 33287 5293
rect 33229 5284 33241 5287
rect 33192 5256 33241 5284
rect 33192 5244 33198 5256
rect 33229 5253 33241 5256
rect 33275 5253 33287 5287
rect 34330 5284 34336 5296
rect 33229 5247 33287 5253
rect 33336 5256 34336 5284
rect 33336 5225 33364 5256
rect 34330 5244 34336 5256
rect 34388 5244 34394 5296
rect 35250 5244 35256 5296
rect 35308 5284 35314 5296
rect 36633 5287 36691 5293
rect 36633 5284 36645 5287
rect 35308 5256 36645 5284
rect 35308 5244 35314 5256
rect 36633 5253 36645 5256
rect 36679 5253 36691 5287
rect 36633 5247 36691 5253
rect 36814 5244 36820 5296
rect 36872 5284 36878 5296
rect 37384 5284 37412 5324
rect 38930 5312 38936 5324
rect 38988 5312 38994 5364
rect 41509 5355 41567 5361
rect 41509 5321 41521 5355
rect 41555 5352 41567 5355
rect 42702 5352 42708 5364
rect 41555 5324 42708 5352
rect 41555 5321 41567 5324
rect 41509 5315 41567 5321
rect 42702 5312 42708 5324
rect 42760 5312 42766 5364
rect 36872 5256 37412 5284
rect 36872 5244 36878 5256
rect 37458 5244 37464 5296
rect 37516 5284 37522 5296
rect 37516 5256 41000 5284
rect 37516 5244 37522 5256
rect 32585 5219 32643 5225
rect 32585 5216 32597 5219
rect 32180 5188 32597 5216
rect 32180 5176 32186 5188
rect 32585 5185 32597 5188
rect 32631 5185 32643 5219
rect 32585 5179 32643 5185
rect 32861 5219 32919 5225
rect 32861 5185 32873 5219
rect 32907 5185 32919 5219
rect 32861 5179 32919 5185
rect 33045 5219 33103 5225
rect 33045 5185 33057 5219
rect 33091 5185 33103 5219
rect 33045 5179 33103 5185
rect 33321 5219 33379 5225
rect 33321 5185 33333 5219
rect 33367 5185 33379 5219
rect 33321 5179 33379 5185
rect 28261 5151 28319 5157
rect 27816 5120 28120 5148
rect 26237 5083 26295 5089
rect 26237 5049 26249 5083
rect 26283 5080 26295 5083
rect 27890 5080 27896 5092
rect 26283 5052 27896 5080
rect 26283 5049 26295 5052
rect 26237 5043 26295 5049
rect 27890 5040 27896 5052
rect 27948 5040 27954 5092
rect 28092 5080 28120 5120
rect 28261 5117 28273 5151
rect 28307 5148 28319 5151
rect 28350 5148 28356 5160
rect 28307 5120 28356 5148
rect 28307 5117 28319 5120
rect 28261 5111 28319 5117
rect 28350 5108 28356 5120
rect 28408 5108 28414 5160
rect 28810 5108 28816 5160
rect 28868 5148 28874 5160
rect 28905 5151 28963 5157
rect 28905 5148 28917 5151
rect 28868 5120 28917 5148
rect 28868 5108 28874 5120
rect 28905 5117 28917 5120
rect 28951 5117 28963 5151
rect 28905 5111 28963 5117
rect 29733 5151 29791 5157
rect 29733 5117 29745 5151
rect 29779 5117 29791 5151
rect 29733 5111 29791 5117
rect 30561 5151 30619 5157
rect 30561 5117 30573 5151
rect 30607 5148 30619 5151
rect 32030 5148 32036 5160
rect 30607 5120 32036 5148
rect 30607 5117 30619 5120
rect 30561 5111 30619 5117
rect 29638 5080 29644 5092
rect 28092 5052 29644 5080
rect 29638 5040 29644 5052
rect 29696 5040 29702 5092
rect 29748 5080 29776 5111
rect 32030 5108 32036 5120
rect 32088 5108 32094 5160
rect 32876 5148 32904 5179
rect 33410 5176 33416 5228
rect 33468 5176 33474 5228
rect 34790 5216 34796 5228
rect 33520 5188 34796 5216
rect 33520 5148 33548 5188
rect 34790 5176 34796 5188
rect 34848 5176 34854 5228
rect 35069 5219 35127 5225
rect 35069 5185 35081 5219
rect 35115 5216 35127 5219
rect 35526 5216 35532 5228
rect 35115 5188 35532 5216
rect 35115 5185 35127 5188
rect 35069 5179 35127 5185
rect 35526 5176 35532 5188
rect 35584 5176 35590 5228
rect 35802 5176 35808 5228
rect 35860 5176 35866 5228
rect 35897 5219 35955 5225
rect 35897 5185 35909 5219
rect 35943 5185 35955 5219
rect 35897 5179 35955 5185
rect 32876 5120 33548 5148
rect 33686 5108 33692 5160
rect 33744 5108 33750 5160
rect 34146 5108 34152 5160
rect 34204 5148 34210 5160
rect 35912 5148 35940 5179
rect 36078 5176 36084 5228
rect 36136 5176 36142 5228
rect 36170 5176 36176 5228
rect 36228 5176 36234 5228
rect 36265 5219 36323 5225
rect 36265 5185 36277 5219
rect 36311 5216 36323 5219
rect 36906 5216 36912 5228
rect 36311 5188 36912 5216
rect 36311 5185 36323 5188
rect 36265 5179 36323 5185
rect 36906 5176 36912 5188
rect 36964 5176 36970 5228
rect 37016 5188 38056 5216
rect 36538 5148 36544 5160
rect 34204 5120 34560 5148
rect 35912 5120 36544 5148
rect 34204 5108 34210 5120
rect 29748 5052 30696 5080
rect 26878 5012 26884 5024
rect 25700 4984 26884 5012
rect 24581 4975 24639 4981
rect 26878 4972 26884 4984
rect 26936 4972 26942 5024
rect 26970 4972 26976 5024
rect 27028 4972 27034 5024
rect 27706 4972 27712 5024
rect 27764 4972 27770 5024
rect 28077 5015 28135 5021
rect 28077 4981 28089 5015
rect 28123 5012 28135 5015
rect 28258 5012 28264 5024
rect 28123 4984 28264 5012
rect 28123 4981 28135 4984
rect 28077 4975 28135 4981
rect 28258 4972 28264 4984
rect 28316 4972 28322 5024
rect 28813 5015 28871 5021
rect 28813 4981 28825 5015
rect 28859 5012 28871 5015
rect 30466 5012 30472 5024
rect 28859 4984 30472 5012
rect 28859 4981 28871 4984
rect 28813 4975 28871 4981
rect 30466 4972 30472 4984
rect 30524 4972 30530 5024
rect 30668 5012 30696 5052
rect 32214 5040 32220 5092
rect 32272 5080 32278 5092
rect 34425 5083 34483 5089
rect 34425 5080 34437 5083
rect 32272 5052 34437 5080
rect 32272 5040 32278 5052
rect 34425 5049 34437 5052
rect 34471 5049 34483 5083
rect 34532 5080 34560 5120
rect 36538 5108 36544 5120
rect 36596 5108 36602 5160
rect 37016 5080 37044 5188
rect 37277 5151 37335 5157
rect 37277 5117 37289 5151
rect 37323 5117 37335 5151
rect 37277 5111 37335 5117
rect 34532 5052 37044 5080
rect 37292 5080 37320 5111
rect 37734 5108 37740 5160
rect 37792 5148 37798 5160
rect 37921 5151 37979 5157
rect 37921 5148 37933 5151
rect 37792 5120 37933 5148
rect 37792 5108 37798 5120
rect 37921 5117 37933 5120
rect 37967 5117 37979 5151
rect 38028 5148 38056 5188
rect 38194 5176 38200 5228
rect 38252 5176 38258 5228
rect 38381 5219 38439 5225
rect 38381 5185 38393 5219
rect 38427 5216 38439 5219
rect 39485 5219 39543 5225
rect 38427 5188 39252 5216
rect 38427 5185 38439 5188
rect 38381 5179 38439 5185
rect 38657 5151 38715 5157
rect 38657 5148 38669 5151
rect 38028 5120 38669 5148
rect 37921 5111 37979 5117
rect 38657 5117 38669 5120
rect 38703 5117 38715 5151
rect 38657 5111 38715 5117
rect 38565 5083 38623 5089
rect 38565 5080 38577 5083
rect 37292 5052 38577 5080
rect 34425 5043 34483 5049
rect 38565 5049 38577 5052
rect 38611 5049 38623 5083
rect 38565 5043 38623 5049
rect 32030 5012 32036 5024
rect 30668 4984 32036 5012
rect 32030 4972 32036 4984
rect 32088 4972 32094 5024
rect 32766 4972 32772 5024
rect 32824 5012 32830 5024
rect 33410 5012 33416 5024
rect 32824 4984 33416 5012
rect 32824 4972 32830 4984
rect 33410 4972 33416 4984
rect 33468 4972 33474 5024
rect 34333 5015 34391 5021
rect 34333 4981 34345 5015
rect 34379 5012 34391 5015
rect 37274 5012 37280 5024
rect 34379 4984 37280 5012
rect 34379 4981 34391 4984
rect 34333 4975 34391 4981
rect 37274 4972 37280 4984
rect 37332 4972 37338 5024
rect 37366 4972 37372 5024
rect 37424 4972 37430 5024
rect 39224 5012 39252 5188
rect 39485 5185 39497 5219
rect 39531 5216 39543 5219
rect 39942 5216 39948 5228
rect 39531 5188 39948 5216
rect 39531 5185 39543 5188
rect 39485 5179 39543 5185
rect 39942 5176 39948 5188
rect 40000 5176 40006 5228
rect 40770 5176 40776 5228
rect 40828 5216 40834 5228
rect 40865 5219 40923 5225
rect 40865 5216 40877 5219
rect 40828 5188 40877 5216
rect 40828 5176 40834 5188
rect 40865 5185 40877 5188
rect 40911 5185 40923 5219
rect 40865 5179 40923 5185
rect 39301 5151 39359 5157
rect 39301 5117 39313 5151
rect 39347 5117 39359 5151
rect 39301 5111 39359 5117
rect 40037 5151 40095 5157
rect 40037 5117 40049 5151
rect 40083 5148 40095 5151
rect 40681 5151 40739 5157
rect 40681 5148 40693 5151
rect 40083 5120 40693 5148
rect 40083 5117 40095 5120
rect 40037 5111 40095 5117
rect 40681 5117 40693 5120
rect 40727 5117 40739 5151
rect 40972 5148 41000 5256
rect 41322 5176 41328 5228
rect 41380 5216 41386 5228
rect 42337 5219 42395 5225
rect 42337 5216 42349 5219
rect 41380 5188 42349 5216
rect 41380 5176 41386 5188
rect 42337 5185 42349 5188
rect 42383 5185 42395 5219
rect 42337 5179 42395 5185
rect 43993 5219 44051 5225
rect 43993 5185 44005 5219
rect 44039 5216 44051 5219
rect 44174 5216 44180 5228
rect 44039 5188 44180 5216
rect 44039 5185 44051 5188
rect 43993 5179 44051 5185
rect 44174 5176 44180 5188
rect 44232 5176 44238 5228
rect 45465 5219 45523 5225
rect 45465 5185 45477 5219
rect 45511 5216 45523 5219
rect 46750 5216 46756 5228
rect 45511 5188 46756 5216
rect 45511 5185 45523 5188
rect 45465 5179 45523 5185
rect 46750 5176 46756 5188
rect 46808 5176 46814 5228
rect 47026 5176 47032 5228
rect 47084 5176 47090 5228
rect 41601 5151 41659 5157
rect 41601 5148 41613 5151
rect 40972 5120 41613 5148
rect 40681 5111 40739 5117
rect 41601 5117 41613 5120
rect 41647 5117 41659 5151
rect 41601 5111 41659 5117
rect 39316 5080 39344 5111
rect 41690 5108 41696 5160
rect 41748 5148 41754 5160
rect 42889 5151 42947 5157
rect 42889 5148 42901 5151
rect 41748 5120 42901 5148
rect 41748 5108 41754 5120
rect 42889 5117 42901 5120
rect 42935 5117 42947 5151
rect 42889 5111 42947 5117
rect 44085 5151 44143 5157
rect 44085 5117 44097 5151
rect 44131 5117 44143 5151
rect 44085 5111 44143 5117
rect 40129 5083 40187 5089
rect 40129 5080 40141 5083
rect 39316 5052 40141 5080
rect 40129 5049 40141 5052
rect 40175 5049 40187 5083
rect 40129 5043 40187 5049
rect 42702 5040 42708 5092
rect 42760 5080 42766 5092
rect 44100 5080 44128 5111
rect 45554 5108 45560 5160
rect 45612 5108 45618 5160
rect 46934 5108 46940 5160
rect 46992 5108 46998 5160
rect 76926 5108 76932 5160
rect 76984 5148 76990 5160
rect 77481 5151 77539 5157
rect 77481 5148 77493 5151
rect 76984 5120 77493 5148
rect 76984 5108 76990 5120
rect 77481 5117 77493 5120
rect 77527 5117 77539 5151
rect 77481 5111 77539 5117
rect 42760 5052 44128 5080
rect 42760 5040 42766 5052
rect 44818 5040 44824 5092
rect 44876 5040 44882 5092
rect 46201 5083 46259 5089
rect 46201 5049 46213 5083
rect 46247 5080 46259 5083
rect 47946 5080 47952 5092
rect 46247 5052 47952 5080
rect 46247 5049 46259 5052
rect 46201 5043 46259 5049
rect 47946 5040 47952 5052
rect 48004 5040 48010 5092
rect 42058 5012 42064 5024
rect 39224 4984 42064 5012
rect 42058 4972 42064 4984
rect 42116 4972 42122 5024
rect 42245 5015 42303 5021
rect 42245 4981 42257 5015
rect 42291 5012 42303 5015
rect 43254 5012 43260 5024
rect 42291 4984 43260 5012
rect 42291 4981 42303 4984
rect 42245 4975 42303 4981
rect 43254 4972 43260 4984
rect 43312 4972 43318 5024
rect 43346 4972 43352 5024
rect 43404 4972 43410 5024
rect 44729 5015 44787 5021
rect 44729 4981 44741 5015
rect 44775 5012 44787 5015
rect 45738 5012 45744 5024
rect 44775 4984 45744 5012
rect 44775 4981 44787 4984
rect 44729 4975 44787 4981
rect 45738 4972 45744 4984
rect 45796 4972 45802 5024
rect 46293 5015 46351 5021
rect 46293 4981 46305 5015
rect 46339 5012 46351 5015
rect 47210 5012 47216 5024
rect 46339 4984 47216 5012
rect 46339 4981 46351 4984
rect 46293 4975 46351 4981
rect 47210 4972 47216 4984
rect 47268 4972 47274 5024
rect 47673 5015 47731 5021
rect 47673 4981 47685 5015
rect 47719 5012 47731 5015
rect 49602 5012 49608 5024
rect 47719 4984 49608 5012
rect 47719 4981 47731 4984
rect 47673 4975 47731 4981
rect 49602 4972 49608 4984
rect 49660 4972 49666 5024
rect 76650 4972 76656 5024
rect 76708 5012 76714 5024
rect 76929 5015 76987 5021
rect 76929 5012 76941 5015
rect 76708 4984 76941 5012
rect 76708 4972 76714 4984
rect 76929 4981 76941 4984
rect 76975 4981 76987 5015
rect 76929 4975 76987 4981
rect 2024 4922 77924 4944
rect 2024 4870 5134 4922
rect 5186 4870 5198 4922
rect 5250 4870 5262 4922
rect 5314 4870 5326 4922
rect 5378 4870 5390 4922
rect 5442 4870 35854 4922
rect 35906 4870 35918 4922
rect 35970 4870 35982 4922
rect 36034 4870 36046 4922
rect 36098 4870 36110 4922
rect 36162 4870 66574 4922
rect 66626 4870 66638 4922
rect 66690 4870 66702 4922
rect 66754 4870 66766 4922
rect 66818 4870 66830 4922
rect 66882 4870 77924 4922
rect 2024 4848 77924 4870
rect 8941 4811 8999 4817
rect 8941 4777 8953 4811
rect 8987 4808 8999 4811
rect 9766 4808 9772 4820
rect 8987 4780 9772 4808
rect 8987 4777 8999 4780
rect 8941 4771 8999 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10229 4811 10287 4817
rect 10229 4777 10241 4811
rect 10275 4808 10287 4811
rect 11238 4808 11244 4820
rect 10275 4780 11244 4808
rect 10275 4777 10287 4780
rect 10229 4771 10287 4777
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 11885 4811 11943 4817
rect 11885 4777 11897 4811
rect 11931 4808 11943 4811
rect 15746 4808 15752 4820
rect 11931 4780 15752 4808
rect 11931 4777 11943 4780
rect 11885 4771 11943 4777
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 16114 4768 16120 4820
rect 16172 4808 16178 4820
rect 16485 4811 16543 4817
rect 16485 4808 16497 4811
rect 16172 4780 16497 4808
rect 16172 4768 16178 4780
rect 16485 4777 16497 4780
rect 16531 4777 16543 4811
rect 16485 4771 16543 4777
rect 19058 4768 19064 4820
rect 19116 4768 19122 4820
rect 19426 4768 19432 4820
rect 19484 4808 19490 4820
rect 21450 4808 21456 4820
rect 19484 4780 21456 4808
rect 19484 4768 19490 4780
rect 21450 4768 21456 4780
rect 21508 4768 21514 4820
rect 23198 4768 23204 4820
rect 23256 4808 23262 4820
rect 23385 4811 23443 4817
rect 23385 4808 23397 4811
rect 23256 4780 23397 4808
rect 23256 4768 23262 4780
rect 23385 4777 23397 4780
rect 23431 4777 23443 4811
rect 23385 4771 23443 4777
rect 24305 4811 24363 4817
rect 24305 4777 24317 4811
rect 24351 4808 24363 4811
rect 24486 4808 24492 4820
rect 24351 4780 24492 4808
rect 24351 4777 24363 4780
rect 24305 4771 24363 4777
rect 24486 4768 24492 4780
rect 24544 4768 24550 4820
rect 27893 4811 27951 4817
rect 27893 4777 27905 4811
rect 27939 4808 27951 4811
rect 27982 4808 27988 4820
rect 27939 4780 27988 4808
rect 27939 4777 27951 4780
rect 27893 4771 27951 4777
rect 27982 4768 27988 4780
rect 28040 4768 28046 4820
rect 29638 4768 29644 4820
rect 29696 4768 29702 4820
rect 30190 4768 30196 4820
rect 30248 4808 30254 4820
rect 30558 4808 30564 4820
rect 30248 4780 30564 4808
rect 30248 4768 30254 4780
rect 30558 4768 30564 4780
rect 30616 4768 30622 4820
rect 31202 4768 31208 4820
rect 31260 4808 31266 4820
rect 31389 4811 31447 4817
rect 31389 4808 31401 4811
rect 31260 4780 31401 4808
rect 31260 4768 31266 4780
rect 31389 4777 31401 4780
rect 31435 4777 31447 4811
rect 31389 4771 31447 4777
rect 32677 4811 32735 4817
rect 32677 4777 32689 4811
rect 32723 4808 32735 4811
rect 32766 4808 32772 4820
rect 32723 4780 32772 4808
rect 32723 4777 32735 4780
rect 32677 4771 32735 4777
rect 32766 4768 32772 4780
rect 32824 4768 32830 4820
rect 32858 4768 32864 4820
rect 32916 4768 32922 4820
rect 33321 4811 33379 4817
rect 33321 4777 33333 4811
rect 33367 4808 33379 4811
rect 33686 4808 33692 4820
rect 33367 4780 33692 4808
rect 33367 4777 33379 4780
rect 33321 4771 33379 4777
rect 33686 4768 33692 4780
rect 33744 4768 33750 4820
rect 36262 4768 36268 4820
rect 36320 4808 36326 4820
rect 37093 4811 37151 4817
rect 37093 4808 37105 4811
rect 36320 4780 37105 4808
rect 36320 4768 36326 4780
rect 37093 4777 37105 4780
rect 37139 4777 37151 4811
rect 37093 4771 37151 4777
rect 37274 4768 37280 4820
rect 37332 4808 37338 4820
rect 41417 4811 41475 4817
rect 37332 4780 40356 4808
rect 37332 4768 37338 4780
rect 9677 4743 9735 4749
rect 9677 4709 9689 4743
rect 9723 4740 9735 4743
rect 11054 4740 11060 4752
rect 9723 4712 11060 4740
rect 9723 4709 9735 4712
rect 9677 4703 9735 4709
rect 11054 4700 11060 4712
rect 11112 4700 11118 4752
rect 12342 4700 12348 4752
rect 12400 4740 12406 4752
rect 12400 4700 12434 4740
rect 12618 4700 12624 4752
rect 12676 4700 12682 4752
rect 14093 4743 14151 4749
rect 14093 4709 14105 4743
rect 14139 4740 14151 4743
rect 16758 4740 16764 4752
rect 14139 4712 16764 4740
rect 14139 4709 14151 4712
rect 14093 4703 14151 4709
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 17221 4743 17279 4749
rect 17221 4709 17233 4743
rect 17267 4740 17279 4743
rect 19518 4740 19524 4752
rect 17267 4712 19012 4740
rect 17267 4709 17279 4712
rect 17221 4703 17279 4709
rect 8294 4632 8300 4684
rect 8352 4632 8358 4684
rect 12406 4672 12434 4700
rect 13357 4675 13415 4681
rect 13357 4672 13369 4675
rect 9048 4644 12296 4672
rect 12406 4644 13369 4672
rect 6730 4564 6736 4616
rect 6788 4564 6794 4616
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4604 7711 4607
rect 9048 4604 9076 4644
rect 7699 4576 9076 4604
rect 7699 4573 7711 4576
rect 7653 4567 7711 4573
rect 7484 4536 7512 4567
rect 9122 4564 9128 4616
rect 9180 4564 9186 4616
rect 10594 4564 10600 4616
rect 10652 4564 10658 4616
rect 11149 4607 11207 4613
rect 11149 4573 11161 4607
rect 11195 4604 11207 4607
rect 11330 4604 11336 4616
rect 11195 4576 11336 4604
rect 11195 4573 11207 4576
rect 11149 4567 11207 4573
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 11974 4564 11980 4616
rect 12032 4564 12038 4616
rect 12268 4604 12296 4644
rect 13357 4641 13369 4644
rect 13403 4641 13415 4675
rect 13357 4635 13415 4641
rect 13538 4632 13544 4684
rect 13596 4632 13602 4684
rect 14274 4632 14280 4684
rect 14332 4672 14338 4684
rect 15841 4675 15899 4681
rect 15841 4672 15853 4675
rect 14332 4644 15853 4672
rect 14332 4632 14338 4644
rect 15841 4641 15853 4644
rect 15887 4641 15899 4675
rect 15841 4635 15899 4641
rect 16206 4632 16212 4684
rect 16264 4672 16270 4684
rect 16577 4675 16635 4681
rect 16577 4672 16589 4675
rect 16264 4644 16589 4672
rect 16264 4632 16270 4644
rect 16577 4641 16589 4644
rect 16623 4641 16635 4675
rect 17126 4672 17132 4684
rect 16577 4635 16635 4641
rect 16684 4644 17132 4672
rect 12342 4604 12348 4616
rect 12268 4576 12348 4604
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 12802 4564 12808 4616
rect 12860 4564 12866 4616
rect 14185 4607 14243 4613
rect 14185 4573 14197 4607
rect 14231 4604 14243 4607
rect 15010 4604 15016 4616
rect 14231 4576 15016 4604
rect 14231 4573 14243 4576
rect 14185 4567 14243 4573
rect 15010 4564 15016 4576
rect 15068 4564 15074 4616
rect 15105 4607 15163 4613
rect 15105 4573 15117 4607
rect 15151 4604 15163 4607
rect 16684 4604 16712 4644
rect 17126 4632 17132 4644
rect 17184 4632 17190 4684
rect 18984 4672 19012 4712
rect 19168 4712 19524 4740
rect 19168 4672 19196 4712
rect 19518 4700 19524 4712
rect 19576 4700 19582 4752
rect 19886 4740 19892 4752
rect 19720 4712 19892 4740
rect 19720 4681 19748 4712
rect 19886 4700 19892 4712
rect 19944 4740 19950 4752
rect 21726 4740 21732 4752
rect 19944 4712 21732 4740
rect 19944 4700 19950 4712
rect 21726 4700 21732 4712
rect 21784 4700 21790 4752
rect 21818 4700 21824 4752
rect 21876 4700 21882 4752
rect 26237 4743 26295 4749
rect 22480 4712 26188 4740
rect 19705 4675 19763 4681
rect 18984 4644 19196 4672
rect 19352 4644 19656 4672
rect 15151 4576 16712 4604
rect 17405 4607 17463 4613
rect 15151 4573 15163 4576
rect 15105 4567 15163 4573
rect 17405 4573 17417 4607
rect 17451 4604 17463 4607
rect 17451 4576 17540 4604
rect 17451 4573 17463 4576
rect 17405 4567 17463 4573
rect 9766 4536 9772 4548
rect 7484 4508 9772 4536
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 10321 4539 10379 4545
rect 10321 4505 10333 4539
rect 10367 4536 10379 4539
rect 12710 4536 12716 4548
rect 10367 4508 12716 4536
rect 10367 4505 10379 4508
rect 10321 4499 10379 4505
rect 12710 4496 12716 4508
rect 12768 4496 12774 4548
rect 15749 4539 15807 4545
rect 15749 4505 15761 4539
rect 15795 4536 15807 4539
rect 15838 4536 15844 4548
rect 15795 4508 15844 4536
rect 15795 4505 15807 4508
rect 15749 4499 15807 4505
rect 15838 4496 15844 4508
rect 15896 4496 15902 4548
rect 17512 4536 17540 4576
rect 17586 4564 17592 4616
rect 17644 4604 17650 4616
rect 19352 4604 19380 4644
rect 17644 4576 19380 4604
rect 19628 4604 19656 4644
rect 19705 4641 19717 4675
rect 19751 4641 19763 4675
rect 19705 4635 19763 4641
rect 20533 4675 20591 4681
rect 20533 4641 20545 4675
rect 20579 4672 20591 4675
rect 20622 4672 20628 4684
rect 20579 4644 20628 4672
rect 20579 4641 20591 4644
rect 20533 4635 20591 4641
rect 20622 4632 20628 4644
rect 20680 4632 20686 4684
rect 21085 4675 21143 4681
rect 21085 4641 21097 4675
rect 21131 4672 21143 4675
rect 22480 4672 22508 4712
rect 21131 4644 22508 4672
rect 22557 4675 22615 4681
rect 21131 4641 21143 4644
rect 21085 4635 21143 4641
rect 22557 4641 22569 4675
rect 22603 4672 22615 4675
rect 23566 4672 23572 4684
rect 22603 4644 23572 4672
rect 22603 4641 22615 4644
rect 22557 4635 22615 4641
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 23937 4675 23995 4681
rect 23937 4641 23949 4675
rect 23983 4672 23995 4675
rect 24302 4672 24308 4684
rect 23983 4644 24308 4672
rect 23983 4641 23995 4644
rect 23937 4635 23995 4641
rect 24302 4632 24308 4644
rect 24360 4632 24366 4684
rect 24762 4632 24768 4684
rect 24820 4632 24826 4684
rect 24949 4675 25007 4681
rect 24949 4641 24961 4675
rect 24995 4672 25007 4675
rect 25038 4672 25044 4684
rect 24995 4644 25044 4672
rect 24995 4641 25007 4644
rect 24949 4635 25007 4641
rect 25038 4632 25044 4644
rect 25096 4632 25102 4684
rect 26160 4672 26188 4712
rect 26237 4709 26249 4743
rect 26283 4740 26295 4743
rect 32490 4740 32496 4752
rect 26283 4712 32496 4740
rect 26283 4709 26295 4712
rect 26237 4703 26295 4709
rect 32490 4700 32496 4712
rect 32548 4700 32554 4752
rect 36814 4740 36820 4752
rect 32600 4712 36820 4740
rect 26326 4672 26332 4684
rect 26160 4644 26332 4672
rect 26326 4632 26332 4644
rect 26384 4632 26390 4684
rect 26418 4632 26424 4684
rect 26476 4632 26482 4684
rect 26878 4632 26884 4684
rect 26936 4672 26942 4684
rect 26936 4644 27660 4672
rect 26936 4632 26942 4644
rect 20898 4604 20904 4616
rect 19628 4576 20904 4604
rect 17644 4564 17650 4576
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 21269 4607 21327 4613
rect 21269 4573 21281 4607
rect 21315 4604 21327 4607
rect 21542 4604 21548 4616
rect 21315 4576 21548 4604
rect 21315 4573 21327 4576
rect 21269 4567 21327 4573
rect 21542 4564 21548 4576
rect 21600 4564 21606 4616
rect 21910 4564 21916 4616
rect 21968 4564 21974 4616
rect 22646 4564 22652 4616
rect 22704 4564 22710 4616
rect 23014 4564 23020 4616
rect 23072 4604 23078 4616
rect 23382 4604 23388 4616
rect 23072 4576 23388 4604
rect 23072 4564 23078 4576
rect 23382 4564 23388 4576
rect 23440 4604 23446 4616
rect 23753 4607 23811 4613
rect 23753 4604 23765 4607
rect 23440 4576 23765 4604
rect 23440 4564 23446 4576
rect 23753 4573 23765 4576
rect 23799 4573 23811 4607
rect 23753 4567 23811 4573
rect 23845 4607 23903 4613
rect 23845 4573 23857 4607
rect 23891 4604 23903 4607
rect 24026 4604 24032 4616
rect 23891 4576 24032 4604
rect 23891 4573 23903 4576
rect 23845 4567 23903 4573
rect 24026 4564 24032 4576
rect 24084 4564 24090 4616
rect 24670 4564 24676 4616
rect 24728 4564 24734 4616
rect 25685 4607 25743 4613
rect 25685 4573 25697 4607
rect 25731 4604 25743 4607
rect 27430 4604 27436 4616
rect 25731 4576 27436 4604
rect 25731 4573 25743 4576
rect 25685 4567 25743 4573
rect 27430 4564 27436 4576
rect 27488 4564 27494 4616
rect 17862 4536 17868 4548
rect 17512 4508 17868 4536
rect 17862 4496 17868 4508
rect 17920 4496 17926 4548
rect 18046 4496 18052 4548
rect 18104 4496 18110 4548
rect 19429 4539 19487 4545
rect 19429 4505 19441 4539
rect 19475 4505 19487 4539
rect 19429 4499 19487 4505
rect 19521 4539 19579 4545
rect 19521 4505 19533 4539
rect 19567 4536 19579 4539
rect 20162 4536 20168 4548
rect 19567 4508 20168 4536
rect 19567 4505 19579 4508
rect 19521 4499 19579 4505
rect 6089 4471 6147 4477
rect 6089 4437 6101 4471
rect 6135 4468 6147 4471
rect 6454 4468 6460 4480
rect 6135 4440 6460 4468
rect 6135 4437 6147 4440
rect 6089 4431 6147 4437
rect 6454 4428 6460 4440
rect 6512 4428 6518 4480
rect 6822 4428 6828 4480
rect 6880 4428 6886 4480
rect 8205 4471 8263 4477
rect 8205 4437 8217 4471
rect 8251 4468 8263 4471
rect 9582 4468 9588 4480
rect 8251 4440 9588 4468
rect 8251 4437 8263 4440
rect 8205 4431 8263 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 12894 4468 12900 4480
rect 12492 4440 12900 4468
rect 12492 4428 12498 4440
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 14829 4471 14887 4477
rect 14829 4437 14841 4471
rect 14875 4468 14887 4471
rect 15654 4468 15660 4480
rect 14875 4440 15660 4468
rect 14875 4437 14887 4440
rect 14829 4431 14887 4437
rect 15654 4428 15660 4440
rect 15712 4428 15718 4480
rect 17957 4471 18015 4477
rect 17957 4437 17969 4471
rect 18003 4468 18015 4471
rect 18322 4468 18328 4480
rect 18003 4440 18328 4468
rect 18003 4437 18015 4440
rect 17957 4431 18015 4437
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 18414 4428 18420 4480
rect 18472 4468 18478 4480
rect 19444 4468 19472 4499
rect 20162 4496 20168 4508
rect 20220 4496 20226 4548
rect 22572 4508 24900 4536
rect 18472 4440 19472 4468
rect 18472 4428 18478 4440
rect 19610 4428 19616 4480
rect 19668 4468 19674 4480
rect 19886 4468 19892 4480
rect 19668 4440 19892 4468
rect 19668 4428 19674 4440
rect 19886 4428 19892 4440
rect 19944 4428 19950 4480
rect 22278 4428 22284 4480
rect 22336 4468 22342 4480
rect 22572 4468 22600 4508
rect 22336 4440 22600 4468
rect 23293 4471 23351 4477
rect 22336 4428 22342 4440
rect 23293 4437 23305 4471
rect 23339 4468 23351 4471
rect 24762 4468 24768 4480
rect 23339 4440 24768 4468
rect 23339 4437 23351 4440
rect 23293 4431 23351 4437
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 24872 4468 24900 4508
rect 24946 4496 24952 4548
rect 25004 4536 25010 4548
rect 26234 4536 26240 4548
rect 25004 4508 26240 4536
rect 25004 4496 25010 4508
rect 26234 4496 26240 4508
rect 26292 4496 26298 4548
rect 26973 4539 27031 4545
rect 26973 4505 26985 4539
rect 27019 4536 27031 4539
rect 27522 4536 27528 4548
rect 27019 4508 27528 4536
rect 27019 4505 27031 4508
rect 26973 4499 27031 4505
rect 27522 4496 27528 4508
rect 27580 4496 27586 4548
rect 27632 4536 27660 4644
rect 28166 4632 28172 4684
rect 28224 4672 28230 4684
rect 28353 4675 28411 4681
rect 28353 4672 28365 4675
rect 28224 4644 28365 4672
rect 28224 4632 28230 4644
rect 28353 4641 28365 4644
rect 28399 4641 28411 4675
rect 28353 4635 28411 4641
rect 28445 4675 28503 4681
rect 28445 4641 28457 4675
rect 28491 4641 28503 4675
rect 28445 4635 28503 4641
rect 27709 4607 27767 4613
rect 27709 4573 27721 4607
rect 27755 4604 27767 4607
rect 27982 4604 27988 4616
rect 27755 4576 27988 4604
rect 27755 4573 27767 4576
rect 27709 4567 27767 4573
rect 27982 4564 27988 4576
rect 28040 4564 28046 4616
rect 28258 4564 28264 4616
rect 28316 4604 28322 4616
rect 28460 4604 28488 4635
rect 28902 4632 28908 4684
rect 28960 4632 28966 4684
rect 30466 4672 30472 4684
rect 29196 4644 30472 4672
rect 28316 4576 28488 4604
rect 28316 4564 28322 4576
rect 29196 4536 29224 4644
rect 30466 4632 30472 4644
rect 30524 4632 30530 4684
rect 30742 4632 30748 4684
rect 30800 4632 30806 4684
rect 31202 4632 31208 4684
rect 31260 4672 31266 4684
rect 31570 4672 31576 4684
rect 31260 4644 31576 4672
rect 31260 4632 31266 4644
rect 31570 4632 31576 4644
rect 31628 4632 31634 4684
rect 31846 4632 31852 4684
rect 31904 4632 31910 4684
rect 31938 4632 31944 4684
rect 31996 4632 32002 4684
rect 32600 4681 32628 4712
rect 36814 4700 36820 4712
rect 36872 4700 36878 4752
rect 37001 4743 37059 4749
rect 37001 4709 37013 4743
rect 37047 4740 37059 4743
rect 37458 4740 37464 4752
rect 37047 4712 37464 4740
rect 37047 4709 37059 4712
rect 37001 4703 37059 4709
rect 37458 4700 37464 4712
rect 37516 4700 37522 4752
rect 32585 4675 32643 4681
rect 32585 4641 32597 4675
rect 32631 4641 32643 4675
rect 32585 4635 32643 4641
rect 32858 4632 32864 4684
rect 32916 4672 32922 4684
rect 33042 4672 33048 4684
rect 32916 4644 33048 4672
rect 32916 4632 32922 4644
rect 33042 4632 33048 4644
rect 33100 4632 33106 4684
rect 33226 4632 33232 4684
rect 33284 4672 33290 4684
rect 35621 4675 35679 4681
rect 35621 4672 35633 4675
rect 33284 4644 35633 4672
rect 33284 4632 33290 4644
rect 35621 4641 35633 4644
rect 35667 4641 35679 4675
rect 35621 4635 35679 4641
rect 36449 4675 36507 4681
rect 36449 4641 36461 4675
rect 36495 4672 36507 4675
rect 37366 4672 37372 4684
rect 36495 4644 37372 4672
rect 36495 4641 36507 4644
rect 36449 4635 36507 4641
rect 37366 4632 37372 4644
rect 37424 4632 37430 4684
rect 37734 4632 37740 4684
rect 37792 4632 37798 4684
rect 37826 4632 37832 4684
rect 37884 4672 37890 4684
rect 38197 4675 38255 4681
rect 38197 4672 38209 4675
rect 37884 4644 38209 4672
rect 37884 4632 37890 4644
rect 38197 4641 38209 4644
rect 38243 4641 38255 4675
rect 38197 4635 38255 4641
rect 38930 4632 38936 4684
rect 38988 4672 38994 4684
rect 38988 4644 40264 4672
rect 38988 4632 38994 4644
rect 29362 4564 29368 4616
rect 29420 4604 29426 4616
rect 29914 4604 29920 4616
rect 29420 4576 29920 4604
rect 29420 4564 29426 4576
rect 29914 4564 29920 4576
rect 29972 4564 29978 4616
rect 30282 4564 30288 4616
rect 30340 4564 30346 4616
rect 32677 4607 32735 4613
rect 30392 4576 32168 4604
rect 27632 4508 29224 4536
rect 29270 4496 29276 4548
rect 29328 4536 29334 4548
rect 30392 4536 30420 4576
rect 29328 4508 30420 4536
rect 29328 4496 29334 4508
rect 30742 4496 30748 4548
rect 30800 4536 30806 4548
rect 31297 4539 31355 4545
rect 31297 4536 31309 4539
rect 30800 4508 31309 4536
rect 30800 4496 30806 4508
rect 31297 4505 31309 4508
rect 31343 4505 31355 4539
rect 31297 4499 31355 4505
rect 31754 4496 31760 4548
rect 31812 4496 31818 4548
rect 32140 4536 32168 4576
rect 32677 4573 32689 4607
rect 32723 4604 32735 4607
rect 33318 4604 33324 4616
rect 32723 4576 33324 4604
rect 32723 4573 32735 4576
rect 32677 4567 32735 4573
rect 33318 4564 33324 4576
rect 33376 4564 33382 4616
rect 33965 4607 34023 4613
rect 33965 4573 33977 4607
rect 34011 4573 34023 4607
rect 33965 4567 34023 4573
rect 34149 4607 34207 4613
rect 34149 4573 34161 4607
rect 34195 4604 34207 4607
rect 34606 4604 34612 4616
rect 34195 4576 34612 4604
rect 34195 4573 34207 4576
rect 34149 4567 34207 4573
rect 32217 4539 32275 4545
rect 32217 4536 32229 4539
rect 32140 4508 32229 4536
rect 32217 4505 32229 4508
rect 32263 4505 32275 4539
rect 32217 4499 32275 4505
rect 27065 4471 27123 4477
rect 27065 4468 27077 4471
rect 24872 4440 27077 4468
rect 27065 4437 27077 4440
rect 27111 4437 27123 4471
rect 27065 4431 27123 4437
rect 27614 4428 27620 4480
rect 27672 4468 27678 4480
rect 28261 4471 28319 4477
rect 28261 4468 28273 4471
rect 27672 4440 28273 4468
rect 27672 4428 27678 4440
rect 28261 4437 28273 4440
rect 28307 4468 28319 4471
rect 28442 4468 28448 4480
rect 28307 4440 28448 4468
rect 28307 4437 28319 4440
rect 28261 4431 28319 4437
rect 28442 4428 28448 4440
rect 28500 4428 28506 4480
rect 29546 4428 29552 4480
rect 29604 4428 29610 4480
rect 30466 4428 30472 4480
rect 30524 4468 30530 4480
rect 31662 4468 31668 4480
rect 30524 4440 31668 4468
rect 30524 4428 30530 4440
rect 31662 4428 31668 4440
rect 31720 4428 31726 4480
rect 32232 4468 32260 4499
rect 32582 4496 32588 4548
rect 32640 4536 32646 4548
rect 32953 4539 33011 4545
rect 32953 4536 32965 4539
rect 32640 4508 32965 4536
rect 32640 4496 32646 4508
rect 32953 4505 32965 4508
rect 32999 4505 33011 4539
rect 32953 4499 33011 4505
rect 33134 4496 33140 4548
rect 33192 4496 33198 4548
rect 33980 4536 34008 4567
rect 34606 4564 34612 4576
rect 34664 4564 34670 4616
rect 34885 4607 34943 4613
rect 34885 4573 34897 4607
rect 34931 4604 34943 4607
rect 35250 4604 35256 4616
rect 34931 4576 35256 4604
rect 34931 4573 34943 4576
rect 34885 4567 34943 4573
rect 35250 4564 35256 4576
rect 35308 4564 35314 4616
rect 35360 4576 37688 4604
rect 34701 4539 34759 4545
rect 33980 4508 34652 4536
rect 34514 4468 34520 4480
rect 32232 4440 34520 4468
rect 34514 4428 34520 4440
rect 34572 4428 34578 4480
rect 34624 4468 34652 4508
rect 34701 4505 34713 4539
rect 34747 4536 34759 4539
rect 35360 4536 35388 4576
rect 34747 4508 35388 4536
rect 35437 4539 35495 4545
rect 34747 4505 34759 4508
rect 34701 4499 34759 4505
rect 35437 4505 35449 4539
rect 35483 4536 35495 4539
rect 35483 4508 36492 4536
rect 35483 4505 35495 4508
rect 35437 4499 35495 4505
rect 36078 4468 36084 4480
rect 34624 4440 36084 4468
rect 36078 4428 36084 4440
rect 36136 4428 36142 4480
rect 36262 4428 36268 4480
rect 36320 4428 36326 4480
rect 36464 4468 36492 4508
rect 37461 4471 37519 4477
rect 37461 4468 37473 4471
rect 36464 4440 37473 4468
rect 37461 4437 37473 4440
rect 37507 4437 37519 4471
rect 37461 4431 37519 4437
rect 37550 4428 37556 4480
rect 37608 4428 37614 4480
rect 37660 4468 37688 4576
rect 37918 4564 37924 4616
rect 37976 4564 37982 4616
rect 40236 4613 40264 4644
rect 40328 4613 40356 4780
rect 41417 4777 41429 4811
rect 41463 4808 41475 4811
rect 41690 4808 41696 4820
rect 41463 4780 41696 4808
rect 41463 4777 41475 4780
rect 41417 4771 41475 4777
rect 41690 4768 41696 4780
rect 41748 4768 41754 4820
rect 42058 4768 42064 4820
rect 42116 4808 42122 4820
rect 42797 4811 42855 4817
rect 42797 4808 42809 4811
rect 42116 4780 42809 4808
rect 42116 4768 42122 4780
rect 42797 4777 42809 4780
rect 42843 4777 42855 4811
rect 42797 4771 42855 4777
rect 42886 4768 42892 4820
rect 42944 4808 42950 4820
rect 43533 4811 43591 4817
rect 43533 4808 43545 4811
rect 42944 4780 43545 4808
rect 42944 4768 42950 4780
rect 43533 4777 43545 4780
rect 43579 4777 43591 4811
rect 43533 4771 43591 4777
rect 43622 4768 43628 4820
rect 43680 4808 43686 4820
rect 45005 4811 45063 4817
rect 45005 4808 45017 4811
rect 43680 4780 45017 4808
rect 43680 4768 43686 4780
rect 45005 4777 45017 4780
rect 45051 4777 45063 4811
rect 45005 4771 45063 4777
rect 45830 4768 45836 4820
rect 45888 4808 45894 4820
rect 46661 4811 46719 4817
rect 46661 4808 46673 4811
rect 45888 4780 46673 4808
rect 45888 4768 45894 4780
rect 46661 4777 46673 4780
rect 46707 4777 46719 4811
rect 46661 4771 46719 4777
rect 76926 4768 76932 4820
rect 76984 4768 76990 4820
rect 44269 4743 44327 4749
rect 44269 4740 44281 4743
rect 41386 4712 44281 4740
rect 40865 4675 40923 4681
rect 40865 4641 40877 4675
rect 40911 4672 40923 4675
rect 41386 4672 41414 4712
rect 44269 4709 44281 4712
rect 44315 4709 44327 4743
rect 44269 4703 44327 4709
rect 40911 4644 41414 4672
rect 40911 4641 40923 4644
rect 40865 4635 40923 4641
rect 43254 4632 43260 4684
rect 43312 4672 43318 4684
rect 44821 4675 44879 4681
rect 44821 4672 44833 4675
rect 43312 4644 44833 4672
rect 43312 4632 43318 4644
rect 44821 4641 44833 4644
rect 44867 4641 44879 4675
rect 44821 4635 44879 4641
rect 45462 4632 45468 4684
rect 45520 4672 45526 4684
rect 45925 4675 45983 4681
rect 45925 4672 45937 4675
rect 45520 4644 45937 4672
rect 45520 4632 45526 4644
rect 45925 4641 45937 4644
rect 45971 4641 45983 4675
rect 45925 4635 45983 4641
rect 47210 4632 47216 4684
rect 47268 4632 47274 4684
rect 48314 4632 48320 4684
rect 48372 4672 48378 4684
rect 48869 4675 48927 4681
rect 48869 4672 48881 4675
rect 48372 4644 48881 4672
rect 48372 4632 48378 4644
rect 48869 4641 48881 4644
rect 48915 4641 48927 4675
rect 48869 4635 48927 4641
rect 40221 4607 40279 4613
rect 40221 4573 40233 4607
rect 40267 4573 40279 4607
rect 40221 4567 40279 4573
rect 40313 4607 40371 4613
rect 40313 4573 40325 4607
rect 40359 4573 40371 4607
rect 40313 4567 40371 4573
rect 40494 4564 40500 4616
rect 40552 4604 40558 4616
rect 40589 4607 40647 4613
rect 40589 4604 40601 4607
rect 40552 4576 40601 4604
rect 40552 4564 40558 4576
rect 40589 4573 40601 4576
rect 40635 4573 40647 4607
rect 40589 4567 40647 4573
rect 41138 4564 41144 4616
rect 41196 4604 41202 4616
rect 42245 4607 42303 4613
rect 42245 4604 42257 4607
rect 41196 4576 42257 4604
rect 41196 4564 41202 4576
rect 42245 4573 42257 4576
rect 42291 4573 42303 4607
rect 42245 4567 42303 4573
rect 43441 4607 43499 4613
rect 43441 4573 43453 4607
rect 43487 4604 43499 4607
rect 43990 4604 43996 4616
rect 43487 4576 43996 4604
rect 43487 4573 43499 4576
rect 43441 4567 43499 4573
rect 43990 4564 43996 4576
rect 44048 4564 44054 4616
rect 44177 4607 44235 4613
rect 44177 4573 44189 4607
rect 44223 4604 44235 4607
rect 44223 4576 44312 4604
rect 44223 4573 44235 4576
rect 44177 4567 44235 4573
rect 39574 4536 39580 4548
rect 39422 4508 39580 4536
rect 39574 4496 39580 4508
rect 39632 4496 39638 4548
rect 39942 4496 39948 4548
rect 40000 4496 40006 4548
rect 40405 4539 40463 4545
rect 40405 4505 40417 4539
rect 40451 4536 40463 4539
rect 40770 4536 40776 4548
rect 40451 4508 40776 4536
rect 40451 4505 40463 4508
rect 40405 4499 40463 4505
rect 40770 4496 40776 4508
rect 40828 4496 40834 4548
rect 41046 4496 41052 4548
rect 41104 4536 41110 4548
rect 43622 4536 43628 4548
rect 41104 4508 43628 4536
rect 41104 4496 41110 4508
rect 43622 4496 43628 4508
rect 43680 4496 43686 4548
rect 38562 4468 38568 4480
rect 37660 4440 38568 4468
rect 38562 4428 38568 4440
rect 38620 4428 38626 4480
rect 39022 4428 39028 4480
rect 39080 4468 39086 4480
rect 40037 4471 40095 4477
rect 40037 4468 40049 4471
rect 39080 4440 40049 4468
rect 39080 4428 39086 4440
rect 40037 4437 40049 4440
rect 40083 4437 40095 4471
rect 40037 4431 40095 4437
rect 41690 4428 41696 4480
rect 41748 4428 41754 4480
rect 41874 4428 41880 4480
rect 41932 4468 41938 4480
rect 44284 4468 44312 4576
rect 45278 4564 45284 4616
rect 45336 4604 45342 4616
rect 45557 4607 45615 4613
rect 45557 4604 45569 4607
rect 45336 4576 45569 4604
rect 45336 4564 45342 4576
rect 45557 4573 45569 4576
rect 45603 4573 45615 4607
rect 45557 4567 45615 4573
rect 47397 4607 47455 4613
rect 47397 4573 47409 4607
rect 47443 4573 47455 4607
rect 47397 4567 47455 4573
rect 47412 4536 47440 4567
rect 48774 4564 48780 4616
rect 48832 4564 48838 4616
rect 77570 4564 77576 4616
rect 77628 4564 77634 4616
rect 45112 4508 47440 4536
rect 48041 4539 48099 4545
rect 41932 4440 44312 4468
rect 41932 4428 41938 4440
rect 44450 4428 44456 4480
rect 44508 4468 44514 4480
rect 45112 4468 45140 4508
rect 48041 4505 48053 4539
rect 48087 4536 48099 4539
rect 48498 4536 48504 4548
rect 48087 4508 48504 4536
rect 48087 4505 48099 4508
rect 48041 4499 48099 4505
rect 48498 4496 48504 4508
rect 48556 4496 48562 4548
rect 44508 4440 45140 4468
rect 46569 4471 46627 4477
rect 44508 4428 44514 4440
rect 46569 4437 46581 4471
rect 46615 4468 46627 4471
rect 47854 4468 47860 4480
rect 46615 4440 47860 4468
rect 46615 4437 46627 4440
rect 46569 4431 46627 4437
rect 47854 4428 47860 4440
rect 47912 4428 47918 4480
rect 48133 4471 48191 4477
rect 48133 4437 48145 4471
rect 48179 4468 48191 4471
rect 48406 4468 48412 4480
rect 48179 4440 48412 4468
rect 48179 4437 48191 4440
rect 48133 4431 48191 4437
rect 48406 4428 48412 4440
rect 48464 4428 48470 4480
rect 49513 4471 49571 4477
rect 49513 4437 49525 4471
rect 49559 4468 49571 4471
rect 49694 4468 49700 4480
rect 49559 4440 49700 4468
rect 49559 4437 49571 4440
rect 49513 4431 49571 4437
rect 49694 4428 49700 4440
rect 49752 4428 49758 4480
rect 2024 4378 77924 4400
rect 2024 4326 5794 4378
rect 5846 4326 5858 4378
rect 5910 4326 5922 4378
rect 5974 4326 5986 4378
rect 6038 4326 6050 4378
rect 6102 4326 36514 4378
rect 36566 4326 36578 4378
rect 36630 4326 36642 4378
rect 36694 4326 36706 4378
rect 36758 4326 36770 4378
rect 36822 4326 67234 4378
rect 67286 4326 67298 4378
rect 67350 4326 67362 4378
rect 67414 4326 67426 4378
rect 67478 4326 67490 4378
rect 67542 4326 77924 4378
rect 2024 4304 77924 4326
rect 7101 4267 7159 4273
rect 7101 4233 7113 4267
rect 7147 4264 7159 4267
rect 7466 4264 7472 4276
rect 7147 4236 7472 4264
rect 7147 4233 7159 4236
rect 7101 4227 7159 4233
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 9122 4224 9128 4276
rect 9180 4264 9186 4276
rect 13998 4264 14004 4276
rect 9180 4236 14004 4264
rect 9180 4224 9186 4236
rect 13998 4224 14004 4236
rect 14056 4224 14062 4276
rect 17126 4224 17132 4276
rect 17184 4264 17190 4276
rect 17770 4264 17776 4276
rect 17184 4236 17776 4264
rect 17184 4224 17190 4236
rect 17770 4224 17776 4236
rect 17828 4264 17834 4276
rect 19978 4264 19984 4276
rect 17828 4236 19984 4264
rect 17828 4224 17834 4236
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 20073 4267 20131 4273
rect 20073 4233 20085 4267
rect 20119 4264 20131 4267
rect 20530 4264 20536 4276
rect 20119 4236 20536 4264
rect 20119 4233 20131 4236
rect 20073 4227 20131 4233
rect 20530 4224 20536 4236
rect 20588 4224 20594 4276
rect 20809 4267 20867 4273
rect 20809 4233 20821 4267
rect 20855 4264 20867 4267
rect 21910 4264 21916 4276
rect 20855 4236 21916 4264
rect 20855 4233 20867 4236
rect 20809 4227 20867 4233
rect 21910 4224 21916 4236
rect 21968 4224 21974 4276
rect 22462 4224 22468 4276
rect 22520 4264 22526 4276
rect 22899 4267 22957 4273
rect 22899 4264 22911 4267
rect 22520 4236 22911 4264
rect 22520 4224 22526 4236
rect 22899 4233 22911 4236
rect 22945 4233 22957 4267
rect 23198 4264 23204 4276
rect 22899 4227 22957 4233
rect 23124 4236 23204 4264
rect 8570 4196 8576 4208
rect 7668 4168 8576 4196
rect 6362 4088 6368 4140
rect 6420 4088 6426 4140
rect 6454 4088 6460 4140
rect 6512 4088 6518 4140
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4128 7619 4131
rect 7668 4128 7696 4168
rect 8570 4156 8576 4168
rect 8628 4156 8634 4208
rect 9766 4156 9772 4208
rect 9824 4196 9830 4208
rect 12434 4196 12440 4208
rect 9824 4168 12440 4196
rect 9824 4156 9830 4168
rect 12434 4156 12440 4168
rect 12492 4156 12498 4208
rect 12529 4199 12587 4205
rect 12529 4165 12541 4199
rect 12575 4196 12587 4199
rect 12802 4196 12808 4208
rect 12575 4168 12808 4196
rect 12575 4165 12587 4168
rect 12529 4159 12587 4165
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 13170 4156 13176 4208
rect 13228 4196 13234 4208
rect 13357 4199 13415 4205
rect 13357 4196 13369 4199
rect 13228 4168 13369 4196
rect 13228 4156 13234 4168
rect 13357 4165 13369 4168
rect 13403 4165 13415 4199
rect 13357 4159 13415 4165
rect 14826 4156 14832 4208
rect 14884 4196 14890 4208
rect 16298 4196 16304 4208
rect 14884 4168 16304 4196
rect 14884 4156 14890 4168
rect 16298 4156 16304 4168
rect 16356 4156 16362 4208
rect 16758 4156 16764 4208
rect 16816 4196 16822 4208
rect 17405 4199 17463 4205
rect 17405 4196 17417 4199
rect 16816 4168 17417 4196
rect 16816 4156 16822 4168
rect 17405 4165 17417 4168
rect 17451 4165 17463 4199
rect 19797 4199 19855 4205
rect 17405 4159 17463 4165
rect 17512 4168 19334 4196
rect 7607 4100 7696 4128
rect 7607 4097 7619 4100
rect 7561 4091 7619 4097
rect 7742 4088 7748 4140
rect 7800 4088 7806 4140
rect 7834 4088 7840 4140
rect 7892 4088 7898 4140
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8067 4100 9812 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 9784 4072 9812 4100
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 10008 4100 10149 4128
rect 10008 4088 10014 4100
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 10781 4131 10839 4137
rect 10781 4128 10793 4131
rect 10560 4100 10793 4128
rect 10560 4088 10566 4100
rect 10781 4097 10793 4100
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 10962 4088 10968 4140
rect 11020 4088 11026 4140
rect 11514 4088 11520 4140
rect 11572 4088 11578 4140
rect 12250 4088 12256 4140
rect 12308 4088 12314 4140
rect 12621 4131 12679 4137
rect 12621 4097 12633 4131
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4126 12771 4131
rect 14090 4128 14096 4140
rect 12912 4126 14096 4128
rect 12759 4100 14096 4126
rect 12759 4098 12940 4100
rect 12759 4097 12771 4098
rect 12713 4091 12771 4097
rect 3786 4020 3792 4072
rect 3844 4060 3850 4072
rect 5721 4063 5779 4069
rect 5721 4060 5733 4063
rect 3844 4032 5733 4060
rect 3844 4020 3850 4032
rect 5721 4029 5733 4032
rect 5767 4029 5779 4063
rect 5721 4023 5779 4029
rect 8757 4063 8815 4069
rect 8757 4029 8769 4063
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 8772 3992 8800 4023
rect 9306 4020 9312 4072
rect 9364 4020 9370 4072
rect 9490 4020 9496 4072
rect 9548 4020 9554 4072
rect 9766 4020 9772 4072
rect 9824 4020 9830 4072
rect 10042 4020 10048 4072
rect 10100 4020 10106 4072
rect 10410 4020 10416 4072
rect 10468 4060 10474 4072
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 10468 4032 11621 4060
rect 10468 4020 10474 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 12644 4060 12672 4091
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 14182 4088 14188 4140
rect 14240 4128 14246 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14240 4100 14657 4128
rect 14240 4088 14246 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 14734 4088 14740 4140
rect 14792 4128 14798 4140
rect 17512 4128 17540 4168
rect 14792 4100 17540 4128
rect 14792 4088 14798 4100
rect 17586 4088 17592 4140
rect 17644 4088 17650 4140
rect 17773 4131 17831 4137
rect 17773 4097 17785 4131
rect 17819 4128 17831 4131
rect 18414 4128 18420 4140
rect 17819 4100 18420 4128
rect 17819 4097 17831 4100
rect 17773 4091 17831 4097
rect 18414 4088 18420 4100
rect 18472 4088 18478 4140
rect 13722 4060 13728 4072
rect 12644 4032 13728 4060
rect 11609 4023 11667 4029
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 14366 4020 14372 4072
rect 14424 4020 14430 4072
rect 15102 4020 15108 4072
rect 15160 4020 15166 4072
rect 15930 4020 15936 4072
rect 15988 4020 15994 4072
rect 16853 4063 16911 4069
rect 16853 4029 16865 4063
rect 16899 4060 16911 4063
rect 17494 4060 17500 4072
rect 16899 4032 17500 4060
rect 16899 4029 16911 4032
rect 16853 4023 16911 4029
rect 17494 4020 17500 4032
rect 17552 4020 17558 4072
rect 19306 4060 19334 4168
rect 19797 4165 19809 4199
rect 19843 4196 19855 4199
rect 22738 4196 22744 4208
rect 19843 4168 22744 4196
rect 19843 4165 19855 4168
rect 19797 4159 19855 4165
rect 22738 4156 22744 4168
rect 22796 4156 22802 4208
rect 23124 4205 23152 4236
rect 23198 4224 23204 4236
rect 23256 4224 23262 4276
rect 23937 4267 23995 4273
rect 23937 4233 23949 4267
rect 23983 4233 23995 4267
rect 23937 4227 23995 4233
rect 23109 4199 23167 4205
rect 23109 4165 23121 4199
rect 23155 4165 23167 4199
rect 23109 4159 23167 4165
rect 23216 4168 23520 4196
rect 19886 4088 19892 4140
rect 19944 4088 19950 4140
rect 21082 4128 21088 4140
rect 19996 4100 21088 4128
rect 19996 4060 20024 4100
rect 21082 4088 21088 4100
rect 21140 4128 21146 4140
rect 21269 4131 21327 4137
rect 21269 4128 21281 4131
rect 21140 4100 21281 4128
rect 21140 4088 21146 4100
rect 21269 4097 21281 4100
rect 21315 4097 21327 4131
rect 21269 4091 21327 4097
rect 21634 4088 21640 4140
rect 21692 4128 21698 4140
rect 23216 4128 23244 4168
rect 21692 4100 23244 4128
rect 21692 4088 21698 4100
rect 23382 4088 23388 4140
rect 23440 4088 23446 4140
rect 23492 4137 23520 4168
rect 23842 4156 23848 4208
rect 23900 4196 23906 4208
rect 23952 4196 23980 4227
rect 24302 4224 24308 4276
rect 24360 4264 24366 4276
rect 24360 4236 26464 4264
rect 24360 4224 24366 4236
rect 23900 4168 23980 4196
rect 23900 4156 23906 4168
rect 24026 4156 24032 4208
rect 24084 4196 24090 4208
rect 24946 4196 24952 4208
rect 24084 4168 24952 4196
rect 24084 4156 24090 4168
rect 24946 4156 24952 4168
rect 25004 4156 25010 4208
rect 26436 4140 26464 4236
rect 27706 4224 27712 4276
rect 27764 4264 27770 4276
rect 35618 4264 35624 4276
rect 27764 4236 35624 4264
rect 27764 4224 27770 4236
rect 35618 4224 35624 4236
rect 35676 4224 35682 4276
rect 35894 4224 35900 4276
rect 35952 4264 35958 4276
rect 36725 4267 36783 4273
rect 36725 4264 36737 4267
rect 35952 4236 36737 4264
rect 35952 4224 35958 4236
rect 36725 4233 36737 4236
rect 36771 4264 36783 4267
rect 37366 4264 37372 4276
rect 36771 4236 37372 4264
rect 36771 4233 36783 4236
rect 36725 4227 36783 4233
rect 37366 4224 37372 4236
rect 37424 4224 37430 4276
rect 37550 4224 37556 4276
rect 37608 4264 37614 4276
rect 42334 4264 42340 4276
rect 37608 4236 42340 4264
rect 37608 4224 37614 4236
rect 42334 4224 42340 4236
rect 42392 4224 42398 4276
rect 42518 4224 42524 4276
rect 42576 4264 42582 4276
rect 43717 4267 43775 4273
rect 43717 4264 43729 4267
rect 42576 4236 43729 4264
rect 42576 4224 42582 4236
rect 43717 4233 43729 4236
rect 43763 4233 43775 4267
rect 43717 4227 43775 4233
rect 43990 4224 43996 4276
rect 44048 4264 44054 4276
rect 47121 4267 47179 4273
rect 47121 4264 47133 4267
rect 44048 4236 47133 4264
rect 44048 4224 44054 4236
rect 47121 4233 47133 4236
rect 47167 4233 47179 4267
rect 47121 4227 47179 4233
rect 48314 4224 48320 4276
rect 48372 4224 48378 4276
rect 48774 4224 48780 4276
rect 48832 4264 48838 4276
rect 49145 4267 49203 4273
rect 49145 4264 49157 4267
rect 48832 4236 49157 4264
rect 48832 4224 48838 4236
rect 49145 4233 49157 4236
rect 49191 4233 49203 4267
rect 49145 4227 49203 4233
rect 26970 4156 26976 4208
rect 27028 4196 27034 4208
rect 27893 4199 27951 4205
rect 27893 4196 27905 4199
rect 27028 4168 27905 4196
rect 27028 4156 27034 4168
rect 27893 4165 27905 4168
rect 27939 4165 27951 4199
rect 28258 4196 28264 4208
rect 27893 4159 27951 4165
rect 28000 4168 28264 4196
rect 23477 4131 23535 4137
rect 23477 4097 23489 4131
rect 23523 4097 23535 4131
rect 23477 4091 23535 4097
rect 23753 4131 23811 4137
rect 23753 4097 23765 4131
rect 23799 4128 23811 4131
rect 23799 4100 23888 4128
rect 23799 4097 23811 4100
rect 23753 4091 23811 4097
rect 19306 4032 20024 4060
rect 20254 4020 20260 4072
rect 20312 4020 20318 4072
rect 21358 4020 21364 4072
rect 21416 4020 21422 4072
rect 21545 4063 21603 4069
rect 21545 4029 21557 4063
rect 21591 4060 21603 4063
rect 21726 4060 21732 4072
rect 21591 4032 21732 4060
rect 21591 4029 21603 4032
rect 21545 4023 21603 4029
rect 21726 4020 21732 4032
rect 21784 4020 21790 4072
rect 22005 4063 22063 4069
rect 22005 4029 22017 4063
rect 22051 4060 22063 4063
rect 22278 4060 22284 4072
rect 22051 4032 22284 4060
rect 22051 4029 22063 4032
rect 22005 4023 22063 4029
rect 22278 4020 22284 4032
rect 22336 4020 22342 4072
rect 22557 4063 22615 4069
rect 22557 4029 22569 4063
rect 22603 4060 22615 4063
rect 23658 4060 23664 4072
rect 22603 4032 23664 4060
rect 22603 4029 22615 4032
rect 22557 4023 22615 4029
rect 23658 4020 23664 4032
rect 23716 4020 23722 4072
rect 11974 3992 11980 4004
rect 8772 3964 11980 3992
rect 11974 3952 11980 3964
rect 12032 3952 12038 4004
rect 17310 3992 17316 4004
rect 15672 3964 17316 3992
rect 7377 3927 7435 3933
rect 7377 3893 7389 3927
rect 7423 3924 7435 3927
rect 8478 3924 8484 3936
rect 7423 3896 8484 3924
rect 7423 3893 7435 3896
rect 7377 3887 7435 3893
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 8570 3884 8576 3936
rect 8628 3884 8634 3936
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 15672 3924 15700 3964
rect 17310 3952 17316 3964
rect 17368 3952 17374 4004
rect 17957 3995 18015 4001
rect 17957 3961 17969 3995
rect 18003 3992 18015 3995
rect 18138 3992 18144 4004
rect 18003 3964 18144 3992
rect 18003 3961 18015 3964
rect 17957 3955 18015 3961
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 18509 3995 18567 4001
rect 18509 3961 18521 3995
rect 18555 3992 18567 3995
rect 18598 3992 18604 4004
rect 18555 3964 18604 3992
rect 18555 3961 18567 3964
rect 18509 3955 18567 3961
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 22370 3992 22376 4004
rect 19306 3964 22376 3992
rect 9180 3896 15700 3924
rect 9180 3884 9186 3896
rect 15746 3884 15752 3936
rect 15804 3884 15810 3936
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 16485 3927 16543 3933
rect 16485 3924 16497 3927
rect 16172 3896 16497 3924
rect 16172 3884 16178 3896
rect 16485 3893 16497 3896
rect 16531 3893 16543 3927
rect 16485 3887 16543 3893
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 17589 3927 17647 3933
rect 17589 3924 17601 3927
rect 16632 3896 17601 3924
rect 16632 3884 16638 3896
rect 17589 3893 17601 3896
rect 17635 3924 17647 3927
rect 19306 3924 19334 3964
rect 22370 3952 22376 3964
rect 22428 3952 22434 4004
rect 22738 3952 22744 4004
rect 22796 3952 22802 4004
rect 17635 3896 19334 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 20438 3884 20444 3936
rect 20496 3924 20502 3936
rect 20901 3927 20959 3933
rect 20901 3924 20913 3927
rect 20496 3896 20913 3924
rect 20496 3884 20502 3896
rect 20901 3893 20913 3896
rect 20947 3893 20959 3927
rect 20901 3887 20959 3893
rect 21818 3884 21824 3936
rect 21876 3884 21882 3936
rect 21910 3884 21916 3936
rect 21968 3924 21974 3936
rect 22925 3927 22983 3933
rect 22925 3924 22937 3927
rect 21968 3896 22937 3924
rect 21968 3884 21974 3896
rect 22925 3893 22937 3896
rect 22971 3924 22983 3927
rect 23106 3924 23112 3936
rect 22971 3896 23112 3924
rect 22971 3893 22983 3896
rect 22925 3887 22983 3893
rect 23106 3884 23112 3896
rect 23164 3884 23170 3936
rect 23860 3924 23888 4100
rect 23934 4088 23940 4140
rect 23992 4088 23998 4140
rect 24210 4088 24216 4140
rect 24268 4088 24274 4140
rect 26329 4131 26387 4137
rect 26329 4128 26341 4131
rect 25700 4100 26341 4128
rect 24118 4020 24124 4072
rect 24176 4060 24182 4072
rect 24489 4063 24547 4069
rect 24489 4060 24501 4063
rect 24176 4032 24501 4060
rect 24176 4020 24182 4032
rect 24489 4029 24501 4032
rect 24535 4029 24547 4063
rect 24489 4023 24547 4029
rect 24578 4020 24584 4072
rect 24636 4060 24642 4072
rect 25700 4060 25728 4100
rect 26329 4097 26341 4100
rect 26375 4097 26387 4131
rect 26329 4091 26387 4097
rect 26418 4088 26424 4140
rect 26476 4128 26482 4140
rect 28000 4128 28028 4168
rect 28258 4156 28264 4168
rect 28316 4156 28322 4208
rect 28534 4156 28540 4208
rect 28592 4196 28598 4208
rect 28592 4168 29500 4196
rect 28592 4156 28598 4168
rect 26476 4100 28028 4128
rect 26476 4088 26482 4100
rect 28074 4088 28080 4140
rect 28132 4088 28138 4140
rect 28169 4131 28227 4137
rect 28169 4097 28181 4131
rect 28215 4097 28227 4131
rect 28169 4091 28227 4097
rect 28629 4131 28687 4137
rect 28629 4097 28641 4131
rect 28675 4128 28687 4131
rect 28718 4128 28724 4140
rect 28675 4100 28724 4128
rect 28675 4097 28687 4100
rect 28629 4091 28687 4097
rect 24636 4032 25728 4060
rect 24636 4020 24642 4032
rect 26142 4020 26148 4072
rect 26200 4060 26206 4072
rect 26237 4063 26295 4069
rect 26237 4060 26249 4063
rect 26200 4032 26249 4060
rect 26200 4020 26206 4032
rect 26237 4029 26249 4032
rect 26283 4029 26295 4063
rect 26237 4023 26295 4029
rect 26878 4020 26884 4072
rect 26936 4020 26942 4072
rect 28184 4060 28212 4091
rect 28718 4088 28724 4100
rect 28776 4088 28782 4140
rect 28994 4088 29000 4140
rect 29052 4128 29058 4140
rect 29362 4128 29368 4140
rect 29052 4100 29368 4128
rect 29052 4088 29058 4100
rect 29362 4088 29368 4100
rect 29420 4088 29426 4140
rect 29472 4128 29500 4168
rect 29546 4156 29552 4208
rect 29604 4196 29610 4208
rect 35158 4196 35164 4208
rect 29604 4168 35164 4196
rect 29604 4156 29610 4168
rect 35158 4156 35164 4168
rect 35216 4156 35222 4208
rect 35250 4156 35256 4208
rect 35308 4196 35314 4208
rect 38102 4196 38108 4208
rect 35308 4168 38108 4196
rect 35308 4156 35314 4168
rect 38102 4156 38108 4168
rect 38160 4156 38166 4208
rect 38194 4156 38200 4208
rect 38252 4196 38258 4208
rect 38378 4196 38384 4208
rect 38252 4168 38384 4196
rect 38252 4156 38258 4168
rect 38378 4156 38384 4168
rect 38436 4156 38442 4208
rect 38488 4168 38700 4196
rect 30285 4131 30343 4137
rect 30285 4128 30297 4131
rect 29472 4100 30297 4128
rect 30285 4097 30297 4100
rect 30331 4097 30343 4131
rect 30285 4091 30343 4097
rect 30834 4088 30840 4140
rect 30892 4088 30898 4140
rect 30926 4088 30932 4140
rect 30984 4128 30990 4140
rect 31481 4131 31539 4137
rect 31481 4128 31493 4131
rect 30984 4100 31493 4128
rect 30984 4088 30990 4100
rect 31481 4097 31493 4100
rect 31527 4097 31539 4131
rect 33045 4131 33103 4137
rect 33045 4128 33057 4131
rect 31481 4091 31539 4097
rect 31726 4100 33057 4128
rect 28902 4060 28908 4072
rect 26988 4032 28120 4060
rect 28184 4032 28908 4060
rect 26988 3992 27016 4032
rect 28092 3992 28120 4032
rect 28902 4020 28908 4032
rect 28960 4020 28966 4072
rect 29086 4020 29092 4072
rect 29144 4020 29150 4072
rect 29730 4020 29736 4072
rect 29788 4060 29794 4072
rect 30377 4063 30435 4069
rect 30377 4060 30389 4063
rect 29788 4032 30389 4060
rect 29788 4020 29794 4032
rect 30377 4029 30389 4032
rect 30423 4029 30435 4063
rect 30377 4023 30435 4029
rect 30469 4063 30527 4069
rect 30469 4029 30481 4063
rect 30515 4029 30527 4063
rect 30469 4023 30527 4029
rect 28353 3995 28411 4001
rect 28353 3992 28365 3995
rect 25516 3964 27016 3992
rect 27080 3964 28028 3992
rect 28092 3964 28365 3992
rect 25516 3924 25544 3964
rect 23860 3896 25544 3924
rect 25590 3884 25596 3936
rect 25648 3924 25654 3936
rect 27080 3924 27108 3964
rect 25648 3896 27108 3924
rect 25648 3884 25654 3896
rect 27890 3884 27896 3936
rect 27948 3884 27954 3936
rect 28000 3924 28028 3964
rect 28353 3961 28365 3964
rect 28399 3961 28411 3995
rect 30190 3992 30196 4004
rect 28353 3955 28411 3961
rect 28966 3964 30196 3992
rect 28966 3924 28994 3964
rect 30190 3952 30196 3964
rect 30248 3952 30254 4004
rect 30484 3992 30512 4023
rect 30742 4020 30748 4072
rect 30800 4060 30806 4072
rect 31726 4060 31754 4100
rect 33045 4097 33057 4100
rect 33091 4097 33103 4131
rect 33045 4091 33103 4097
rect 33229 4131 33287 4137
rect 33229 4097 33241 4131
rect 33275 4097 33287 4131
rect 33229 4091 33287 4097
rect 30800 4032 31754 4060
rect 30800 4020 30806 4032
rect 31938 4020 31944 4072
rect 31996 4020 32002 4072
rect 32398 4020 32404 4072
rect 32456 4060 32462 4072
rect 33244 4060 33272 4091
rect 33778 4088 33784 4140
rect 33836 4128 33842 4140
rect 33965 4131 34023 4137
rect 33965 4128 33977 4131
rect 33836 4100 33977 4128
rect 33836 4088 33842 4100
rect 33965 4097 33977 4100
rect 34011 4097 34023 4131
rect 33965 4091 34023 4097
rect 34054 4088 34060 4140
rect 34112 4088 34118 4140
rect 36265 4131 36323 4137
rect 36265 4097 36277 4131
rect 36311 4128 36323 4131
rect 36630 4128 36636 4140
rect 36311 4100 36636 4128
rect 36311 4097 36323 4100
rect 36265 4091 36323 4097
rect 36630 4088 36636 4100
rect 36688 4088 36694 4140
rect 36817 4131 36875 4137
rect 36817 4097 36829 4131
rect 36863 4128 36875 4131
rect 37458 4128 37464 4140
rect 36863 4100 37464 4128
rect 36863 4097 36875 4100
rect 36817 4091 36875 4097
rect 37458 4088 37464 4100
rect 37516 4088 37522 4140
rect 37550 4088 37556 4140
rect 37608 4128 37614 4140
rect 38488 4137 38516 4168
rect 38013 4131 38071 4137
rect 38013 4128 38025 4131
rect 37608 4100 38025 4128
rect 37608 4088 37614 4100
rect 38013 4097 38025 4100
rect 38059 4097 38071 4131
rect 38013 4091 38071 4097
rect 38473 4131 38531 4137
rect 38473 4097 38485 4131
rect 38519 4097 38531 4131
rect 38473 4091 38531 4097
rect 38562 4088 38568 4140
rect 38620 4088 38626 4140
rect 38672 4128 38700 4168
rect 40328 4168 40632 4196
rect 39206 4128 39212 4140
rect 38672 4100 39212 4128
rect 39206 4088 39212 4100
rect 39264 4088 39270 4140
rect 39482 4088 39488 4140
rect 39540 4128 39546 4140
rect 40328 4128 40356 4168
rect 39540 4100 40356 4128
rect 39540 4088 39546 4100
rect 40402 4088 40408 4140
rect 40460 4088 40466 4140
rect 40494 4088 40500 4140
rect 40552 4088 40558 4140
rect 40604 4128 40632 4168
rect 43346 4156 43352 4208
rect 43404 4196 43410 4208
rect 43404 4168 47072 4196
rect 43404 4156 43410 4168
rect 41049 4131 41107 4137
rect 40604 4100 40724 4128
rect 32456 4032 33272 4060
rect 32456 4020 32462 4032
rect 33410 4020 33416 4072
rect 33468 4020 33474 4072
rect 35250 4020 35256 4072
rect 35308 4020 35314 4072
rect 35713 4063 35771 4069
rect 35713 4029 35725 4063
rect 35759 4029 35771 4063
rect 35713 4023 35771 4029
rect 31846 3992 31852 4004
rect 30395 3964 31852 3992
rect 28000 3896 28994 3924
rect 29914 3884 29920 3936
rect 29972 3884 29978 3936
rect 30098 3884 30104 3936
rect 30156 3924 30162 3936
rect 30395 3924 30423 3964
rect 31846 3952 31852 3964
rect 31904 3952 31910 4004
rect 33226 3952 33232 4004
rect 33284 3952 33290 4004
rect 33318 3952 33324 4004
rect 33376 3992 33382 4004
rect 35728 3992 35756 4023
rect 36078 4020 36084 4072
rect 36136 4060 36142 4072
rect 36722 4060 36728 4072
rect 36136 4032 36728 4060
rect 36136 4020 36142 4032
rect 36722 4020 36728 4032
rect 36780 4020 36786 4072
rect 36906 4020 36912 4072
rect 36964 4020 36970 4072
rect 37734 4020 37740 4072
rect 37792 4020 37798 4072
rect 38102 4020 38108 4072
rect 38160 4060 38166 4072
rect 39025 4063 39083 4069
rect 39025 4060 39037 4063
rect 38160 4032 39037 4060
rect 38160 4020 38166 4032
rect 39025 4029 39037 4032
rect 39071 4029 39083 4063
rect 39025 4023 39083 4029
rect 40310 4020 40316 4072
rect 40368 4060 40374 4072
rect 40589 4063 40647 4069
rect 40589 4060 40601 4063
rect 40368 4032 40601 4060
rect 40368 4020 40374 4032
rect 40589 4029 40601 4032
rect 40635 4029 40647 4063
rect 40696 4060 40724 4100
rect 41049 4097 41061 4131
rect 41095 4128 41107 4131
rect 41095 4100 42472 4128
rect 41095 4097 41107 4100
rect 41049 4091 41107 4097
rect 41141 4063 41199 4069
rect 41141 4060 41153 4063
rect 40696 4032 41153 4060
rect 40589 4023 40647 4029
rect 41141 4029 41153 4032
rect 41187 4029 41199 4063
rect 41141 4023 41199 4029
rect 41785 4063 41843 4069
rect 41785 4029 41797 4063
rect 41831 4060 41843 4063
rect 42058 4060 42064 4072
rect 41831 4032 42064 4060
rect 41831 4029 41843 4032
rect 41785 4023 41843 4029
rect 42058 4020 42064 4032
rect 42116 4020 42122 4072
rect 42444 4060 42472 4100
rect 42518 4088 42524 4140
rect 42576 4088 42582 4140
rect 42702 4088 42708 4140
rect 42760 4128 42766 4140
rect 42981 4131 43039 4137
rect 42981 4128 42993 4131
rect 42760 4100 42993 4128
rect 42760 4088 42766 4100
rect 42981 4097 42993 4100
rect 43027 4097 43039 4131
rect 42981 4091 43039 4097
rect 43254 4088 43260 4140
rect 43312 4128 43318 4140
rect 46385 4131 46443 4137
rect 46385 4128 46397 4131
rect 43312 4100 46397 4128
rect 43312 4088 43318 4100
rect 46385 4097 46397 4100
rect 46431 4097 46443 4131
rect 46385 4091 46443 4097
rect 46474 4088 46480 4140
rect 46532 4128 46538 4140
rect 46937 4131 46995 4137
rect 46937 4128 46949 4131
rect 46532 4100 46949 4128
rect 46532 4088 46538 4100
rect 46937 4097 46949 4100
rect 46983 4097 46995 4131
rect 47044 4128 47072 4168
rect 47044 4100 47900 4128
rect 46937 4091 46995 4097
rect 42794 4060 42800 4072
rect 42444 4032 42800 4060
rect 42794 4020 42800 4032
rect 42852 4020 42858 4072
rect 42886 4020 42892 4072
rect 42944 4020 42950 4072
rect 43070 4020 43076 4072
rect 43128 4060 43134 4072
rect 43441 4063 43499 4069
rect 43441 4060 43453 4063
rect 43128 4032 43453 4060
rect 43128 4020 43134 4032
rect 43441 4029 43453 4032
rect 43487 4029 43499 4063
rect 43441 4023 43499 4029
rect 43625 4063 43683 4069
rect 43625 4029 43637 4063
rect 43671 4060 43683 4063
rect 43671 4032 44036 4060
rect 43671 4029 43683 4032
rect 43625 4023 43683 4029
rect 33376 3964 34100 3992
rect 35728 3964 36492 3992
rect 33376 3952 33382 3964
rect 30156 3896 30423 3924
rect 30156 3884 30162 3896
rect 31386 3884 31392 3936
rect 31444 3884 31450 3936
rect 32490 3884 32496 3936
rect 32548 3924 32554 3936
rect 33870 3924 33876 3936
rect 32548 3896 33876 3924
rect 32548 3884 32554 3896
rect 33870 3884 33876 3896
rect 33928 3884 33934 3936
rect 34072 3924 34100 3964
rect 36357 3927 36415 3933
rect 36357 3924 36369 3927
rect 34072 3896 36369 3924
rect 36357 3893 36369 3896
rect 36403 3893 36415 3927
rect 36464 3924 36492 3964
rect 36648 3964 40172 3992
rect 36648 3924 36676 3964
rect 36464 3896 36676 3924
rect 36357 3887 36415 3893
rect 36722 3884 36728 3936
rect 36780 3924 36786 3936
rect 38289 3927 38347 3933
rect 38289 3924 38301 3927
rect 36780 3896 38301 3924
rect 36780 3884 36786 3896
rect 38289 3893 38301 3896
rect 38335 3893 38347 3927
rect 38289 3887 38347 3893
rect 39942 3884 39948 3936
rect 40000 3924 40006 3936
rect 40037 3927 40095 3933
rect 40037 3924 40049 3927
rect 40000 3896 40049 3924
rect 40000 3884 40006 3896
rect 40037 3893 40049 3896
rect 40083 3893 40095 3927
rect 40144 3924 40172 3964
rect 40865 3927 40923 3933
rect 40865 3924 40877 3927
rect 40144 3896 40877 3924
rect 40037 3887 40095 3893
rect 40865 3893 40877 3896
rect 40911 3893 40923 3927
rect 40865 3887 40923 3893
rect 41230 3884 41236 3936
rect 41288 3924 41294 3936
rect 41877 3927 41935 3933
rect 41877 3924 41889 3927
rect 41288 3896 41889 3924
rect 41288 3884 41294 3896
rect 41877 3893 41889 3896
rect 41923 3893 41935 3927
rect 41877 3887 41935 3893
rect 42334 3884 42340 3936
rect 42392 3924 42398 3936
rect 42705 3927 42763 3933
rect 42705 3924 42717 3927
rect 42392 3896 42717 3924
rect 42392 3884 42398 3896
rect 42705 3893 42717 3896
rect 42751 3893 42763 3927
rect 42705 3887 42763 3893
rect 42794 3884 42800 3936
rect 42852 3924 42858 3936
rect 43806 3924 43812 3936
rect 42852 3896 43812 3924
rect 42852 3884 42858 3896
rect 43806 3884 43812 3896
rect 43864 3884 43870 3936
rect 44008 3924 44036 4032
rect 44174 4020 44180 4072
rect 44232 4020 44238 4072
rect 44284 4032 44680 4060
rect 44085 3995 44143 4001
rect 44085 3961 44097 3995
rect 44131 3992 44143 3995
rect 44284 3992 44312 4032
rect 44131 3964 44312 3992
rect 44652 3992 44680 4032
rect 44726 4020 44732 4072
rect 44784 4020 44790 4072
rect 45557 4063 45615 4069
rect 45557 4029 45569 4063
rect 45603 4029 45615 4063
rect 45557 4023 45615 4029
rect 45572 3992 45600 4023
rect 45646 4020 45652 4072
rect 45704 4020 45710 4072
rect 46293 4063 46351 4069
rect 46293 4029 46305 4063
rect 46339 4029 46351 4063
rect 46293 4023 46351 4029
rect 47765 4063 47823 4069
rect 47765 4029 47777 4063
rect 47811 4029 47823 4063
rect 47872 4060 47900 4100
rect 48038 4088 48044 4140
rect 48096 4088 48102 4140
rect 48133 4131 48191 4137
rect 48133 4097 48145 4131
rect 48179 4097 48191 4131
rect 48133 4091 48191 4097
rect 48148 4060 48176 4091
rect 48498 4088 48504 4140
rect 48556 4088 48562 4140
rect 74626 4088 74632 4140
rect 74684 4128 74690 4140
rect 74721 4131 74779 4137
rect 74721 4128 74733 4131
rect 74684 4100 74733 4128
rect 74684 4088 74690 4100
rect 74721 4097 74733 4100
rect 74767 4097 74779 4131
rect 76193 4131 76251 4137
rect 76193 4128 76205 4131
rect 74721 4091 74779 4097
rect 75288 4100 76205 4128
rect 47872 4032 48176 4060
rect 49237 4063 49295 4069
rect 47765 4023 47823 4029
rect 49237 4029 49249 4063
rect 49283 4029 49295 4063
rect 49237 4023 49295 4029
rect 52181 4063 52239 4069
rect 52181 4029 52193 4063
rect 52227 4060 52239 4063
rect 53190 4060 53196 4072
rect 52227 4032 53196 4060
rect 52227 4029 52239 4032
rect 52181 4023 52239 4029
rect 44652 3964 45600 3992
rect 46308 3992 46336 4023
rect 47578 3992 47584 4004
rect 46308 3964 47584 3992
rect 44131 3961 44143 3964
rect 44085 3955 44143 3961
rect 47578 3952 47584 3964
rect 47636 3952 47642 4004
rect 47780 3992 47808 4023
rect 47857 3995 47915 4001
rect 47857 3992 47869 3995
rect 47780 3964 47869 3992
rect 47857 3961 47869 3964
rect 47903 3961 47915 3995
rect 47857 3955 47915 3961
rect 44818 3924 44824 3936
rect 44008 3896 44824 3924
rect 44818 3884 44824 3896
rect 44876 3884 44882 3936
rect 44910 3884 44916 3936
rect 44968 3884 44974 3936
rect 46382 3884 46388 3936
rect 46440 3924 46446 3936
rect 49252 3924 49280 4023
rect 53190 4020 53196 4032
rect 53248 4020 53254 4072
rect 53834 4020 53840 4072
rect 53892 4020 53898 4072
rect 65426 4020 65432 4072
rect 65484 4060 65490 4072
rect 65521 4063 65579 4069
rect 65521 4060 65533 4063
rect 65484 4032 65533 4060
rect 65484 4020 65490 4032
rect 65521 4029 65533 4032
rect 65567 4029 65579 4063
rect 65521 4023 65579 4029
rect 67637 4063 67695 4069
rect 67637 4029 67649 4063
rect 67683 4060 67695 4063
rect 68646 4060 68652 4072
rect 67683 4032 68652 4060
rect 67683 4029 67695 4032
rect 67637 4023 67695 4029
rect 68646 4020 68652 4032
rect 68704 4020 68710 4072
rect 69290 4020 69296 4072
rect 69348 4020 69354 4072
rect 71501 4063 71559 4069
rect 71501 4029 71513 4063
rect 71547 4060 71559 4063
rect 71682 4060 71688 4072
rect 71547 4032 71688 4060
rect 71547 4029 71559 4032
rect 71501 4023 71559 4029
rect 71682 4020 71688 4032
rect 71740 4020 71746 4072
rect 74258 4020 74264 4072
rect 74316 4060 74322 4072
rect 75288 4060 75316 4100
rect 76193 4097 76205 4100
rect 76239 4097 76251 4131
rect 76193 4091 76251 4097
rect 74316 4032 75316 4060
rect 75917 4063 75975 4069
rect 74316 4020 74322 4032
rect 75917 4029 75929 4063
rect 75963 4060 75975 4063
rect 76558 4060 76564 4072
rect 75963 4032 76564 4060
rect 75963 4029 75975 4032
rect 75917 4023 75975 4029
rect 76558 4020 76564 4032
rect 76616 4020 76622 4072
rect 77018 4020 77024 4072
rect 77076 4020 77082 4072
rect 46440 3896 49280 3924
rect 49881 3927 49939 3933
rect 46440 3884 46446 3896
rect 49881 3893 49893 3927
rect 49927 3924 49939 3927
rect 51350 3924 51356 3936
rect 49927 3896 51356 3924
rect 49927 3893 49939 3896
rect 49881 3887 49939 3893
rect 51350 3884 51356 3896
rect 51408 3884 51414 3936
rect 52733 3927 52791 3933
rect 52733 3893 52745 3927
rect 52779 3924 52791 3927
rect 52822 3924 52828 3936
rect 52779 3896 52828 3924
rect 52779 3893 52791 3896
rect 52733 3887 52791 3893
rect 52822 3884 52828 3896
rect 52880 3884 52886 3936
rect 54018 3884 54024 3936
rect 54076 3924 54082 3936
rect 54389 3927 54447 3933
rect 54389 3924 54401 3927
rect 54076 3896 54401 3924
rect 54076 3884 54082 3896
rect 54389 3893 54401 3896
rect 54435 3893 54447 3927
rect 54389 3887 54447 3893
rect 66165 3927 66223 3933
rect 66165 3893 66177 3927
rect 66211 3924 66223 3927
rect 66254 3924 66260 3936
rect 66211 3896 66260 3924
rect 66211 3893 66223 3896
rect 66165 3887 66223 3893
rect 66254 3884 66260 3896
rect 66312 3884 66318 3936
rect 68189 3927 68247 3933
rect 68189 3893 68201 3927
rect 68235 3924 68247 3927
rect 68278 3924 68284 3936
rect 68235 3896 68284 3924
rect 68235 3893 68247 3896
rect 68189 3887 68247 3893
rect 68278 3884 68284 3896
rect 68336 3884 68342 3936
rect 69474 3884 69480 3936
rect 69532 3924 69538 3936
rect 69845 3927 69903 3933
rect 69845 3924 69857 3927
rect 69532 3896 69857 3924
rect 69532 3884 69538 3896
rect 69845 3893 69857 3896
rect 69891 3893 69903 3927
rect 69845 3887 69903 3893
rect 72053 3927 72111 3933
rect 72053 3893 72065 3927
rect 72099 3924 72111 3927
rect 73706 3924 73712 3936
rect 72099 3896 73712 3924
rect 72099 3893 72111 3896
rect 72053 3887 72111 3893
rect 73706 3884 73712 3896
rect 73764 3884 73770 3936
rect 2024 3834 77924 3856
rect 2024 3782 5134 3834
rect 5186 3782 5198 3834
rect 5250 3782 5262 3834
rect 5314 3782 5326 3834
rect 5378 3782 5390 3834
rect 5442 3782 35854 3834
rect 35906 3782 35918 3834
rect 35970 3782 35982 3834
rect 36034 3782 36046 3834
rect 36098 3782 36110 3834
rect 36162 3782 66574 3834
rect 66626 3782 66638 3834
rect 66690 3782 66702 3834
rect 66754 3782 66766 3834
rect 66818 3782 66830 3834
rect 66882 3782 77924 3834
rect 2024 3760 77924 3782
rect 5813 3723 5871 3729
rect 5813 3689 5825 3723
rect 5859 3720 5871 3723
rect 6638 3720 6644 3732
rect 5859 3692 6644 3720
rect 5859 3689 5871 3692
rect 5813 3683 5871 3689
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 8628 3692 13676 3720
rect 8628 3680 8634 3692
rect 7285 3655 7343 3661
rect 7285 3621 7297 3655
rect 7331 3652 7343 3655
rect 13648 3652 13676 3692
rect 13722 3680 13728 3732
rect 13780 3680 13786 3732
rect 14826 3680 14832 3732
rect 14884 3680 14890 3732
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15344 3692 15516 3720
rect 15344 3680 15350 3692
rect 15488 3652 15516 3692
rect 15930 3680 15936 3732
rect 15988 3720 15994 3732
rect 15988 3692 19012 3720
rect 15988 3680 15994 3692
rect 16117 3655 16175 3661
rect 16117 3652 16129 3655
rect 7331 3624 11744 3652
rect 13648 3624 15424 3652
rect 15488 3624 16129 3652
rect 7331 3621 7343 3624
rect 7285 3615 7343 3621
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 6822 3584 6828 3596
rect 6595 3556 6828 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 9677 3587 9735 3593
rect 8251 3556 9628 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 5258 3476 5264 3528
rect 5316 3476 5322 3528
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3516 6791 3519
rect 7377 3519 7435 3525
rect 7377 3516 7389 3519
rect 6779 3488 7389 3516
rect 6779 3485 6791 3488
rect 6733 3479 6791 3485
rect 7377 3485 7389 3488
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3516 8079 3519
rect 8754 3516 8760 3528
rect 8067 3488 8760 3516
rect 8067 3485 8079 3488
rect 8021 3479 8079 3485
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 9033 3519 9091 3525
rect 9033 3485 9045 3519
rect 9079 3485 9091 3519
rect 9600 3516 9628 3556
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 9858 3584 9864 3596
rect 9723 3556 9864 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 9858 3544 9864 3556
rect 9916 3544 9922 3596
rect 10229 3587 10287 3593
rect 10229 3553 10241 3587
rect 10275 3584 10287 3587
rect 10410 3584 10416 3596
rect 10275 3556 10416 3584
rect 10275 3553 10287 3556
rect 10229 3547 10287 3553
rect 10410 3544 10416 3556
rect 10468 3544 10474 3596
rect 10870 3544 10876 3596
rect 10928 3544 10934 3596
rect 11716 3584 11744 3624
rect 12253 3587 12311 3593
rect 12253 3584 12265 3587
rect 11716 3556 12265 3584
rect 12253 3553 12265 3556
rect 12299 3553 12311 3587
rect 12253 3547 12311 3553
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 12400 3556 13860 3584
rect 12400 3544 12406 3556
rect 10042 3516 10048 3528
rect 9600 3488 10048 3516
rect 9033 3479 9091 3485
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 5905 3451 5963 3457
rect 5905 3448 5917 3451
rect 4212 3420 5917 3448
rect 4212 3408 4218 3420
rect 5905 3417 5917 3420
rect 5951 3417 5963 3451
rect 5905 3411 5963 3417
rect 9048 3392 9076 3479
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 11977 3519 12035 3525
rect 11977 3485 11989 3519
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 10502 3408 10508 3460
rect 10560 3448 10566 3460
rect 11992 3448 12020 3479
rect 10560 3420 12020 3448
rect 10560 3408 10566 3420
rect 8757 3383 8815 3389
rect 8757 3349 8769 3383
rect 8803 3380 8815 3383
rect 8846 3380 8852 3392
rect 8803 3352 8852 3380
rect 8803 3349 8815 3352
rect 8757 3343 8815 3349
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 8941 3383 8999 3389
rect 8941 3349 8953 3383
rect 8987 3380 8999 3383
rect 9030 3380 9036 3392
rect 8987 3352 9036 3380
rect 8987 3349 8999 3352
rect 8941 3343 8999 3349
rect 9030 3340 9036 3352
rect 9088 3340 9094 3392
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 10410 3380 10416 3392
rect 9640 3352 10416 3380
rect 9640 3340 9646 3352
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 10781 3383 10839 3389
rect 10781 3349 10793 3383
rect 10827 3380 10839 3383
rect 10962 3380 10968 3392
rect 10827 3352 10968 3380
rect 10827 3349 10839 3352
rect 10781 3343 10839 3349
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11514 3340 11520 3392
rect 11572 3340 11578 3392
rect 11992 3380 12020 3420
rect 12342 3408 12348 3460
rect 12400 3448 12406 3460
rect 12400 3420 12742 3448
rect 12400 3408 12406 3420
rect 13078 3380 13084 3392
rect 11992 3352 13084 3380
rect 13078 3340 13084 3352
rect 13136 3340 13142 3392
rect 13832 3389 13860 3556
rect 14090 3544 14096 3596
rect 14148 3584 14154 3596
rect 14369 3587 14427 3593
rect 14369 3584 14381 3587
rect 14148 3556 14381 3584
rect 14148 3544 14154 3556
rect 14369 3553 14381 3556
rect 14415 3584 14427 3587
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 14415 3556 15301 3584
rect 14415 3553 14427 3556
rect 14369 3547 14427 3553
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 15396 3584 15424 3624
rect 16117 3621 16129 3624
rect 16163 3652 16175 3655
rect 16390 3652 16396 3664
rect 16163 3624 16396 3652
rect 16163 3621 16175 3624
rect 16117 3615 16175 3621
rect 16390 3612 16396 3624
rect 16448 3612 16454 3664
rect 18984 3652 19012 3692
rect 19886 3680 19892 3732
rect 19944 3720 19950 3732
rect 19981 3723 20039 3729
rect 19981 3720 19993 3723
rect 19944 3692 19993 3720
rect 19944 3680 19950 3692
rect 19981 3689 19993 3692
rect 20027 3689 20039 3723
rect 19981 3683 20039 3689
rect 20070 3680 20076 3732
rect 20128 3720 20134 3732
rect 22005 3723 22063 3729
rect 22005 3720 22017 3723
rect 20128 3692 22017 3720
rect 20128 3680 20134 3692
rect 22005 3689 22017 3692
rect 22051 3689 22063 3723
rect 22005 3683 22063 3689
rect 25593 3723 25651 3729
rect 25593 3689 25605 3723
rect 25639 3720 25651 3723
rect 27706 3720 27712 3732
rect 25639 3692 27712 3720
rect 25639 3689 25651 3692
rect 25593 3683 25651 3689
rect 27706 3680 27712 3692
rect 27764 3680 27770 3732
rect 28074 3680 28080 3732
rect 28132 3720 28138 3732
rect 29546 3720 29552 3732
rect 28132 3692 29552 3720
rect 28132 3680 28138 3692
rect 29546 3680 29552 3692
rect 29604 3720 29610 3732
rect 31294 3720 31300 3732
rect 29604 3692 31300 3720
rect 29604 3680 29610 3692
rect 31294 3680 31300 3692
rect 31352 3720 31358 3732
rect 33042 3720 33048 3732
rect 31352 3692 33048 3720
rect 31352 3680 31358 3692
rect 33042 3680 33048 3692
rect 33100 3680 33106 3732
rect 33962 3680 33968 3732
rect 34020 3720 34026 3732
rect 34057 3723 34115 3729
rect 34057 3720 34069 3723
rect 34020 3692 34069 3720
rect 34020 3680 34026 3692
rect 34057 3689 34069 3692
rect 34103 3689 34115 3723
rect 34057 3683 34115 3689
rect 34698 3680 34704 3732
rect 34756 3680 34762 3732
rect 36906 3720 36912 3732
rect 35268 3692 36912 3720
rect 17696 3624 18736 3652
rect 18984 3624 22324 3652
rect 16669 3587 16727 3593
rect 16669 3584 16681 3587
rect 15396 3556 16681 3584
rect 15289 3547 15347 3553
rect 16669 3553 16681 3556
rect 16715 3553 16727 3587
rect 16669 3547 16727 3553
rect 16758 3544 16764 3596
rect 16816 3584 16822 3596
rect 17696 3584 17724 3624
rect 16816 3556 17724 3584
rect 16816 3544 16822 3556
rect 17862 3544 17868 3596
rect 17920 3544 17926 3596
rect 18138 3544 18144 3596
rect 18196 3544 18202 3596
rect 18708 3593 18736 3624
rect 18693 3587 18751 3593
rect 18693 3553 18705 3587
rect 18739 3553 18751 3587
rect 18693 3547 18751 3553
rect 20070 3544 20076 3596
rect 20128 3584 20134 3596
rect 20809 3587 20867 3593
rect 20809 3584 20821 3587
rect 20128 3556 20821 3584
rect 20128 3544 20134 3556
rect 20809 3553 20821 3556
rect 20855 3553 20867 3587
rect 20809 3547 20867 3553
rect 20990 3544 20996 3596
rect 21048 3584 21054 3596
rect 22296 3584 22324 3624
rect 22370 3612 22376 3664
rect 22428 3652 22434 3664
rect 24946 3652 24952 3664
rect 22428 3624 24952 3652
rect 22428 3612 22434 3624
rect 24946 3612 24952 3624
rect 25004 3612 25010 3664
rect 25314 3612 25320 3664
rect 25372 3652 25378 3664
rect 25682 3652 25688 3664
rect 25372 3624 25688 3652
rect 25372 3612 25378 3624
rect 25682 3612 25688 3624
rect 25740 3612 25746 3664
rect 26510 3612 26516 3664
rect 26568 3612 26574 3664
rect 27982 3612 27988 3664
rect 28040 3652 28046 3664
rect 28040 3624 28396 3652
rect 28040 3612 28046 3624
rect 23937 3587 23995 3593
rect 23937 3584 23949 3587
rect 21048 3556 22094 3584
rect 22296 3556 23949 3584
rect 21048 3544 21054 3556
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14185 3519 14243 3525
rect 14185 3516 14197 3519
rect 14056 3488 14197 3516
rect 14056 3476 14062 3488
rect 14185 3485 14197 3488
rect 14231 3485 14243 3519
rect 14185 3479 14243 3485
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 14458 3516 14464 3528
rect 14323 3488 14464 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 14200 3448 14228 3479
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14642 3476 14648 3528
rect 14700 3476 14706 3528
rect 15194 3476 15200 3528
rect 15252 3516 15258 3528
rect 15562 3516 15568 3528
rect 15252 3488 15568 3516
rect 15252 3476 15258 3488
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 16298 3476 16304 3528
rect 16356 3476 16362 3528
rect 16393 3519 16451 3525
rect 16393 3485 16405 3519
rect 16439 3485 16451 3519
rect 17880 3516 17908 3544
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 17880 3488 18245 3516
rect 16393 3479 16451 3485
rect 18233 3485 18245 3488
rect 18279 3485 18291 3519
rect 18233 3479 18291 3485
rect 19797 3519 19855 3525
rect 19797 3485 19809 3519
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 14734 3448 14740 3460
rect 14200 3420 14740 3448
rect 14734 3408 14740 3420
rect 14792 3408 14798 3460
rect 14918 3408 14924 3460
rect 14976 3448 14982 3460
rect 16408 3448 16436 3479
rect 19812 3448 19840 3479
rect 19886 3476 19892 3528
rect 19944 3516 19950 3528
rect 20349 3519 20407 3525
rect 20349 3516 20361 3519
rect 19944 3488 20361 3516
rect 19944 3476 19950 3488
rect 20349 3485 20361 3488
rect 20395 3485 20407 3519
rect 22066 3516 22094 3556
rect 23937 3553 23949 3556
rect 23983 3553 23995 3587
rect 23937 3547 23995 3553
rect 26329 3587 26387 3593
rect 26329 3553 26341 3587
rect 26375 3584 26387 3587
rect 26418 3584 26424 3596
rect 26375 3556 26424 3584
rect 26375 3553 26387 3556
rect 26329 3547 26387 3553
rect 26418 3544 26424 3556
rect 26476 3544 26482 3596
rect 27430 3544 27436 3596
rect 27488 3584 27494 3596
rect 27488 3556 28304 3584
rect 27488 3544 27494 3556
rect 22281 3519 22339 3525
rect 22281 3516 22293 3519
rect 22066 3488 22293 3516
rect 20349 3479 20407 3485
rect 22281 3485 22293 3488
rect 22327 3485 22339 3519
rect 22281 3479 22339 3485
rect 23382 3476 23388 3528
rect 23440 3516 23446 3528
rect 24026 3516 24032 3528
rect 23440 3488 24032 3516
rect 23440 3476 23446 3488
rect 24026 3476 24032 3488
rect 24084 3476 24090 3528
rect 25133 3519 25191 3525
rect 25133 3485 25145 3519
rect 25179 3516 25191 3519
rect 25222 3516 25228 3528
rect 25179 3488 25228 3516
rect 25179 3485 25191 3488
rect 25133 3479 25191 3485
rect 25222 3476 25228 3488
rect 25280 3476 25286 3528
rect 25314 3476 25320 3528
rect 25372 3476 25378 3528
rect 26697 3519 26755 3525
rect 26697 3516 26709 3519
rect 25424 3488 26709 3516
rect 20254 3448 20260 3460
rect 14976 3420 16436 3448
rect 17894 3420 19334 3448
rect 19812 3420 20260 3448
rect 14976 3408 14982 3420
rect 13817 3383 13875 3389
rect 13817 3349 13829 3383
rect 13863 3349 13875 3383
rect 13817 3343 13875 3349
rect 14550 3340 14556 3392
rect 14608 3380 14614 3392
rect 15473 3383 15531 3389
rect 15473 3380 15485 3383
rect 14608 3352 15485 3380
rect 14608 3340 14614 3352
rect 15473 3349 15485 3352
rect 15519 3349 15531 3383
rect 15473 3343 15531 3349
rect 15930 3340 15936 3392
rect 15988 3340 15994 3392
rect 16408 3380 16436 3420
rect 19306 3392 19334 3420
rect 20254 3408 20260 3420
rect 20312 3408 20318 3460
rect 21266 3408 21272 3460
rect 21324 3448 21330 3460
rect 21910 3448 21916 3460
rect 21324 3420 21916 3448
rect 21324 3408 21330 3420
rect 21910 3408 21916 3420
rect 21968 3457 21974 3460
rect 21968 3451 22031 3457
rect 21968 3417 21985 3451
rect 22019 3417 22031 3451
rect 21968 3411 22031 3417
rect 21968 3408 21974 3411
rect 22186 3408 22192 3460
rect 22244 3408 22250 3460
rect 22462 3408 22468 3460
rect 22520 3448 22526 3460
rect 23201 3451 23259 3457
rect 23201 3448 23213 3451
rect 22520 3420 23213 3448
rect 22520 3408 22526 3420
rect 23201 3417 23213 3420
rect 23247 3417 23259 3451
rect 25424 3448 25452 3488
rect 26697 3485 26709 3488
rect 26743 3485 26755 3519
rect 26697 3479 26755 3485
rect 28074 3476 28080 3528
rect 28132 3476 28138 3528
rect 23201 3411 23259 3417
rect 24780 3420 25452 3448
rect 24780 3392 24808 3420
rect 25590 3408 25596 3460
rect 25648 3408 25654 3460
rect 25866 3408 25872 3460
rect 25924 3448 25930 3460
rect 26053 3451 26111 3457
rect 26053 3448 26065 3451
rect 25924 3420 26065 3448
rect 25924 3408 25930 3420
rect 26053 3417 26065 3420
rect 26099 3417 26111 3451
rect 26053 3411 26111 3417
rect 26142 3408 26148 3460
rect 26200 3408 26206 3460
rect 26973 3451 27031 3457
rect 26973 3417 26985 3451
rect 27019 3448 27031 3451
rect 27246 3448 27252 3460
rect 27019 3420 27252 3448
rect 27019 3417 27031 3420
rect 26973 3411 27031 3417
rect 27246 3408 27252 3420
rect 27304 3408 27310 3460
rect 28276 3448 28304 3556
rect 28368 3516 28396 3624
rect 28442 3612 28448 3664
rect 28500 3612 28506 3664
rect 30374 3652 30380 3664
rect 28644 3624 30380 3652
rect 28644 3516 28672 3624
rect 30374 3612 30380 3624
rect 30432 3612 30438 3664
rect 32030 3612 32036 3664
rect 32088 3612 32094 3664
rect 34609 3655 34667 3661
rect 34609 3621 34621 3655
rect 34655 3652 34667 3655
rect 34974 3652 34980 3664
rect 34655 3624 34980 3652
rect 34655 3621 34667 3624
rect 34609 3615 34667 3621
rect 34974 3612 34980 3624
rect 35032 3612 35038 3664
rect 29362 3544 29368 3596
rect 29420 3544 29426 3596
rect 30098 3544 30104 3596
rect 30156 3584 30162 3596
rect 30650 3584 30656 3596
rect 30156 3556 30656 3584
rect 30156 3544 30162 3556
rect 30650 3544 30656 3556
rect 30708 3544 30714 3596
rect 31202 3544 31208 3596
rect 31260 3584 31266 3596
rect 32122 3584 32128 3596
rect 31260 3556 32128 3584
rect 31260 3544 31266 3556
rect 32122 3544 32128 3556
rect 32180 3584 32186 3596
rect 32309 3587 32367 3593
rect 32309 3584 32321 3587
rect 32180 3556 32321 3584
rect 32180 3544 32186 3556
rect 32309 3553 32321 3556
rect 32355 3584 32367 3587
rect 32582 3584 32588 3596
rect 32355 3556 32588 3584
rect 32355 3553 32367 3556
rect 32309 3547 32367 3553
rect 32582 3544 32588 3556
rect 32640 3544 32646 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 35268 3593 35296 3692
rect 36906 3680 36912 3692
rect 36964 3720 36970 3732
rect 40310 3720 40316 3732
rect 36964 3692 40316 3720
rect 36964 3680 36970 3692
rect 40310 3680 40316 3692
rect 40368 3680 40374 3732
rect 41233 3723 41291 3729
rect 41233 3689 41245 3723
rect 41279 3720 41291 3723
rect 41506 3720 41512 3732
rect 41279 3692 41512 3720
rect 41279 3689 41291 3692
rect 41233 3683 41291 3689
rect 41506 3680 41512 3692
rect 41564 3680 41570 3732
rect 41874 3680 41880 3732
rect 41932 3720 41938 3732
rect 41969 3723 42027 3729
rect 41969 3720 41981 3723
rect 41932 3692 41981 3720
rect 41932 3680 41938 3692
rect 41969 3689 41981 3692
rect 42015 3689 42027 3723
rect 41969 3683 42027 3689
rect 43551 3723 43609 3729
rect 43551 3689 43563 3723
rect 43597 3720 43609 3723
rect 44910 3720 44916 3732
rect 43597 3692 44916 3720
rect 43597 3689 43609 3692
rect 43551 3683 43609 3689
rect 44910 3680 44916 3692
rect 44968 3680 44974 3732
rect 45554 3680 45560 3732
rect 45612 3680 45618 3732
rect 46750 3680 46756 3732
rect 46808 3720 46814 3732
rect 47397 3723 47455 3729
rect 47397 3720 47409 3723
rect 46808 3692 47409 3720
rect 46808 3680 46814 3692
rect 47397 3689 47409 3692
rect 47443 3689 47455 3723
rect 47397 3683 47455 3689
rect 48038 3680 48044 3732
rect 48096 3720 48102 3732
rect 49605 3723 49663 3729
rect 49605 3720 49617 3723
rect 48096 3692 49617 3720
rect 48096 3680 48102 3692
rect 49605 3689 49617 3692
rect 49651 3689 49663 3723
rect 49605 3683 49663 3689
rect 53190 3680 53196 3732
rect 53248 3680 53254 3732
rect 68646 3680 68652 3732
rect 68704 3680 68710 3732
rect 71682 3680 71688 3732
rect 71740 3680 71746 3732
rect 77570 3680 77576 3732
rect 77628 3680 77634 3732
rect 42061 3655 42119 3661
rect 37200 3624 38700 3652
rect 35253 3587 35311 3593
rect 35253 3584 35265 3587
rect 33652 3556 35265 3584
rect 33652 3544 33658 3556
rect 35253 3553 35265 3556
rect 35299 3553 35311 3587
rect 37200 3584 37228 3624
rect 35253 3547 35311 3553
rect 35544 3556 37228 3584
rect 28368 3488 28672 3516
rect 28718 3476 28724 3528
rect 28776 3476 28782 3528
rect 29086 3476 29092 3528
rect 29144 3476 29150 3528
rect 31110 3516 31116 3528
rect 30300 3488 31116 3516
rect 30300 3448 30328 3488
rect 31110 3476 31116 3488
rect 31168 3476 31174 3528
rect 31662 3476 31668 3528
rect 31720 3476 31726 3528
rect 32217 3519 32275 3525
rect 32217 3485 32229 3519
rect 32263 3516 32275 3519
rect 32263 3488 32352 3516
rect 32263 3485 32275 3488
rect 32217 3479 32275 3485
rect 28276 3420 30328 3448
rect 30374 3408 30380 3460
rect 30432 3448 30438 3460
rect 30653 3451 30711 3457
rect 30653 3448 30665 3451
rect 30432 3420 30665 3448
rect 30432 3408 30438 3420
rect 30653 3417 30665 3420
rect 30699 3417 30711 3451
rect 30653 3411 30711 3417
rect 18046 3380 18052 3392
rect 16408 3352 18052 3380
rect 18046 3340 18052 3352
rect 18104 3380 18110 3392
rect 18598 3380 18604 3392
rect 18104 3352 18604 3380
rect 18104 3340 18110 3352
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 19306 3352 19340 3392
rect 19334 3340 19340 3352
rect 19392 3380 19398 3392
rect 20806 3380 20812 3392
rect 19392 3352 20812 3380
rect 19392 3340 19398 3352
rect 20806 3340 20812 3352
rect 20864 3340 20870 3392
rect 21450 3340 21456 3392
rect 21508 3380 21514 3392
rect 21821 3383 21879 3389
rect 21821 3380 21833 3383
rect 21508 3352 21833 3380
rect 21508 3340 21514 3352
rect 21821 3349 21833 3352
rect 21867 3349 21879 3383
rect 21821 3343 21879 3349
rect 24210 3340 24216 3392
rect 24268 3380 24274 3392
rect 24762 3380 24768 3392
rect 24268 3352 24768 3380
rect 24268 3340 24274 3352
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 25406 3340 25412 3392
rect 25464 3340 25470 3392
rect 25682 3340 25688 3392
rect 25740 3340 25746 3392
rect 26234 3340 26240 3392
rect 26292 3380 26298 3392
rect 28629 3383 28687 3389
rect 28629 3380 28641 3383
rect 26292 3352 28641 3380
rect 26292 3340 26298 3352
rect 28629 3349 28641 3352
rect 28675 3349 28687 3383
rect 28629 3343 28687 3349
rect 29454 3340 29460 3392
rect 29512 3380 29518 3392
rect 30834 3380 30840 3392
rect 29512 3352 30840 3380
rect 29512 3340 29518 3352
rect 30834 3340 30840 3352
rect 30892 3340 30898 3392
rect 32324 3380 32352 3488
rect 34146 3476 34152 3528
rect 34204 3476 34210 3528
rect 34425 3519 34483 3525
rect 34425 3485 34437 3519
rect 34471 3516 34483 3519
rect 34882 3516 34888 3528
rect 34471 3488 34888 3516
rect 34471 3485 34483 3488
rect 34425 3479 34483 3485
rect 34882 3476 34888 3488
rect 34940 3516 34946 3528
rect 35544 3516 35572 3556
rect 34940 3488 35572 3516
rect 35621 3519 35679 3525
rect 34940 3476 34946 3488
rect 35621 3485 35633 3519
rect 35667 3485 35679 3519
rect 35621 3479 35679 3485
rect 32585 3451 32643 3457
rect 32585 3417 32597 3451
rect 32631 3448 32643 3451
rect 32674 3448 32680 3460
rect 32631 3420 32680 3448
rect 32631 3417 32643 3420
rect 32585 3411 32643 3417
rect 32674 3408 32680 3420
rect 32732 3408 32738 3460
rect 33042 3408 33048 3460
rect 33100 3408 33106 3460
rect 33870 3408 33876 3460
rect 33928 3448 33934 3460
rect 34241 3451 34299 3457
rect 34241 3448 34253 3451
rect 33928 3420 34253 3448
rect 33928 3408 33934 3420
rect 34241 3417 34253 3420
rect 34287 3448 34299 3451
rect 35636 3448 35664 3479
rect 35710 3476 35716 3528
rect 35768 3476 35774 3528
rect 35912 3525 35940 3556
rect 38562 3544 38568 3596
rect 38620 3544 38626 3596
rect 38672 3584 38700 3624
rect 42061 3621 42073 3655
rect 42107 3652 42119 3655
rect 42518 3652 42524 3664
rect 42107 3624 42524 3652
rect 42107 3621 42119 3624
rect 42061 3615 42119 3621
rect 42518 3612 42524 3624
rect 42576 3612 42582 3664
rect 43806 3612 43812 3664
rect 43864 3652 43870 3664
rect 46661 3655 46719 3661
rect 46661 3652 46673 3655
rect 43864 3624 46673 3652
rect 43864 3612 43870 3624
rect 46661 3621 46673 3624
rect 46707 3621 46719 3655
rect 46661 3615 46719 3621
rect 41690 3584 41696 3596
rect 38672 3556 40908 3584
rect 35897 3519 35955 3525
rect 35897 3485 35909 3519
rect 35943 3485 35955 3519
rect 35897 3479 35955 3485
rect 36081 3519 36139 3525
rect 36081 3485 36093 3519
rect 36127 3516 36139 3519
rect 36262 3516 36268 3528
rect 36127 3488 36268 3516
rect 36127 3485 36139 3488
rect 36081 3479 36139 3485
rect 36262 3476 36268 3488
rect 36320 3476 36326 3528
rect 36357 3519 36415 3525
rect 36357 3485 36369 3519
rect 36403 3516 36415 3519
rect 37182 3516 37188 3528
rect 36403 3488 37188 3516
rect 36403 3485 36415 3488
rect 36357 3479 36415 3485
rect 37182 3476 37188 3488
rect 37240 3476 37246 3528
rect 37274 3476 37280 3528
rect 37332 3476 37338 3528
rect 39114 3476 39120 3528
rect 39172 3476 39178 3528
rect 40586 3476 40592 3528
rect 40644 3476 40650 3528
rect 38470 3448 38476 3460
rect 34287 3420 35572 3448
rect 35636 3420 38476 3448
rect 34287 3417 34299 3420
rect 34241 3411 34299 3417
rect 33502 3380 33508 3392
rect 32324 3352 33508 3380
rect 33502 3340 33508 3352
rect 33560 3340 33566 3392
rect 34146 3340 34152 3392
rect 34204 3380 34210 3392
rect 35069 3383 35127 3389
rect 35069 3380 35081 3383
rect 34204 3352 35081 3380
rect 34204 3340 34210 3352
rect 35069 3349 35081 3352
rect 35115 3349 35127 3383
rect 35069 3343 35127 3349
rect 35158 3340 35164 3392
rect 35216 3340 35222 3392
rect 35544 3380 35572 3420
rect 38470 3408 38476 3420
rect 38528 3408 38534 3460
rect 39390 3408 39396 3460
rect 39448 3408 39454 3460
rect 35710 3380 35716 3392
rect 35544 3352 35716 3380
rect 35710 3340 35716 3352
rect 35768 3340 35774 3392
rect 36078 3340 36084 3392
rect 36136 3380 36142 3392
rect 40678 3380 40684 3392
rect 36136 3352 40684 3380
rect 36136 3340 36142 3352
rect 40678 3340 40684 3352
rect 40736 3340 40742 3392
rect 40770 3340 40776 3392
rect 40828 3340 40834 3392
rect 40880 3380 40908 3556
rect 40972 3556 41696 3584
rect 40972 3525 41000 3556
rect 41690 3544 41696 3556
rect 41748 3544 41754 3596
rect 42242 3544 42248 3596
rect 42300 3584 42306 3596
rect 45925 3587 45983 3593
rect 45925 3584 45937 3587
rect 42300 3556 45937 3584
rect 42300 3544 42306 3556
rect 45925 3553 45937 3556
rect 45971 3553 45983 3587
rect 45925 3547 45983 3553
rect 46842 3544 46848 3596
rect 46900 3584 46906 3596
rect 47213 3587 47271 3593
rect 47213 3584 47225 3587
rect 46900 3556 47225 3584
rect 46900 3544 46906 3556
rect 47213 3553 47225 3556
rect 47259 3553 47271 3587
rect 47213 3547 47271 3553
rect 47854 3544 47860 3596
rect 47912 3584 47918 3596
rect 48685 3587 48743 3593
rect 48685 3584 48697 3587
rect 47912 3556 48697 3584
rect 47912 3544 47918 3556
rect 48685 3553 48697 3556
rect 48731 3553 48743 3587
rect 48685 3547 48743 3553
rect 48866 3544 48872 3596
rect 48924 3544 48930 3596
rect 52365 3587 52423 3593
rect 52365 3553 52377 3587
rect 52411 3584 52423 3587
rect 53837 3587 53895 3593
rect 53837 3584 53849 3587
rect 52411 3556 53849 3584
rect 52411 3553 52423 3556
rect 52365 3547 52423 3553
rect 53837 3553 53849 3556
rect 53883 3553 53895 3587
rect 53837 3547 53895 3553
rect 54018 3544 54024 3596
rect 54076 3544 54082 3596
rect 67821 3587 67879 3593
rect 67821 3553 67833 3587
rect 67867 3584 67879 3587
rect 69201 3587 69259 3593
rect 69201 3584 69213 3587
rect 67867 3556 69213 3584
rect 67867 3553 67879 3556
rect 67821 3547 67879 3553
rect 69201 3553 69213 3556
rect 69247 3553 69259 3587
rect 69201 3547 69259 3553
rect 69474 3544 69480 3596
rect 69532 3544 69538 3596
rect 73706 3544 73712 3596
rect 73764 3544 73770 3596
rect 77018 3544 77024 3596
rect 77076 3544 77082 3596
rect 40957 3519 41015 3525
rect 40957 3485 40969 3519
rect 41003 3485 41015 3519
rect 40957 3479 41015 3485
rect 41046 3476 41052 3528
rect 41104 3476 41110 3528
rect 41230 3476 41236 3528
rect 41288 3476 41294 3528
rect 41322 3476 41328 3528
rect 41380 3476 41386 3528
rect 43809 3519 43867 3525
rect 43809 3485 43821 3519
rect 43855 3485 43867 3519
rect 43809 3479 43867 3485
rect 42518 3408 42524 3460
rect 42576 3408 42582 3460
rect 43254 3380 43260 3392
rect 40880 3352 43260 3380
rect 43254 3340 43260 3352
rect 43312 3340 43318 3392
rect 43346 3340 43352 3392
rect 43404 3380 43410 3392
rect 43824 3380 43852 3479
rect 43898 3476 43904 3528
rect 43956 3476 43962 3528
rect 45373 3519 45431 3525
rect 45373 3485 45385 3519
rect 45419 3485 45431 3519
rect 45373 3479 45431 3485
rect 46569 3519 46627 3525
rect 46569 3485 46581 3519
rect 46615 3516 46627 3519
rect 47118 3516 47124 3528
rect 46615 3488 47124 3516
rect 46615 3485 46627 3488
rect 46569 3479 46627 3485
rect 45097 3451 45155 3457
rect 45097 3417 45109 3451
rect 45143 3448 45155 3451
rect 45186 3448 45192 3460
rect 45143 3420 45192 3448
rect 45143 3417 45155 3420
rect 45097 3411 45155 3417
rect 45186 3408 45192 3420
rect 45244 3408 45250 3460
rect 45388 3448 45416 3479
rect 47118 3476 47124 3488
rect 47176 3476 47182 3528
rect 47946 3476 47952 3528
rect 48004 3476 48010 3528
rect 50249 3519 50307 3525
rect 50249 3485 50261 3519
rect 50295 3516 50307 3519
rect 50798 3516 50804 3528
rect 50295 3488 50804 3516
rect 50295 3485 50307 3488
rect 50249 3479 50307 3485
rect 50798 3476 50804 3488
rect 50856 3476 50862 3528
rect 51813 3519 51871 3525
rect 51813 3485 51825 3519
rect 51859 3516 51871 3519
rect 52457 3519 52515 3525
rect 52457 3516 52469 3519
rect 51859 3488 52469 3516
rect 51859 3485 51871 3488
rect 51813 3479 51871 3485
rect 52457 3485 52469 3488
rect 52503 3485 52515 3519
rect 52457 3479 52515 3485
rect 53006 3476 53012 3528
rect 53064 3476 53070 3528
rect 54573 3519 54631 3525
rect 54573 3485 54585 3519
rect 54619 3516 54631 3519
rect 54665 3519 54723 3525
rect 54665 3516 54677 3519
rect 54619 3488 54677 3516
rect 54619 3485 54631 3488
rect 54573 3479 54631 3485
rect 54665 3485 54677 3488
rect 54711 3485 54723 3519
rect 54665 3479 54723 3485
rect 58069 3519 58127 3525
rect 58069 3485 58081 3519
rect 58115 3516 58127 3519
rect 58161 3519 58219 3525
rect 58161 3516 58173 3519
rect 58115 3488 58173 3516
rect 58115 3485 58127 3488
rect 58069 3479 58127 3485
rect 58161 3485 58173 3488
rect 58207 3485 58219 3519
rect 58161 3479 58219 3485
rect 58713 3519 58771 3525
rect 58713 3485 58725 3519
rect 58759 3485 58771 3519
rect 58713 3479 58771 3485
rect 49513 3451 49571 3457
rect 45388 3420 49464 3448
rect 43404 3352 43852 3380
rect 43404 3340 43410 3352
rect 48130 3340 48136 3392
rect 48188 3340 48194 3392
rect 49436 3380 49464 3420
rect 49513 3417 49525 3451
rect 49559 3448 49571 3451
rect 50522 3448 50528 3460
rect 49559 3420 50528 3448
rect 49559 3417 49571 3420
rect 49513 3411 49571 3417
rect 50522 3408 50528 3420
rect 50580 3408 50586 3460
rect 57330 3408 57336 3460
rect 57388 3448 57394 3460
rect 58728 3448 58756 3479
rect 59446 3476 59452 3528
rect 59504 3476 59510 3528
rect 62025 3519 62083 3525
rect 62025 3485 62037 3519
rect 62071 3516 62083 3519
rect 62117 3519 62175 3525
rect 62117 3516 62129 3519
rect 62071 3488 62129 3516
rect 62071 3485 62083 3488
rect 62025 3479 62083 3485
rect 62117 3485 62129 3488
rect 62163 3485 62175 3519
rect 62117 3479 62175 3485
rect 62669 3519 62727 3525
rect 62669 3485 62681 3519
rect 62715 3485 62727 3519
rect 62669 3479 62727 3485
rect 57388 3420 58756 3448
rect 57388 3408 57394 3420
rect 60918 3408 60924 3460
rect 60976 3448 60982 3460
rect 62684 3448 62712 3479
rect 63402 3476 63408 3528
rect 63460 3476 63466 3528
rect 64506 3476 64512 3528
rect 64564 3476 64570 3528
rect 65061 3519 65119 3525
rect 65061 3485 65073 3519
rect 65107 3516 65119 3519
rect 65705 3519 65763 3525
rect 65705 3516 65717 3519
rect 65107 3488 65717 3516
rect 65107 3485 65119 3488
rect 65061 3479 65119 3485
rect 65705 3485 65717 3488
rect 65751 3485 65763 3519
rect 65705 3479 65763 3485
rect 67269 3519 67327 3525
rect 67269 3485 67281 3519
rect 67315 3516 67327 3519
rect 67913 3519 67971 3525
rect 67913 3516 67925 3519
rect 67315 3488 67925 3516
rect 67315 3485 67327 3488
rect 67269 3479 67327 3485
rect 67913 3485 67925 3488
rect 67959 3485 67971 3519
rect 67913 3479 67971 3485
rect 68462 3476 68468 3528
rect 68520 3476 68526 3528
rect 70029 3519 70087 3525
rect 70029 3485 70041 3519
rect 70075 3516 70087 3519
rect 70121 3519 70179 3525
rect 70121 3516 70133 3519
rect 70075 3488 70133 3516
rect 70075 3485 70087 3488
rect 70029 3479 70087 3485
rect 70121 3485 70133 3488
rect 70167 3485 70179 3519
rect 70121 3479 70179 3485
rect 72329 3519 72387 3525
rect 72329 3485 72341 3519
rect 72375 3516 72387 3519
rect 72421 3519 72479 3525
rect 72421 3516 72433 3519
rect 72375 3488 72433 3516
rect 72375 3485 72387 3488
rect 72329 3479 72387 3485
rect 72421 3485 72433 3488
rect 72467 3485 72479 3519
rect 72421 3479 72479 3485
rect 72970 3476 72976 3528
rect 73028 3476 73034 3528
rect 74442 3476 74448 3528
rect 74500 3516 74506 3528
rect 75089 3519 75147 3525
rect 75089 3516 75101 3519
rect 74500 3488 75101 3516
rect 74500 3476 74506 3488
rect 75089 3485 75101 3488
rect 75135 3485 75147 3519
rect 75089 3479 75147 3485
rect 76650 3476 76656 3528
rect 76708 3476 76714 3528
rect 60976 3420 62712 3448
rect 60976 3408 60982 3420
rect 75454 3408 75460 3460
rect 75512 3408 75518 3460
rect 49970 3380 49976 3392
rect 49436 3352 49976 3380
rect 49970 3340 49976 3352
rect 50028 3340 50034 3392
rect 55309 3383 55367 3389
rect 55309 3349 55321 3383
rect 55355 3380 55367 3383
rect 56042 3380 56048 3392
rect 55355 3352 56048 3380
rect 55355 3349 55367 3352
rect 55309 3343 55367 3349
rect 56042 3340 56048 3352
rect 56100 3340 56106 3392
rect 57422 3340 57428 3392
rect 57480 3340 57486 3392
rect 58618 3340 58624 3392
rect 58676 3380 58682 3392
rect 58897 3383 58955 3389
rect 58897 3380 58909 3383
rect 58676 3352 58909 3380
rect 58676 3340 58682 3352
rect 58897 3349 58909 3352
rect 58943 3349 58955 3383
rect 58897 3343 58955 3349
rect 61102 3340 61108 3392
rect 61160 3380 61166 3392
rect 61381 3383 61439 3389
rect 61381 3380 61393 3383
rect 61160 3352 61393 3380
rect 61160 3340 61166 3352
rect 61381 3349 61393 3352
rect 61427 3349 61439 3383
rect 61381 3343 61439 3349
rect 62758 3340 62764 3392
rect 62816 3380 62822 3392
rect 62853 3383 62911 3389
rect 62853 3380 62865 3383
rect 62816 3352 62865 3380
rect 62816 3340 62822 3352
rect 62853 3349 62865 3352
rect 62899 3349 62911 3383
rect 62853 3343 62911 3349
rect 64874 3340 64880 3392
rect 64932 3380 64938 3392
rect 65153 3383 65211 3389
rect 65153 3380 65165 3383
rect 64932 3352 65165 3380
rect 64932 3340 64938 3352
rect 65153 3349 65165 3352
rect 65199 3349 65211 3383
rect 65153 3343 65211 3349
rect 70765 3383 70823 3389
rect 70765 3349 70777 3383
rect 70811 3380 70823 3383
rect 71498 3380 71504 3392
rect 70811 3352 71504 3380
rect 70811 3349 70823 3352
rect 70765 3343 70823 3349
rect 71498 3340 71504 3352
rect 71556 3340 71562 3392
rect 73157 3383 73215 3389
rect 73157 3349 73169 3383
rect 73203 3380 73215 3383
rect 73246 3380 73252 3392
rect 73203 3352 73252 3380
rect 73203 3349 73215 3352
rect 73157 3343 73215 3349
rect 73246 3340 73252 3352
rect 73304 3340 73310 3392
rect 74534 3340 74540 3392
rect 74592 3340 74598 3392
rect 2024 3290 77924 3312
rect 2024 3238 5794 3290
rect 5846 3238 5858 3290
rect 5910 3238 5922 3290
rect 5974 3238 5986 3290
rect 6038 3238 6050 3290
rect 6102 3238 36514 3290
rect 36566 3238 36578 3290
rect 36630 3238 36642 3290
rect 36694 3238 36706 3290
rect 36758 3238 36770 3290
rect 36822 3238 67234 3290
rect 67286 3238 67298 3290
rect 67350 3238 67362 3290
rect 67414 3238 67426 3290
rect 67478 3238 67490 3290
rect 67542 3238 77924 3290
rect 2024 3216 77924 3238
rect 3786 3136 3792 3188
rect 3844 3136 3850 3188
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 7285 3179 7343 3185
rect 7285 3176 7297 3179
rect 5316 3148 7297 3176
rect 5316 3136 5322 3148
rect 7285 3145 7297 3148
rect 7331 3145 7343 3179
rect 7285 3139 7343 3145
rect 8202 3136 8208 3188
rect 8260 3136 8266 3188
rect 8941 3179 8999 3185
rect 8941 3145 8953 3179
rect 8987 3176 8999 3179
rect 9214 3176 9220 3188
rect 8987 3148 9220 3176
rect 8987 3145 8999 3148
rect 8941 3139 8999 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9677 3179 9735 3185
rect 9677 3145 9689 3179
rect 9723 3176 9735 3179
rect 9950 3176 9956 3188
rect 9723 3148 9956 3176
rect 9723 3145 9735 3148
rect 9677 3139 9735 3145
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 10410 3136 10416 3188
rect 10468 3176 10474 3188
rect 10468 3148 12112 3176
rect 10468 3136 10474 3148
rect 10134 3108 10140 3120
rect 3252 3080 10140 3108
rect 3252 3049 3280 3080
rect 10134 3068 10140 3080
rect 10192 3068 10198 3120
rect 10778 3068 10784 3120
rect 10836 3068 10842 3120
rect 11238 3068 11244 3120
rect 11296 3068 11302 3120
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3040 4951 3043
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 4939 3012 7481 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 7558 3000 7564 3052
rect 7616 3000 7622 3052
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 9769 3043 9827 3049
rect 9769 3040 9781 3043
rect 8536 3012 9781 3040
rect 8536 3000 8542 3012
rect 9769 3009 9781 3012
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 9950 3000 9956 3052
rect 10008 3040 10014 3052
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 10008 3012 10425 3040
rect 10008 3000 10014 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 10502 3000 10508 3052
rect 10560 3000 10566 3052
rect 12084 3040 12112 3148
rect 12158 3136 12164 3188
rect 12216 3176 12222 3188
rect 12253 3179 12311 3185
rect 12253 3176 12265 3179
rect 12216 3148 12265 3176
rect 12216 3136 12222 3148
rect 12253 3145 12265 3148
rect 12299 3145 12311 3179
rect 12253 3139 12311 3145
rect 12342 3136 12348 3188
rect 12400 3176 12406 3188
rect 12897 3179 12955 3185
rect 12400 3148 12848 3176
rect 12400 3136 12406 3148
rect 12618 3068 12624 3120
rect 12676 3068 12682 3120
rect 12820 3108 12848 3148
rect 12897 3145 12909 3179
rect 12943 3176 12955 3179
rect 12986 3176 12992 3188
rect 12943 3148 12992 3176
rect 12943 3145 12955 3148
rect 12897 3139 12955 3145
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 14918 3176 14924 3188
rect 13136 3148 14924 3176
rect 13136 3136 13142 3148
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 15930 3136 15936 3188
rect 15988 3176 15994 3188
rect 16850 3176 16856 3188
rect 15988 3148 16856 3176
rect 15988 3136 15994 3148
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17310 3136 17316 3188
rect 17368 3176 17374 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17368 3148 17417 3176
rect 17368 3136 17374 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17405 3139 17463 3145
rect 17586 3136 17592 3188
rect 17644 3136 17650 3188
rect 18598 3136 18604 3188
rect 18656 3176 18662 3188
rect 18656 3148 19932 3176
rect 18656 3136 18662 3148
rect 13814 3108 13820 3120
rect 12820 3080 13820 3108
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 12084 3012 12296 3040
rect 4341 2975 4399 2981
rect 4341 2941 4353 2975
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 5077 2975 5135 2981
rect 5077 2941 5089 2975
rect 5123 2972 5135 2975
rect 5534 2972 5540 2984
rect 5123 2944 5540 2972
rect 5123 2941 5135 2944
rect 5077 2935 5135 2941
rect 4356 2904 4384 2935
rect 5534 2932 5540 2944
rect 5592 2932 5598 2984
rect 5626 2932 5632 2984
rect 5684 2932 5690 2984
rect 5718 2932 5724 2984
rect 5776 2932 5782 2984
rect 6914 2972 6920 2984
rect 5828 2944 6920 2972
rect 5828 2904 5856 2944
rect 6914 2932 6920 2944
rect 6972 2932 6978 2984
rect 7098 2932 7104 2984
rect 7156 2932 7162 2984
rect 7650 2932 7656 2984
rect 7708 2972 7714 2984
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 7708 2944 8309 2972
rect 7708 2932 7714 2944
rect 8297 2941 8309 2944
rect 8343 2941 8355 2975
rect 8297 2935 8355 2941
rect 9122 2932 9128 2984
rect 9180 2932 9186 2984
rect 12268 2972 12296 3012
rect 13078 3000 13084 3052
rect 13136 3000 13142 3052
rect 14936 3049 14964 3136
rect 15102 3068 15108 3120
rect 15160 3108 15166 3120
rect 15160 3080 15686 3108
rect 15160 3068 15166 3080
rect 14921 3043 14979 3049
rect 14921 3009 14933 3043
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3040 16911 3043
rect 17604 3040 17632 3136
rect 17954 3068 17960 3120
rect 18012 3108 18018 3120
rect 18325 3111 18383 3117
rect 18325 3108 18337 3111
rect 18012 3080 18337 3108
rect 18012 3068 18018 3080
rect 18325 3077 18337 3080
rect 18371 3077 18383 3111
rect 18325 3071 18383 3077
rect 19334 3068 19340 3120
rect 19392 3068 19398 3120
rect 16899 3012 17632 3040
rect 16899 3009 16911 3012
rect 16853 3003 16911 3009
rect 18046 3000 18052 3052
rect 18104 3000 18110 3052
rect 13357 2975 13415 2981
rect 13357 2972 13369 2975
rect 9646 2944 11836 2972
rect 12268 2944 13369 2972
rect 4356 2876 5856 2904
rect 6365 2907 6423 2913
rect 6365 2873 6377 2907
rect 6411 2904 6423 2907
rect 9646 2904 9674 2944
rect 6411 2876 9674 2904
rect 11808 2904 11836 2944
rect 13357 2941 13369 2944
rect 13403 2941 13415 2975
rect 15197 2975 15255 2981
rect 15197 2972 15209 2975
rect 13357 2935 13415 2941
rect 14384 2944 15209 2972
rect 11808 2876 12434 2904
rect 6411 2873 6423 2876
rect 6365 2867 6423 2873
rect 6454 2796 6460 2848
rect 6512 2796 6518 2848
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 12250 2836 12256 2848
rect 10192 2808 12256 2836
rect 10192 2796 10198 2808
rect 12250 2796 12256 2808
rect 12308 2796 12314 2848
rect 12406 2836 12434 2876
rect 14384 2836 14412 2944
rect 15197 2941 15209 2944
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 16669 2975 16727 2981
rect 16669 2972 16681 2975
rect 15620 2944 16681 2972
rect 15620 2932 15626 2944
rect 16669 2941 16681 2944
rect 16715 2941 16727 2975
rect 16669 2935 16727 2941
rect 17310 2932 17316 2984
rect 17368 2972 17374 2984
rect 19352 2972 19380 3068
rect 19904 3049 19932 3148
rect 21082 3136 21088 3188
rect 21140 3176 21146 3188
rect 21637 3179 21695 3185
rect 21637 3176 21649 3179
rect 21140 3148 21649 3176
rect 21140 3136 21146 3148
rect 21637 3145 21649 3148
rect 21683 3145 21695 3179
rect 21637 3139 21695 3145
rect 22557 3179 22615 3185
rect 22557 3145 22569 3179
rect 22603 3176 22615 3179
rect 22646 3176 22652 3188
rect 22603 3148 22652 3176
rect 22603 3145 22615 3148
rect 22557 3139 22615 3145
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 23014 3136 23020 3188
rect 23072 3136 23078 3188
rect 25041 3179 25099 3185
rect 23216 3148 24900 3176
rect 21390 3080 22692 3108
rect 19889 3043 19947 3049
rect 19889 3009 19901 3043
rect 19935 3009 19947 3043
rect 19889 3003 19947 3009
rect 21818 3000 21824 3052
rect 21876 3040 21882 3052
rect 21913 3043 21971 3049
rect 21913 3040 21925 3043
rect 21876 3012 21925 3040
rect 21876 3000 21882 3012
rect 21913 3009 21925 3012
rect 21959 3040 21971 3043
rect 22002 3040 22008 3052
rect 21959 3012 22008 3040
rect 21959 3009 21971 3012
rect 21913 3003 21971 3009
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 17368 2944 19380 2972
rect 17368 2932 17374 2944
rect 19702 2932 19708 2984
rect 19760 2972 19766 2984
rect 20165 2975 20223 2981
rect 20165 2972 20177 2975
rect 19760 2944 20177 2972
rect 19760 2932 19766 2944
rect 20165 2941 20177 2944
rect 20211 2941 20223 2975
rect 22664 2972 22692 3080
rect 22741 3043 22799 3049
rect 22741 3009 22753 3043
rect 22787 3040 22799 3043
rect 23216 3040 23244 3148
rect 24486 3068 24492 3120
rect 24544 3068 24550 3120
rect 24872 3108 24900 3148
rect 25041 3145 25053 3179
rect 25087 3176 25099 3179
rect 25958 3176 25964 3188
rect 25087 3148 25964 3176
rect 25087 3145 25099 3148
rect 25041 3139 25099 3145
rect 25958 3136 25964 3148
rect 26016 3136 26022 3188
rect 26970 3136 26976 3188
rect 27028 3136 27034 3188
rect 27430 3136 27436 3188
rect 27488 3136 27494 3188
rect 27525 3179 27583 3185
rect 27525 3145 27537 3179
rect 27571 3176 27583 3179
rect 28442 3176 28448 3188
rect 27571 3148 28448 3176
rect 27571 3145 27583 3148
rect 27525 3139 27583 3145
rect 28442 3136 28448 3148
rect 28500 3136 28506 3188
rect 28534 3136 28540 3188
rect 28592 3136 28598 3188
rect 30742 3176 30748 3188
rect 28736 3148 30748 3176
rect 28736 3120 28764 3148
rect 30742 3136 30748 3148
rect 30800 3136 30806 3188
rect 30834 3136 30840 3188
rect 30892 3176 30898 3188
rect 33505 3179 33563 3185
rect 33505 3176 33517 3179
rect 30892 3148 33517 3176
rect 30892 3136 30898 3148
rect 33505 3145 33517 3148
rect 33551 3145 33563 3179
rect 33505 3139 33563 3145
rect 34057 3179 34115 3185
rect 34057 3145 34069 3179
rect 34103 3176 34115 3179
rect 36078 3176 36084 3188
rect 34103 3148 36084 3176
rect 34103 3145 34115 3148
rect 34057 3139 34115 3145
rect 36078 3136 36084 3148
rect 36136 3136 36142 3188
rect 37918 3176 37924 3188
rect 36188 3148 37924 3176
rect 25409 3111 25467 3117
rect 24872 3080 25360 3108
rect 22787 3012 23244 3040
rect 22787 3009 22799 3012
rect 22741 3003 22799 3009
rect 23382 3000 23388 3052
rect 23440 3000 23446 3052
rect 24762 3000 24768 3052
rect 24820 3000 24826 3052
rect 24854 3000 24860 3052
rect 24912 3000 24918 3052
rect 25133 3043 25191 3049
rect 25133 3040 25145 3043
rect 24964 3012 25145 3040
rect 23400 2972 23428 3000
rect 22664 2944 23428 2972
rect 20165 2935 20223 2941
rect 23750 2932 23756 2984
rect 23808 2972 23814 2984
rect 24964 2972 24992 3012
rect 25133 3009 25145 3012
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 25222 3000 25228 3052
rect 25280 3000 25286 3052
rect 25332 3040 25360 3080
rect 25409 3077 25421 3111
rect 25455 3108 25467 3111
rect 25498 3108 25504 3120
rect 25455 3080 25504 3108
rect 25455 3077 25467 3080
rect 25409 3071 25467 3077
rect 25498 3068 25504 3080
rect 25556 3108 25562 3120
rect 26050 3108 26056 3120
rect 25556 3080 26056 3108
rect 25556 3068 25562 3080
rect 26050 3068 26056 3080
rect 26108 3068 26114 3120
rect 28718 3068 28724 3120
rect 28776 3068 28782 3120
rect 29546 3068 29552 3120
rect 29604 3068 29610 3120
rect 30006 3068 30012 3120
rect 30064 3068 30070 3120
rect 30098 3068 30104 3120
rect 30156 3108 30162 3120
rect 30469 3111 30527 3117
rect 30156 3080 30420 3108
rect 30156 3068 30162 3080
rect 26694 3040 26700 3052
rect 25332 3012 26700 3040
rect 26694 3000 26700 3012
rect 26752 3000 26758 3052
rect 26878 3000 26884 3052
rect 26936 3000 26942 3052
rect 27338 3000 27344 3052
rect 27396 3000 27402 3052
rect 27982 3000 27988 3052
rect 28040 3000 28046 3052
rect 30392 3049 30420 3080
rect 30469 3077 30481 3111
rect 30515 3108 30527 3111
rect 30558 3108 30564 3120
rect 30515 3080 30564 3108
rect 30515 3077 30527 3080
rect 30469 3071 30527 3077
rect 30558 3068 30564 3080
rect 30616 3068 30622 3120
rect 30926 3108 30932 3120
rect 30668 3080 30932 3108
rect 30668 3049 30696 3080
rect 30926 3068 30932 3080
rect 30984 3068 30990 3120
rect 32306 3068 32312 3120
rect 32364 3108 32370 3120
rect 32401 3111 32459 3117
rect 32401 3108 32413 3111
rect 32364 3080 32413 3108
rect 32364 3068 32370 3080
rect 32401 3077 32413 3080
rect 32447 3077 32459 3111
rect 32401 3071 32459 3077
rect 32766 3068 32772 3120
rect 32824 3108 32830 3120
rect 33413 3111 33471 3117
rect 32824 3080 33364 3108
rect 32824 3068 32830 3080
rect 28169 3043 28227 3049
rect 28169 3009 28181 3043
rect 28215 3040 28227 3043
rect 30377 3043 30435 3049
rect 28215 3012 28856 3040
rect 28215 3009 28227 3012
rect 28169 3003 28227 3009
rect 23808 2944 24992 2972
rect 23808 2932 23814 2944
rect 26418 2932 26424 2984
rect 26476 2932 26482 2984
rect 26786 2932 26792 2984
rect 26844 2972 26850 2984
rect 28077 2975 28135 2981
rect 28077 2972 28089 2975
rect 26844 2944 28089 2972
rect 26844 2932 26850 2944
rect 28077 2941 28089 2944
rect 28123 2941 28135 2975
rect 28077 2935 28135 2941
rect 28261 2975 28319 2981
rect 28261 2941 28273 2975
rect 28307 2972 28319 2975
rect 28626 2972 28632 2984
rect 28307 2944 28632 2972
rect 28307 2941 28319 2944
rect 28261 2935 28319 2941
rect 28626 2932 28632 2944
rect 28684 2932 28690 2984
rect 28828 2972 28856 3012
rect 30377 3009 30389 3043
rect 30423 3009 30435 3043
rect 30377 3003 30435 3009
rect 30653 3043 30711 3049
rect 30653 3009 30665 3043
rect 30699 3009 30711 3043
rect 30653 3003 30711 3009
rect 30837 3043 30895 3049
rect 30837 3009 30849 3043
rect 30883 3040 30895 3043
rect 31018 3040 31024 3052
rect 30883 3012 31024 3040
rect 30883 3009 30895 3012
rect 30837 3003 30895 3009
rect 31018 3000 31024 3012
rect 31076 3000 31082 3052
rect 31294 3000 31300 3052
rect 31352 3000 31358 3052
rect 32674 3000 32680 3052
rect 32732 3000 32738 3052
rect 33336 3040 33364 3080
rect 33413 3077 33425 3111
rect 33459 3108 33471 3111
rect 33962 3108 33968 3120
rect 33459 3080 33968 3108
rect 33459 3077 33471 3080
rect 33413 3071 33471 3077
rect 33962 3068 33968 3080
rect 34020 3068 34026 3120
rect 35526 3108 35532 3120
rect 35190 3080 35532 3108
rect 35526 3068 35532 3080
rect 35584 3068 35590 3120
rect 35618 3068 35624 3120
rect 35676 3068 35682 3120
rect 33870 3040 33876 3052
rect 33336 3012 33876 3040
rect 33870 3000 33876 3012
rect 33928 3000 33934 3052
rect 36188 3049 36216 3148
rect 37918 3136 37924 3148
rect 37976 3176 37982 3188
rect 37976 3148 41414 3176
rect 37976 3136 37982 3148
rect 38396 3049 38424 3148
rect 38654 3068 38660 3120
rect 38712 3068 38718 3120
rect 41386 3108 41414 3148
rect 42058 3136 42064 3188
rect 42116 3136 42122 3188
rect 42705 3179 42763 3185
rect 42705 3145 42717 3179
rect 42751 3176 42763 3179
rect 42978 3176 42984 3188
rect 42751 3148 42984 3176
rect 42751 3145 42763 3148
rect 42705 3139 42763 3145
rect 42978 3136 42984 3148
rect 43036 3136 43042 3188
rect 43165 3179 43223 3185
rect 43165 3145 43177 3179
rect 43211 3176 43223 3179
rect 44358 3176 44364 3188
rect 43211 3148 44364 3176
rect 43211 3145 43223 3148
rect 43165 3139 43223 3145
rect 44358 3136 44364 3148
rect 44416 3136 44422 3188
rect 45097 3179 45155 3185
rect 45097 3145 45109 3179
rect 45143 3176 45155 3179
rect 45278 3176 45284 3188
rect 45143 3148 45284 3176
rect 45143 3145 45155 3148
rect 45097 3139 45155 3145
rect 45278 3136 45284 3148
rect 45336 3136 45342 3188
rect 46934 3136 46940 3188
rect 46992 3176 46998 3188
rect 48133 3179 48191 3185
rect 48133 3176 48145 3179
rect 46992 3148 48145 3176
rect 46992 3136 46998 3148
rect 48133 3145 48145 3148
rect 48179 3145 48191 3179
rect 48133 3139 48191 3145
rect 48314 3136 48320 3188
rect 48372 3176 48378 3188
rect 48372 3148 50200 3176
rect 48372 3136 48378 3148
rect 43625 3111 43683 3117
rect 41386 3080 43392 3108
rect 34057 3043 34115 3049
rect 34057 3009 34069 3043
rect 34103 3009 34115 3043
rect 34057 3003 34115 3009
rect 35897 3043 35955 3049
rect 35897 3009 35909 3043
rect 35943 3040 35955 3043
rect 36173 3043 36231 3049
rect 36173 3040 36185 3043
rect 35943 3012 36185 3040
rect 35943 3009 35955 3012
rect 35897 3003 35955 3009
rect 36173 3009 36185 3012
rect 36219 3009 36231 3043
rect 38381 3043 38439 3049
rect 36173 3003 36231 3009
rect 29914 2972 29920 2984
rect 28828 2944 29920 2972
rect 29914 2932 29920 2944
rect 29972 2932 29978 2984
rect 30296 2975 30354 2981
rect 30296 2941 30308 2975
rect 30342 2972 30354 2975
rect 31202 2972 31208 2984
rect 30342 2944 31208 2972
rect 30342 2941 30354 2944
rect 30296 2935 30354 2941
rect 31202 2932 31208 2944
rect 31260 2932 31266 2984
rect 31846 2932 31852 2984
rect 31904 2972 31910 2984
rect 33594 2972 33600 2984
rect 31904 2944 33600 2972
rect 31904 2932 31910 2944
rect 33594 2932 33600 2944
rect 33652 2932 33658 2984
rect 33778 2932 33784 2984
rect 33836 2972 33842 2984
rect 34072 2972 34100 3003
rect 36449 2975 36507 2981
rect 36449 2972 36461 2975
rect 33836 2944 34100 2972
rect 35820 2944 36461 2972
rect 33836 2932 33842 2944
rect 24854 2864 24860 2916
rect 24912 2904 24918 2916
rect 26510 2904 26516 2916
rect 24912 2876 26516 2904
rect 24912 2864 24918 2876
rect 26510 2864 26516 2876
rect 26568 2864 26574 2916
rect 27157 2907 27215 2913
rect 27157 2873 27169 2907
rect 27203 2873 27215 2907
rect 27157 2867 27215 2873
rect 28445 2907 28503 2913
rect 28445 2873 28457 2907
rect 28491 2904 28503 2907
rect 28994 2904 29000 2916
rect 28491 2876 29000 2904
rect 28491 2873 28503 2876
rect 28445 2867 28503 2873
rect 12406 2808 14412 2836
rect 14734 2796 14740 2848
rect 14792 2836 14798 2848
rect 14829 2839 14887 2845
rect 14829 2836 14841 2839
rect 14792 2808 14841 2836
rect 14792 2796 14798 2808
rect 14829 2805 14841 2808
rect 14875 2805 14887 2839
rect 14829 2799 14887 2805
rect 18414 2796 18420 2848
rect 18472 2836 18478 2848
rect 19797 2839 19855 2845
rect 19797 2836 19809 2839
rect 18472 2808 19809 2836
rect 18472 2796 18478 2808
rect 19797 2805 19809 2808
rect 19843 2805 19855 2839
rect 19797 2799 19855 2805
rect 21818 2796 21824 2848
rect 21876 2796 21882 2848
rect 22830 2796 22836 2848
rect 22888 2836 22894 2848
rect 22925 2839 22983 2845
rect 22925 2836 22937 2839
rect 22888 2808 22937 2836
rect 22888 2796 22894 2808
rect 22925 2805 22937 2808
rect 22971 2805 22983 2839
rect 22925 2799 22983 2805
rect 24394 2796 24400 2848
rect 24452 2836 24458 2848
rect 25409 2839 25467 2845
rect 25409 2836 25421 2839
rect 24452 2808 25421 2836
rect 24452 2796 24458 2808
rect 25409 2805 25421 2808
rect 25455 2805 25467 2839
rect 25409 2799 25467 2805
rect 26970 2796 26976 2848
rect 27028 2836 27034 2848
rect 27172 2836 27200 2867
rect 28994 2864 29000 2876
rect 29052 2864 29058 2916
rect 34146 2904 34152 2916
rect 30300 2876 31432 2904
rect 30300 2848 30328 2876
rect 27028 2808 27200 2836
rect 27709 2839 27767 2845
rect 27028 2796 27034 2808
rect 27709 2805 27721 2839
rect 27755 2836 27767 2839
rect 29270 2836 29276 2848
rect 27755 2808 29276 2836
rect 27755 2805 27767 2808
rect 27709 2799 27767 2805
rect 29270 2796 29276 2808
rect 29328 2796 29334 2848
rect 30282 2796 30288 2848
rect 30340 2796 30346 2848
rect 30466 2796 30472 2848
rect 30524 2836 30530 2848
rect 30929 2839 30987 2845
rect 30929 2836 30941 2839
rect 30524 2808 30941 2836
rect 30524 2796 30530 2808
rect 30929 2805 30941 2808
rect 30975 2805 30987 2839
rect 31404 2836 31432 2876
rect 32968 2876 34152 2904
rect 32968 2836 32996 2876
rect 34146 2864 34152 2876
rect 34204 2864 34210 2916
rect 31404 2808 32996 2836
rect 30929 2799 30987 2805
rect 33042 2796 33048 2848
rect 33100 2796 33106 2848
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 35820 2836 35848 2944
rect 36449 2941 36461 2944
rect 36495 2941 36507 2975
rect 37568 2972 37596 3026
rect 38381 3009 38393 3043
rect 38427 3009 38439 3043
rect 38381 3003 38439 3009
rect 39758 3000 39764 3052
rect 39816 3040 39822 3052
rect 41984 3049 42012 3080
rect 43364 3052 43392 3080
rect 43625 3077 43637 3111
rect 43671 3108 43683 3111
rect 43714 3108 43720 3120
rect 43671 3080 43720 3108
rect 43671 3077 43683 3080
rect 43625 3071 43683 3077
rect 43714 3068 43720 3080
rect 43772 3068 43778 3120
rect 44174 3068 44180 3120
rect 44232 3068 44238 3120
rect 50065 3111 50123 3117
rect 50065 3108 50077 3111
rect 48332 3080 50077 3108
rect 41969 3043 42027 3049
rect 39816 3012 40618 3040
rect 39816 3000 39822 3012
rect 41969 3009 41981 3043
rect 42015 3009 42027 3043
rect 41969 3003 42027 3009
rect 42242 3000 42248 3052
rect 42300 3000 42306 3052
rect 42797 3043 42855 3049
rect 42797 3009 42809 3043
rect 42843 3040 42855 3043
rect 42843 3012 43300 3040
rect 42843 3009 42855 3012
rect 42797 3003 42855 3009
rect 39776 2972 39804 3000
rect 37568 2944 39804 2972
rect 40221 2975 40279 2981
rect 36449 2935 36507 2941
rect 37458 2864 37464 2916
rect 37516 2904 37522 2916
rect 37921 2907 37979 2913
rect 37921 2904 37933 2907
rect 37516 2876 37933 2904
rect 37516 2864 37522 2876
rect 37921 2873 37933 2876
rect 37967 2873 37979 2907
rect 37921 2867 37979 2873
rect 34572 2808 35848 2836
rect 34572 2796 34578 2808
rect 35894 2796 35900 2848
rect 35952 2836 35958 2848
rect 38028 2836 38056 2944
rect 40221 2941 40233 2975
rect 40267 2972 40279 2975
rect 41138 2972 41144 2984
rect 40267 2944 41144 2972
rect 40267 2941 40279 2944
rect 40221 2935 40279 2941
rect 41138 2932 41144 2944
rect 41196 2932 41202 2984
rect 41693 2975 41751 2981
rect 41693 2941 41705 2975
rect 41739 2972 41751 2975
rect 42150 2972 42156 2984
rect 41739 2944 42156 2972
rect 41739 2941 41751 2944
rect 41693 2935 41751 2941
rect 42150 2932 42156 2944
rect 42208 2932 42214 2984
rect 42521 2975 42579 2981
rect 42521 2972 42533 2975
rect 42260 2944 42533 2972
rect 40129 2907 40187 2913
rect 40129 2873 40141 2907
rect 40175 2904 40187 2907
rect 40402 2904 40408 2916
rect 40175 2876 40408 2904
rect 40175 2873 40187 2876
rect 40129 2867 40187 2873
rect 40402 2864 40408 2876
rect 40460 2864 40466 2916
rect 35952 2808 38056 2836
rect 35952 2796 35958 2808
rect 40310 2796 40316 2848
rect 40368 2836 40374 2848
rect 42260 2836 42288 2944
rect 42521 2941 42533 2944
rect 42567 2972 42579 2975
rect 43070 2972 43076 2984
rect 42567 2944 43076 2972
rect 42567 2941 42579 2944
rect 42521 2935 42579 2941
rect 43070 2932 43076 2944
rect 43128 2932 43134 2984
rect 40368 2808 42288 2836
rect 43272 2836 43300 3012
rect 43346 3000 43352 3052
rect 43404 3000 43410 3052
rect 45186 3000 45192 3052
rect 45244 3000 45250 3052
rect 46750 3000 46756 3052
rect 46808 3000 46814 3052
rect 48332 3049 48360 3080
rect 50065 3077 50077 3080
rect 50111 3077 50123 3111
rect 50172 3108 50200 3148
rect 50798 3136 50804 3188
rect 50856 3136 50862 3188
rect 51721 3179 51779 3185
rect 51721 3145 51733 3179
rect 51767 3176 51779 3179
rect 53006 3176 53012 3188
rect 51767 3148 53012 3176
rect 51767 3145 51779 3148
rect 51721 3139 51779 3145
rect 53006 3136 53012 3148
rect 53064 3136 53070 3188
rect 53834 3136 53840 3188
rect 53892 3136 53898 3188
rect 57330 3136 57336 3188
rect 57388 3136 57394 3188
rect 58069 3179 58127 3185
rect 58069 3145 58081 3179
rect 58115 3176 58127 3179
rect 59446 3176 59452 3188
rect 58115 3148 59452 3176
rect 58115 3145 58127 3148
rect 58069 3139 58127 3145
rect 59446 3136 59452 3148
rect 59504 3136 59510 3188
rect 60918 3136 60924 3188
rect 60976 3136 60982 3188
rect 61657 3179 61715 3185
rect 61657 3145 61669 3179
rect 61703 3176 61715 3179
rect 63402 3176 63408 3188
rect 61703 3148 63408 3176
rect 61703 3145 61715 3148
rect 61657 3139 61715 3145
rect 63402 3136 63408 3148
rect 63460 3136 63466 3188
rect 64506 3136 64512 3188
rect 64564 3136 64570 3188
rect 65426 3136 65432 3188
rect 65484 3136 65490 3188
rect 67177 3179 67235 3185
rect 67177 3145 67189 3179
rect 67223 3176 67235 3179
rect 68462 3176 68468 3188
rect 67223 3148 68468 3176
rect 67223 3145 67235 3148
rect 67177 3139 67235 3145
rect 68462 3136 68468 3148
rect 68520 3136 68526 3188
rect 69290 3136 69296 3188
rect 69348 3136 69354 3188
rect 74442 3136 74448 3188
rect 74500 3136 74506 3188
rect 70302 3108 70308 3120
rect 50172 3080 70308 3108
rect 50065 3071 50123 3077
rect 48317 3043 48375 3049
rect 48317 3009 48329 3043
rect 48363 3009 48375 3043
rect 48317 3003 48375 3009
rect 49786 3000 49792 3052
rect 49844 3000 49850 3052
rect 51350 3000 51356 3052
rect 51408 3000 51414 3052
rect 51552 3049 51580 3080
rect 51537 3043 51595 3049
rect 51537 3009 51549 3043
rect 51583 3009 51595 3043
rect 51537 3003 51595 3009
rect 52086 3000 52092 3052
rect 52144 3000 52150 3052
rect 53668 3049 53696 3080
rect 53653 3043 53711 3049
rect 53653 3009 53665 3043
rect 53699 3009 53711 3043
rect 53653 3003 53711 3009
rect 54018 3000 54024 3052
rect 54076 3000 54082 3052
rect 56042 3000 56048 3052
rect 56100 3000 56106 3052
rect 57164 3049 57192 3080
rect 57149 3043 57207 3049
rect 57149 3009 57161 3043
rect 57195 3009 57207 3043
rect 57149 3003 57207 3009
rect 57422 3000 57428 3052
rect 57480 3000 57486 3052
rect 60752 3049 60780 3080
rect 60737 3043 60795 3049
rect 60737 3009 60749 3043
rect 60783 3009 60795 3043
rect 60737 3003 60795 3009
rect 61102 3000 61108 3052
rect 61160 3000 61166 3052
rect 61746 3000 61752 3052
rect 61804 3000 61810 3052
rect 64708 3049 64736 3080
rect 64693 3043 64751 3049
rect 64693 3009 64705 3043
rect 64739 3009 64751 3043
rect 64693 3003 64751 3009
rect 64874 3000 64880 3052
rect 64932 3000 64938 3052
rect 65518 3000 65524 3052
rect 65576 3000 65582 3052
rect 67008 3049 67036 3080
rect 66993 3043 67051 3049
rect 66993 3009 67005 3043
rect 67039 3009 67051 3043
rect 66993 3003 67051 3009
rect 67634 3000 67640 3052
rect 67692 3000 67698 3052
rect 69124 3049 69152 3080
rect 70302 3068 70308 3080
rect 70360 3068 70366 3120
rect 69109 3043 69167 3049
rect 69109 3009 69121 3043
rect 69155 3009 69167 3043
rect 69109 3003 69167 3009
rect 69474 3000 69480 3052
rect 69532 3000 69538 3052
rect 71498 3000 71504 3052
rect 71556 3000 71562 3052
rect 72602 3000 72608 3052
rect 72660 3040 72666 3052
rect 72973 3043 73031 3049
rect 72973 3040 72985 3043
rect 72660 3012 72985 3040
rect 72660 3000 72666 3012
rect 72973 3009 72985 3012
rect 73019 3009 73031 3043
rect 72973 3003 73031 3009
rect 74258 3000 74264 3052
rect 74316 3000 74322 3052
rect 74534 3000 74540 3052
rect 74592 3000 74598 3052
rect 76650 3000 76656 3052
rect 76708 3000 76714 3052
rect 44174 2932 44180 2984
rect 44232 2972 44238 2984
rect 45649 2975 45707 2981
rect 45649 2972 45661 2975
rect 44232 2944 45661 2972
rect 44232 2932 44238 2944
rect 45649 2941 45661 2944
rect 45695 2941 45707 2975
rect 45649 2935 45707 2941
rect 45738 2932 45744 2984
rect 45796 2972 45802 2984
rect 47121 2975 47179 2981
rect 47121 2972 47133 2975
rect 45796 2944 47133 2972
rect 45796 2932 45802 2944
rect 47121 2941 47133 2944
rect 47167 2941 47179 2975
rect 47121 2935 47179 2941
rect 47670 2932 47676 2984
rect 47728 2972 47734 2984
rect 48777 2975 48835 2981
rect 48777 2972 48789 2975
rect 47728 2944 48789 2972
rect 47728 2932 47734 2944
rect 48777 2941 48789 2944
rect 48823 2941 48835 2975
rect 48777 2935 48835 2941
rect 49602 2932 49608 2984
rect 49660 2972 49666 2984
rect 50617 2975 50675 2981
rect 50617 2972 50629 2975
rect 49660 2944 50629 2972
rect 49660 2932 49666 2944
rect 50617 2941 50629 2944
rect 50663 2941 50675 2975
rect 52549 2975 52607 2981
rect 52549 2972 52561 2975
rect 50617 2935 50675 2941
rect 51552 2944 52561 2972
rect 51552 2916 51580 2944
rect 52549 2941 52561 2944
rect 52595 2941 52607 2975
rect 52549 2935 52607 2941
rect 53466 2932 53472 2984
rect 53524 2972 53530 2984
rect 54481 2975 54539 2981
rect 54481 2972 54493 2975
rect 53524 2944 54493 2972
rect 53524 2932 53530 2944
rect 54481 2941 54493 2944
rect 54527 2941 54539 2975
rect 54481 2935 54539 2941
rect 61194 2932 61200 2984
rect 61252 2972 61258 2984
rect 62209 2975 62267 2981
rect 62209 2972 62221 2975
rect 61252 2944 62221 2972
rect 61252 2932 61258 2944
rect 62209 2941 62221 2944
rect 62255 2941 62267 2975
rect 62209 2935 62267 2941
rect 65058 2932 65064 2984
rect 65116 2972 65122 2984
rect 65981 2975 66039 2981
rect 65981 2972 65993 2975
rect 65116 2944 65993 2972
rect 65116 2932 65122 2944
rect 65981 2941 65993 2944
rect 66027 2941 66039 2975
rect 68005 2975 68063 2981
rect 68005 2972 68017 2975
rect 65981 2935 66039 2941
rect 67008 2944 68017 2972
rect 67008 2916 67036 2944
rect 68005 2941 68017 2944
rect 68051 2941 68063 2975
rect 68005 2935 68063 2941
rect 68922 2932 68928 2984
rect 68980 2972 68986 2984
rect 69937 2975 69995 2981
rect 69937 2972 69949 2975
rect 68980 2944 69949 2972
rect 68980 2932 68986 2944
rect 69937 2941 69949 2944
rect 69983 2941 69995 2975
rect 69937 2935 69995 2941
rect 70854 2932 70860 2984
rect 70912 2972 70918 2984
rect 71961 2975 72019 2981
rect 71961 2972 71973 2975
rect 70912 2944 71973 2972
rect 70912 2932 70918 2944
rect 71961 2941 71973 2944
rect 72007 2941 72019 2975
rect 71961 2935 72019 2941
rect 74718 2932 74724 2984
rect 74776 2972 74782 2984
rect 75457 2975 75515 2981
rect 75457 2972 75469 2975
rect 74776 2944 75469 2972
rect 74776 2932 74782 2944
rect 75457 2941 75469 2944
rect 75503 2941 75515 2975
rect 75457 2935 75515 2941
rect 77297 2975 77355 2981
rect 77297 2941 77309 2975
rect 77343 2941 77355 2975
rect 77297 2935 77355 2941
rect 51534 2864 51540 2916
rect 51592 2864 51598 2916
rect 66990 2864 66996 2916
rect 67048 2864 67054 2916
rect 75181 2907 75239 2913
rect 75181 2873 75193 2907
rect 75227 2904 75239 2907
rect 77312 2904 77340 2935
rect 75227 2876 77340 2904
rect 75227 2873 75239 2876
rect 75181 2867 75239 2873
rect 45278 2836 45284 2848
rect 43272 2808 45284 2836
rect 40368 2796 40374 2808
rect 45278 2796 45284 2808
rect 45336 2796 45342 2848
rect 55306 2796 55312 2848
rect 55364 2836 55370 2848
rect 55493 2839 55551 2845
rect 55493 2836 55505 2839
rect 55364 2808 55505 2836
rect 55364 2796 55370 2808
rect 55493 2805 55505 2808
rect 55539 2805 55551 2839
rect 55493 2799 55551 2805
rect 59262 2796 59268 2848
rect 59320 2836 59326 2848
rect 59357 2839 59415 2845
rect 59357 2836 59369 2839
rect 59320 2808 59369 2836
rect 59320 2796 59326 2808
rect 59357 2805 59369 2808
rect 59403 2805 59415 2839
rect 59357 2799 59415 2805
rect 70486 2796 70492 2848
rect 70544 2836 70550 2848
rect 70949 2839 71007 2845
rect 70949 2836 70961 2839
rect 70544 2808 70961 2836
rect 70544 2796 70550 2808
rect 70949 2805 70961 2808
rect 70995 2805 71007 2839
rect 70949 2799 71007 2805
rect 76190 2796 76196 2848
rect 76248 2836 76254 2848
rect 76745 2839 76803 2845
rect 76745 2836 76757 2839
rect 76248 2808 76757 2836
rect 76248 2796 76254 2808
rect 76745 2805 76757 2808
rect 76791 2805 76803 2839
rect 76745 2799 76803 2805
rect 2024 2746 77924 2768
rect 2024 2694 5134 2746
rect 5186 2694 5198 2746
rect 5250 2694 5262 2746
rect 5314 2694 5326 2746
rect 5378 2694 5390 2746
rect 5442 2694 35854 2746
rect 35906 2694 35918 2746
rect 35970 2694 35982 2746
rect 36034 2694 36046 2746
rect 36098 2694 36110 2746
rect 36162 2694 66574 2746
rect 66626 2694 66638 2746
rect 66690 2694 66702 2746
rect 66754 2694 66766 2746
rect 66818 2694 66830 2746
rect 66882 2694 77924 2746
rect 2024 2672 77924 2694
rect 3789 2635 3847 2641
rect 3789 2601 3801 2635
rect 3835 2632 3847 2635
rect 3878 2632 3884 2644
rect 3835 2604 3884 2632
rect 3835 2601 3847 2604
rect 3789 2595 3847 2601
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 7650 2632 7656 2644
rect 6411 2604 7656 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 8570 2592 8576 2644
rect 8628 2592 8634 2644
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 11882 2632 11888 2644
rect 11195 2604 11888 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12066 2592 12072 2644
rect 12124 2632 12130 2644
rect 12437 2635 12495 2641
rect 12437 2632 12449 2635
rect 12124 2604 12449 2632
rect 12124 2592 12130 2604
rect 12437 2601 12449 2604
rect 12483 2601 12495 2635
rect 12437 2595 12495 2601
rect 16666 2592 16672 2644
rect 16724 2632 16730 2644
rect 16853 2635 16911 2641
rect 16853 2632 16865 2635
rect 16724 2604 16865 2632
rect 16724 2592 16730 2604
rect 16853 2601 16865 2604
rect 16899 2632 16911 2635
rect 20714 2632 20720 2644
rect 16899 2604 20720 2632
rect 16899 2601 16911 2604
rect 16853 2595 16911 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 20809 2635 20867 2641
rect 20809 2601 20821 2635
rect 20855 2632 20867 2635
rect 21910 2632 21916 2644
rect 20855 2604 21916 2632
rect 20855 2601 20867 2604
rect 20809 2595 20867 2601
rect 21910 2592 21916 2604
rect 21968 2592 21974 2644
rect 22066 2604 22876 2632
rect 3053 2567 3111 2573
rect 3053 2533 3065 2567
rect 3099 2564 3111 2567
rect 8205 2567 8263 2573
rect 3099 2536 5488 2564
rect 3099 2533 3111 2536
rect 3053 2527 3111 2533
rect 3234 2456 3240 2508
rect 3292 2456 3298 2508
rect 3970 2456 3976 2508
rect 4028 2456 4034 2508
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 4985 2499 5043 2505
rect 4985 2496 4997 2499
rect 4571 2468 4997 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 4985 2465 4997 2468
rect 5031 2465 5043 2499
rect 5460 2496 5488 2536
rect 8205 2533 8217 2567
rect 8251 2564 8263 2567
rect 8846 2564 8852 2576
rect 8251 2536 8852 2564
rect 8251 2533 8263 2536
rect 8205 2527 8263 2533
rect 8846 2524 8852 2536
rect 8904 2524 8910 2576
rect 9048 2536 15332 2564
rect 5460 2468 5856 2496
rect 4985 2459 5043 2465
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 4154 2428 4160 2440
rect 2547 2400 4160 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 4755 2400 5488 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 4890 2252 4896 2304
rect 4948 2252 4954 2304
rect 5460 2292 5488 2400
rect 5626 2388 5632 2440
rect 5684 2388 5690 2440
rect 5718 2388 5724 2440
rect 5776 2388 5782 2440
rect 5828 2428 5856 2468
rect 6546 2456 6552 2508
rect 6604 2456 6610 2508
rect 7101 2499 7159 2505
rect 7101 2465 7113 2499
rect 7147 2496 7159 2499
rect 7653 2499 7711 2505
rect 7147 2468 7604 2496
rect 7147 2465 7159 2468
rect 7101 2459 7159 2465
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 5828 2400 7481 2428
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7576 2428 7604 2468
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 8386 2496 8392 2508
rect 7699 2468 8392 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 9048 2428 9076 2536
rect 10045 2499 10103 2505
rect 10045 2465 10057 2499
rect 10091 2496 10103 2499
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 10091 2468 11805 2496
rect 10091 2465 10103 2468
rect 10045 2459 10103 2465
rect 11793 2465 11805 2468
rect 11839 2496 11851 2499
rect 13081 2499 13139 2505
rect 13081 2496 13093 2499
rect 11839 2468 13093 2496
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 13081 2465 13093 2468
rect 13127 2496 13139 2499
rect 14090 2496 14096 2508
rect 13127 2468 14096 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 14090 2456 14096 2468
rect 14148 2456 14154 2508
rect 7576 2400 9076 2428
rect 9125 2431 9183 2437
rect 7469 2391 7527 2397
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9582 2428 9588 2440
rect 9171 2400 9588 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 10594 2388 10600 2440
rect 10652 2388 10658 2440
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11664 2400 11713 2428
rect 11664 2388 11670 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12066 2388 12072 2440
rect 12124 2388 12130 2440
rect 12805 2431 12863 2437
rect 12805 2397 12817 2431
rect 12851 2428 12863 2431
rect 13722 2428 13728 2440
rect 12851 2400 13728 2428
rect 12851 2397 12863 2400
rect 12805 2391 12863 2397
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 15304 2437 15332 2536
rect 16114 2524 16120 2576
rect 16172 2564 16178 2576
rect 22066 2564 22094 2604
rect 16172 2536 22094 2564
rect 16172 2524 16178 2536
rect 22554 2524 22560 2576
rect 22612 2564 22618 2576
rect 22741 2567 22799 2573
rect 22741 2564 22753 2567
rect 22612 2536 22753 2564
rect 22612 2524 22618 2536
rect 22741 2533 22753 2536
rect 22787 2533 22799 2567
rect 22741 2527 22799 2533
rect 16485 2499 16543 2505
rect 16485 2465 16497 2499
rect 16531 2496 16543 2499
rect 17862 2496 17868 2508
rect 16531 2468 17868 2496
rect 16531 2465 16543 2468
rect 16485 2459 16543 2465
rect 17862 2456 17868 2468
rect 17920 2456 17926 2508
rect 18233 2499 18291 2505
rect 18233 2465 18245 2499
rect 18279 2465 18291 2499
rect 18233 2459 18291 2465
rect 19521 2499 19579 2505
rect 19521 2465 19533 2499
rect 19567 2496 19579 2499
rect 19886 2496 19892 2508
rect 19567 2468 19892 2496
rect 19567 2465 19579 2468
rect 19521 2459 19579 2465
rect 14645 2431 14703 2437
rect 14645 2428 14657 2431
rect 14424 2400 14657 2428
rect 14424 2388 14430 2400
rect 14645 2397 14657 2400
rect 14691 2397 14703 2431
rect 14645 2391 14703 2397
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2397 15347 2431
rect 15289 2391 15347 2397
rect 16022 2388 16028 2440
rect 16080 2428 16086 2440
rect 18049 2431 18107 2437
rect 18049 2428 18061 2431
rect 16080 2400 18061 2428
rect 16080 2388 16086 2400
rect 18049 2397 18061 2400
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 18248 2428 18276 2459
rect 19886 2456 19892 2468
rect 19944 2456 19950 2508
rect 19978 2456 19984 2508
rect 20036 2496 20042 2508
rect 20165 2499 20223 2505
rect 20165 2496 20177 2499
rect 20036 2468 20177 2496
rect 20036 2456 20042 2468
rect 20165 2465 20177 2468
rect 20211 2465 20223 2499
rect 20165 2459 20223 2465
rect 22097 2499 22155 2505
rect 22097 2465 22109 2499
rect 22143 2496 22155 2499
rect 22848 2496 22876 2604
rect 23198 2592 23204 2644
rect 23256 2632 23262 2644
rect 23293 2635 23351 2641
rect 23293 2632 23305 2635
rect 23256 2604 23305 2632
rect 23256 2592 23262 2604
rect 23293 2601 23305 2604
rect 23339 2601 23351 2635
rect 23293 2595 23351 2601
rect 25958 2592 25964 2644
rect 26016 2632 26022 2644
rect 27065 2635 27123 2641
rect 27065 2632 27077 2635
rect 26016 2604 27077 2632
rect 26016 2592 26022 2604
rect 27065 2601 27077 2604
rect 27111 2601 27123 2635
rect 27065 2595 27123 2601
rect 27154 2592 27160 2644
rect 27212 2632 27218 2644
rect 27341 2635 27399 2641
rect 27341 2632 27353 2635
rect 27212 2604 27353 2632
rect 27212 2592 27218 2604
rect 27341 2601 27353 2604
rect 27387 2601 27399 2635
rect 27341 2595 27399 2601
rect 28810 2592 28816 2644
rect 28868 2632 28874 2644
rect 30469 2635 30527 2641
rect 30469 2632 30481 2635
rect 28868 2604 30481 2632
rect 28868 2592 28874 2604
rect 30469 2601 30481 2604
rect 30515 2601 30527 2635
rect 30469 2595 30527 2601
rect 31389 2635 31447 2641
rect 31389 2601 31401 2635
rect 31435 2632 31447 2635
rect 34514 2632 34520 2644
rect 31435 2604 34520 2632
rect 31435 2601 31447 2604
rect 31389 2595 31447 2601
rect 34514 2592 34520 2604
rect 34572 2592 34578 2644
rect 35713 2635 35771 2641
rect 35713 2601 35725 2635
rect 35759 2632 35771 2635
rect 36262 2632 36268 2644
rect 35759 2604 36268 2632
rect 35759 2601 35771 2604
rect 35713 2595 35771 2601
rect 36262 2592 36268 2604
rect 36320 2592 36326 2644
rect 36354 2592 36360 2644
rect 36412 2632 36418 2644
rect 38838 2632 38844 2644
rect 36412 2604 38844 2632
rect 36412 2592 36418 2604
rect 38838 2592 38844 2604
rect 38896 2592 38902 2644
rect 41598 2592 41604 2644
rect 41656 2592 41662 2644
rect 47118 2592 47124 2644
rect 47176 2632 47182 2644
rect 47397 2635 47455 2641
rect 47397 2632 47409 2635
rect 47176 2604 47409 2632
rect 47176 2592 47182 2604
rect 47397 2601 47409 2604
rect 47443 2601 47455 2635
rect 47397 2595 47455 2601
rect 49970 2592 49976 2644
rect 50028 2592 50034 2644
rect 70857 2635 70915 2641
rect 70857 2601 70869 2635
rect 70903 2632 70915 2635
rect 72970 2632 72976 2644
rect 70903 2604 72976 2632
rect 70903 2601 70915 2604
rect 70857 2595 70915 2601
rect 72970 2592 72976 2604
rect 73028 2592 73034 2644
rect 74077 2635 74135 2641
rect 74077 2601 74089 2635
rect 74123 2632 74135 2635
rect 74626 2632 74632 2644
rect 74123 2604 74632 2632
rect 74123 2601 74135 2604
rect 74077 2595 74135 2601
rect 74626 2592 74632 2604
rect 74684 2592 74690 2644
rect 76650 2592 76656 2644
rect 76708 2632 76714 2644
rect 76837 2635 76895 2641
rect 76837 2632 76849 2635
rect 76708 2604 76849 2632
rect 76708 2592 76714 2604
rect 76837 2601 76849 2604
rect 76883 2601 76895 2635
rect 76837 2595 76895 2601
rect 23658 2524 23664 2576
rect 23716 2564 23722 2576
rect 33134 2564 33140 2576
rect 23716 2536 25452 2564
rect 23716 2524 23722 2536
rect 22143 2468 22600 2496
rect 22848 2468 23428 2496
rect 22143 2465 22155 2468
rect 22097 2459 22155 2465
rect 22572 2440 22600 2468
rect 19610 2428 19616 2440
rect 18248 2400 19616 2428
rect 5534 2320 5540 2372
rect 5592 2360 5598 2372
rect 10321 2363 10379 2369
rect 5592 2332 7328 2360
rect 5592 2320 5598 2332
rect 6454 2292 6460 2304
rect 5460 2264 6460 2292
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 7300 2301 7328 2332
rect 10321 2329 10333 2363
rect 10367 2360 10379 2363
rect 11422 2360 11428 2372
rect 10367 2332 11428 2360
rect 10367 2329 10379 2332
rect 10321 2323 10379 2329
rect 11422 2320 11428 2332
rect 11480 2320 11486 2372
rect 12618 2320 12624 2372
rect 12676 2360 12682 2372
rect 12897 2363 12955 2369
rect 12897 2360 12909 2363
rect 12676 2332 12909 2360
rect 12676 2320 12682 2332
rect 12897 2329 12909 2332
rect 12943 2329 12955 2363
rect 12897 2323 12955 2329
rect 13538 2320 13544 2372
rect 13596 2360 13602 2372
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 13596 2332 13645 2360
rect 13596 2320 13602 2332
rect 13633 2329 13645 2332
rect 13679 2329 13691 2363
rect 13633 2323 13691 2329
rect 16945 2363 17003 2369
rect 16945 2329 16957 2363
rect 16991 2360 17003 2363
rect 17126 2360 17132 2372
rect 16991 2332 17132 2360
rect 16991 2329 17003 2332
rect 16945 2323 17003 2329
rect 17126 2320 17132 2332
rect 17184 2320 17190 2372
rect 17310 2320 17316 2372
rect 17368 2320 17374 2372
rect 17957 2363 18015 2369
rect 17420 2332 17724 2360
rect 7285 2295 7343 2301
rect 7285 2261 7297 2295
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 11054 2252 11060 2304
rect 11112 2292 11118 2304
rect 11241 2295 11299 2301
rect 11241 2292 11253 2295
rect 11112 2264 11253 2292
rect 11112 2252 11118 2264
rect 11241 2261 11253 2264
rect 11287 2261 11299 2295
rect 11241 2255 11299 2261
rect 11609 2295 11667 2301
rect 11609 2261 11621 2295
rect 11655 2292 11667 2295
rect 12158 2292 12164 2304
rect 11655 2264 12164 2292
rect 11655 2261 11667 2264
rect 11609 2255 11667 2261
rect 12158 2252 12164 2264
rect 12216 2252 12222 2304
rect 12250 2252 12256 2304
rect 12308 2252 12314 2304
rect 14090 2252 14096 2304
rect 14148 2292 14154 2304
rect 17420 2292 17448 2332
rect 14148 2264 17448 2292
rect 14148 2252 14154 2264
rect 17586 2252 17592 2304
rect 17644 2252 17650 2304
rect 17696 2292 17724 2332
rect 17957 2329 17969 2363
rect 18003 2360 18015 2363
rect 18138 2360 18144 2372
rect 18003 2332 18144 2360
rect 18003 2329 18015 2332
rect 17957 2323 18015 2329
rect 18138 2320 18144 2332
rect 18196 2320 18202 2372
rect 18248 2292 18276 2400
rect 19610 2388 19616 2400
rect 19668 2388 19674 2440
rect 19794 2388 19800 2440
rect 19852 2388 19858 2440
rect 20901 2431 20959 2437
rect 20901 2397 20913 2431
rect 20947 2428 20959 2431
rect 21818 2428 21824 2440
rect 20947 2400 21824 2428
rect 20947 2397 20959 2400
rect 20901 2391 20959 2397
rect 21818 2388 21824 2400
rect 21876 2388 21882 2440
rect 22462 2388 22468 2440
rect 22520 2388 22526 2440
rect 22554 2388 22560 2440
rect 22612 2388 22618 2440
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2428 22983 2431
rect 23014 2428 23020 2440
rect 22971 2400 23020 2428
rect 22971 2397 22983 2400
rect 22925 2391 22983 2397
rect 23014 2388 23020 2400
rect 23072 2388 23078 2440
rect 23400 2437 23428 2468
rect 24762 2456 24768 2508
rect 24820 2496 24826 2508
rect 25317 2499 25375 2505
rect 25317 2496 25329 2499
rect 24820 2468 25329 2496
rect 24820 2456 24826 2468
rect 25317 2465 25329 2468
rect 25363 2465 25375 2499
rect 25424 2496 25452 2536
rect 26620 2536 30696 2564
rect 26620 2496 26648 2536
rect 25424 2468 26648 2496
rect 25317 2459 25375 2465
rect 26786 2456 26792 2508
rect 26844 2456 26850 2508
rect 29825 2499 29883 2505
rect 29825 2465 29837 2499
rect 29871 2496 29883 2499
rect 30190 2496 30196 2508
rect 29871 2468 30196 2496
rect 29871 2465 29883 2468
rect 29825 2459 29883 2465
rect 30190 2456 30196 2468
rect 30248 2456 30254 2508
rect 23385 2431 23443 2437
rect 23385 2397 23397 2431
rect 23431 2397 23443 2431
rect 26804 2428 26832 2456
rect 27525 2431 27583 2437
rect 27525 2428 27537 2431
rect 26804 2400 27537 2428
rect 23385 2391 23443 2397
rect 27525 2397 27537 2400
rect 27571 2397 27583 2431
rect 27525 2391 27583 2397
rect 28077 2431 28135 2437
rect 28077 2397 28089 2431
rect 28123 2428 28135 2431
rect 28258 2428 28264 2440
rect 28123 2400 28264 2428
rect 28123 2397 28135 2400
rect 28077 2391 28135 2397
rect 28258 2388 28264 2400
rect 28316 2388 28322 2440
rect 30285 2431 30343 2437
rect 30285 2397 30297 2431
rect 30331 2428 30343 2431
rect 30374 2428 30380 2440
rect 30331 2400 30380 2428
rect 30331 2397 30343 2400
rect 30285 2391 30343 2397
rect 30374 2388 30380 2400
rect 30432 2388 30438 2440
rect 30668 2437 30696 2536
rect 30852 2536 33140 2564
rect 30852 2505 30880 2536
rect 33134 2524 33140 2536
rect 33192 2524 33198 2576
rect 33410 2524 33416 2576
rect 33468 2564 33474 2576
rect 38197 2567 38255 2573
rect 38197 2564 38209 2567
rect 33468 2536 38209 2564
rect 33468 2524 33474 2536
rect 38197 2533 38209 2536
rect 38243 2533 38255 2567
rect 38197 2527 38255 2533
rect 39117 2567 39175 2573
rect 39117 2533 39129 2567
rect 39163 2564 39175 2567
rect 48130 2564 48136 2576
rect 39163 2536 45416 2564
rect 39163 2533 39175 2536
rect 39117 2527 39175 2533
rect 30837 2499 30895 2505
rect 30837 2465 30849 2499
rect 30883 2465 30895 2499
rect 30837 2459 30895 2465
rect 32214 2456 32220 2508
rect 32272 2456 32278 2508
rect 34698 2456 34704 2508
rect 34756 2496 34762 2508
rect 34756 2468 35388 2496
rect 34756 2456 34762 2468
rect 30653 2431 30711 2437
rect 30653 2397 30665 2431
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 31478 2388 31484 2440
rect 31536 2388 31542 2440
rect 33045 2431 33103 2437
rect 33045 2428 33057 2431
rect 31726 2400 33057 2428
rect 23109 2363 23167 2369
rect 23109 2329 23121 2363
rect 23155 2360 23167 2363
rect 25498 2360 25504 2372
rect 23155 2332 25504 2360
rect 23155 2329 23167 2332
rect 23109 2323 23167 2329
rect 25498 2320 25504 2332
rect 25556 2320 25562 2372
rect 25590 2320 25596 2372
rect 25648 2320 25654 2372
rect 26234 2320 26240 2372
rect 26292 2320 26298 2372
rect 27709 2363 27767 2369
rect 27709 2329 27721 2363
rect 27755 2360 27767 2363
rect 28350 2360 28356 2372
rect 27755 2332 28356 2360
rect 27755 2329 27767 2332
rect 27709 2323 27767 2329
rect 28350 2320 28356 2332
rect 28408 2320 28414 2372
rect 28813 2363 28871 2369
rect 28813 2329 28825 2363
rect 28859 2360 28871 2363
rect 31726 2360 31754 2400
rect 33045 2397 33057 2400
rect 33091 2397 33103 2431
rect 33045 2391 33103 2397
rect 33410 2388 33416 2440
rect 33468 2388 33474 2440
rect 35250 2388 35256 2440
rect 35308 2388 35314 2440
rect 35360 2428 35388 2468
rect 35526 2456 35532 2508
rect 35584 2496 35590 2508
rect 35584 2468 35848 2496
rect 35584 2456 35590 2468
rect 35820 2437 35848 2468
rect 36078 2456 36084 2508
rect 36136 2496 36142 2508
rect 37093 2499 37151 2505
rect 37093 2496 37105 2499
rect 36136 2468 37105 2496
rect 36136 2456 36142 2468
rect 37093 2465 37105 2468
rect 37139 2465 37151 2499
rect 37093 2459 37151 2465
rect 38565 2499 38623 2505
rect 38565 2465 38577 2499
rect 38611 2496 38623 2499
rect 39482 2496 39488 2508
rect 38611 2468 39488 2496
rect 38611 2465 38623 2468
rect 38565 2459 38623 2465
rect 39482 2456 39488 2468
rect 39540 2456 39546 2508
rect 39942 2456 39948 2508
rect 40000 2456 40006 2508
rect 40310 2456 40316 2508
rect 40368 2496 40374 2508
rect 45388 2505 45416 2536
rect 45756 2536 48136 2564
rect 40957 2499 41015 2505
rect 40957 2496 40969 2499
rect 40368 2468 40969 2496
rect 40368 2456 40374 2468
rect 40957 2465 40969 2468
rect 41003 2465 41015 2499
rect 44821 2499 44879 2505
rect 44821 2496 44833 2499
rect 40957 2459 41015 2465
rect 41386 2468 44833 2496
rect 35621 2431 35679 2437
rect 35621 2428 35633 2431
rect 35360 2400 35633 2428
rect 35621 2397 35633 2400
rect 35667 2397 35679 2431
rect 35621 2391 35679 2397
rect 35805 2431 35863 2437
rect 35805 2397 35817 2431
rect 35851 2397 35863 2431
rect 35805 2391 35863 2397
rect 35989 2431 36047 2437
rect 35989 2397 36001 2431
rect 36035 2397 36047 2431
rect 35989 2391 36047 2397
rect 36817 2431 36875 2437
rect 36817 2397 36829 2431
rect 36863 2428 36875 2431
rect 36906 2428 36912 2440
rect 36863 2400 36912 2428
rect 36863 2397 36875 2400
rect 36817 2391 36875 2397
rect 28859 2332 31754 2360
rect 28859 2329 28871 2332
rect 28813 2323 28871 2329
rect 34146 2320 34152 2372
rect 34204 2360 34210 2372
rect 34241 2363 34299 2369
rect 34241 2360 34253 2363
rect 34204 2332 34253 2360
rect 34204 2320 34210 2332
rect 34241 2329 34253 2332
rect 34287 2329 34299 2363
rect 36004 2360 36032 2391
rect 36906 2388 36912 2400
rect 36964 2388 36970 2440
rect 38378 2388 38384 2440
rect 38436 2388 38442 2440
rect 39390 2388 39396 2440
rect 39448 2388 39454 2440
rect 41138 2388 41144 2440
rect 41196 2428 41202 2440
rect 41233 2431 41291 2437
rect 41233 2428 41245 2431
rect 41196 2400 41245 2428
rect 41196 2388 41202 2400
rect 41233 2397 41245 2400
rect 41279 2397 41291 2431
rect 41233 2391 41291 2397
rect 41046 2360 41052 2372
rect 36004 2332 41052 2360
rect 34241 2323 34299 2329
rect 41046 2320 41052 2332
rect 41104 2320 41110 2372
rect 41386 2360 41414 2468
rect 44821 2465 44833 2468
rect 44867 2465 44879 2499
rect 44821 2459 44879 2465
rect 45373 2499 45431 2505
rect 45373 2465 45385 2499
rect 45419 2465 45431 2499
rect 45373 2459 45431 2465
rect 41966 2388 41972 2440
rect 42024 2388 42030 2440
rect 45756 2437 45784 2536
rect 48130 2524 48136 2536
rect 48188 2524 48194 2576
rect 49602 2524 49608 2576
rect 49660 2564 49666 2576
rect 50709 2567 50767 2573
rect 50709 2564 50721 2567
rect 49660 2536 50721 2564
rect 49660 2524 49666 2536
rect 50709 2533 50721 2536
rect 50755 2533 50767 2567
rect 50709 2527 50767 2533
rect 46750 2456 46756 2508
rect 46808 2456 46814 2508
rect 49421 2499 49479 2505
rect 49421 2465 49433 2499
rect 49467 2496 49479 2499
rect 49786 2496 49792 2508
rect 49467 2468 49792 2496
rect 49467 2465 49479 2468
rect 49421 2459 49479 2465
rect 49786 2456 49792 2468
rect 49844 2456 49850 2508
rect 50522 2456 50528 2508
rect 50580 2456 50586 2508
rect 52086 2456 52092 2508
rect 52144 2456 52150 2508
rect 54018 2456 54024 2508
rect 54076 2456 54082 2508
rect 58161 2499 58219 2505
rect 58161 2465 58173 2499
rect 58207 2496 58219 2499
rect 59265 2499 59323 2505
rect 58207 2468 58848 2496
rect 58207 2465 58219 2468
rect 58161 2459 58219 2465
rect 42981 2431 43039 2437
rect 42981 2397 42993 2431
rect 43027 2428 43039 2431
rect 43349 2431 43407 2437
rect 43349 2428 43361 2431
rect 43027 2400 43361 2428
rect 43027 2397 43039 2400
rect 42981 2391 43039 2397
rect 43349 2397 43361 2400
rect 43395 2397 43407 2431
rect 43349 2391 43407 2397
rect 45741 2431 45799 2437
rect 45741 2397 45753 2431
rect 45787 2397 45799 2431
rect 45741 2391 45799 2397
rect 45830 2388 45836 2440
rect 45888 2428 45894 2440
rect 45925 2431 45983 2437
rect 45925 2428 45937 2431
rect 45888 2400 45937 2428
rect 45888 2388 45894 2400
rect 45925 2397 45937 2400
rect 45971 2397 45983 2431
rect 45925 2391 45983 2397
rect 47946 2388 47952 2440
rect 48004 2388 48010 2440
rect 48317 2431 48375 2437
rect 48317 2397 48329 2431
rect 48363 2428 48375 2431
rect 48406 2428 48412 2440
rect 48363 2400 48412 2428
rect 48363 2397 48375 2400
rect 48317 2391 48375 2397
rect 48406 2388 48412 2400
rect 48464 2388 48470 2440
rect 49694 2388 49700 2440
rect 49752 2388 49758 2440
rect 52822 2388 52828 2440
rect 52880 2388 52886 2440
rect 55033 2431 55091 2437
rect 55033 2397 55045 2431
rect 55079 2428 55091 2431
rect 55306 2428 55312 2440
rect 55079 2400 55312 2428
rect 55079 2397 55091 2400
rect 55033 2391 55091 2397
rect 55306 2388 55312 2400
rect 55364 2388 55370 2440
rect 55398 2388 55404 2440
rect 55456 2428 55462 2440
rect 55493 2431 55551 2437
rect 55493 2428 55505 2431
rect 55456 2400 55505 2428
rect 55456 2388 55462 2400
rect 55493 2397 55505 2400
rect 55539 2397 55551 2431
rect 55493 2391 55551 2397
rect 58618 2388 58624 2440
rect 58676 2388 58682 2440
rect 58820 2437 58848 2468
rect 59265 2465 59277 2499
rect 59311 2465 59323 2499
rect 59265 2459 59323 2465
rect 58805 2431 58863 2437
rect 58805 2397 58817 2431
rect 58851 2397 58863 2431
rect 58805 2391 58863 2397
rect 41156 2332 41414 2360
rect 17696 2264 18276 2292
rect 21082 2252 21088 2304
rect 21140 2252 21146 2304
rect 22922 2252 22928 2304
rect 22980 2292 22986 2304
rect 23017 2295 23075 2301
rect 23017 2292 23029 2295
rect 22980 2264 23029 2292
rect 22980 2252 22986 2264
rect 23017 2261 23029 2264
rect 23063 2261 23075 2295
rect 23017 2255 23075 2261
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 24673 2295 24731 2301
rect 24673 2292 24685 2295
rect 24544 2264 24685 2292
rect 24544 2252 24550 2264
rect 24673 2261 24685 2264
rect 24719 2261 24731 2295
rect 24673 2255 24731 2261
rect 33226 2252 33232 2304
rect 33284 2252 33290 2304
rect 33965 2295 34023 2301
rect 33965 2261 33977 2295
rect 34011 2292 34023 2295
rect 36354 2292 36360 2304
rect 34011 2264 36360 2292
rect 34011 2261 34023 2264
rect 33965 2255 34023 2261
rect 36354 2252 36360 2264
rect 36412 2252 36418 2304
rect 36541 2295 36599 2301
rect 36541 2261 36553 2295
rect 36587 2292 36599 2295
rect 38102 2292 38108 2304
rect 36587 2264 38108 2292
rect 36587 2261 36599 2264
rect 36541 2255 36599 2261
rect 38102 2252 38108 2264
rect 38160 2252 38166 2304
rect 41156 2301 41184 2332
rect 41874 2320 41880 2372
rect 41932 2360 41938 2372
rect 44269 2363 44327 2369
rect 44269 2360 44281 2363
rect 41932 2332 44281 2360
rect 41932 2320 41938 2332
rect 44269 2329 44281 2332
rect 44315 2329 44327 2363
rect 44269 2323 44327 2329
rect 57330 2320 57336 2372
rect 57388 2360 57394 2372
rect 59280 2360 59308 2459
rect 61746 2456 61752 2508
rect 61804 2456 61810 2508
rect 65518 2456 65524 2508
rect 65576 2456 65582 2508
rect 67634 2456 67640 2508
rect 67692 2456 67698 2508
rect 69474 2456 69480 2508
rect 69532 2456 69538 2508
rect 70302 2456 70308 2508
rect 70360 2496 70366 2508
rect 70360 2468 70716 2496
rect 70360 2456 70366 2468
rect 62758 2388 62764 2440
rect 62816 2388 62822 2440
rect 63126 2388 63132 2440
rect 63184 2428 63190 2440
rect 63221 2431 63279 2437
rect 63221 2428 63233 2431
rect 63184 2400 63233 2428
rect 63184 2388 63190 2400
rect 63221 2397 63233 2400
rect 63267 2397 63279 2431
rect 63221 2391 63279 2397
rect 66254 2388 66260 2440
rect 66312 2388 66318 2440
rect 68278 2388 68284 2440
rect 68336 2388 68342 2440
rect 70486 2388 70492 2440
rect 70544 2388 70550 2440
rect 70688 2437 70716 2468
rect 72602 2456 72608 2508
rect 72660 2456 72666 2508
rect 72786 2456 72792 2508
rect 72844 2496 72850 2508
rect 73157 2499 73215 2505
rect 73157 2496 73169 2499
rect 72844 2468 73169 2496
rect 72844 2456 72850 2468
rect 73157 2465 73169 2468
rect 73203 2465 73215 2499
rect 73157 2459 73215 2465
rect 73525 2499 73583 2505
rect 73525 2465 73537 2499
rect 73571 2496 73583 2499
rect 75454 2496 75460 2508
rect 73571 2468 75460 2496
rect 73571 2465 73583 2468
rect 73525 2459 73583 2465
rect 75454 2456 75460 2468
rect 75512 2456 75518 2508
rect 75733 2499 75791 2505
rect 75733 2465 75745 2499
rect 75779 2496 75791 2499
rect 77389 2499 77447 2505
rect 77389 2496 77401 2499
rect 75779 2468 77401 2496
rect 75779 2465 75791 2468
rect 75733 2459 75791 2465
rect 77389 2465 77401 2468
rect 77435 2465 77447 2499
rect 77389 2459 77447 2465
rect 70673 2431 70731 2437
rect 70673 2397 70685 2431
rect 70719 2397 70731 2431
rect 70673 2391 70731 2397
rect 73065 2431 73123 2437
rect 73065 2397 73077 2431
rect 73111 2428 73123 2431
rect 73246 2428 73252 2440
rect 73111 2400 73252 2428
rect 73111 2397 73123 2400
rect 73065 2391 73123 2397
rect 73246 2388 73252 2400
rect 73304 2388 73310 2440
rect 76190 2388 76196 2440
rect 76248 2388 76254 2440
rect 57388 2332 59308 2360
rect 57388 2320 57394 2332
rect 41141 2295 41199 2301
rect 41141 2261 41153 2295
rect 41187 2261 41199 2295
rect 41141 2255 41199 2261
rect 41322 2252 41328 2304
rect 41380 2292 41386 2304
rect 45557 2295 45615 2301
rect 45557 2292 45569 2295
rect 41380 2264 45569 2292
rect 41380 2252 41386 2264
rect 45557 2261 45569 2264
rect 45603 2261 45615 2295
rect 45557 2255 45615 2261
rect 47578 2252 47584 2304
rect 47636 2292 47642 2304
rect 48133 2295 48191 2301
rect 48133 2292 48145 2295
rect 47636 2264 48145 2292
rect 47636 2252 47642 2264
rect 48133 2261 48145 2264
rect 48179 2261 48191 2295
rect 48133 2255 48191 2261
rect 2024 2202 77924 2224
rect 2024 2150 5794 2202
rect 5846 2150 5858 2202
rect 5910 2150 5922 2202
rect 5974 2150 5986 2202
rect 6038 2150 6050 2202
rect 6102 2150 36514 2202
rect 36566 2150 36578 2202
rect 36630 2150 36642 2202
rect 36694 2150 36706 2202
rect 36758 2150 36770 2202
rect 36822 2150 67234 2202
rect 67286 2150 67298 2202
rect 67350 2150 67362 2202
rect 67414 2150 67426 2202
rect 67478 2150 67490 2202
rect 67542 2150 77924 2202
rect 2024 2128 77924 2150
rect 12250 2048 12256 2100
rect 12308 2088 12314 2100
rect 17218 2088 17224 2100
rect 12308 2060 17224 2088
rect 12308 2048 12314 2060
rect 17218 2048 17224 2060
rect 17276 2048 17282 2100
rect 20530 2048 20536 2100
rect 20588 2088 20594 2100
rect 30926 2088 30932 2100
rect 20588 2060 30932 2088
rect 20588 2048 20594 2060
rect 30926 2048 30932 2060
rect 30984 2048 30990 2100
rect 38102 2048 38108 2100
rect 38160 2088 38166 2100
rect 47946 2088 47952 2100
rect 38160 2060 47952 2088
rect 38160 2048 38166 2060
rect 47946 2048 47952 2060
rect 48004 2048 48010 2100
rect 10226 1980 10232 2032
rect 10284 2020 10290 2032
rect 12618 2020 12624 2032
rect 10284 1992 12624 2020
rect 10284 1980 10290 1992
rect 12618 1980 12624 1992
rect 12676 1980 12682 2032
rect 18966 1980 18972 2032
rect 19024 2020 19030 2032
rect 32398 2020 32404 2032
rect 19024 1992 32404 2020
rect 19024 1980 19030 1992
rect 32398 1980 32404 1992
rect 32456 1980 32462 2032
rect 33410 1980 33416 2032
rect 33468 2020 33474 2032
rect 40586 2020 40592 2032
rect 33468 1992 40592 2020
rect 33468 1980 33474 1992
rect 40586 1980 40592 1992
rect 40644 1980 40650 2032
rect 9858 1912 9864 1964
rect 9916 1952 9922 1964
rect 17586 1952 17592 1964
rect 9916 1924 17592 1952
rect 9916 1912 9922 1924
rect 17586 1912 17592 1924
rect 17644 1912 17650 1964
rect 27522 1912 27528 1964
rect 27580 1952 27586 1964
rect 38378 1952 38384 1964
rect 27580 1924 38384 1952
rect 27580 1912 27586 1924
rect 38378 1912 38384 1924
rect 38436 1912 38442 1964
rect 12066 1844 12072 1896
rect 12124 1884 12130 1896
rect 17402 1884 17408 1896
rect 12124 1856 17408 1884
rect 12124 1844 12130 1856
rect 17402 1844 17408 1856
rect 17460 1844 17466 1896
rect 21818 1844 21824 1896
rect 21876 1884 21882 1896
rect 21876 1856 33180 1884
rect 21876 1844 21882 1856
rect 5718 1776 5724 1828
rect 5776 1816 5782 1828
rect 13906 1816 13912 1828
rect 5776 1788 13912 1816
rect 5776 1776 5782 1788
rect 13906 1776 13912 1788
rect 13964 1776 13970 1828
rect 18506 1776 18512 1828
rect 18564 1816 18570 1828
rect 31938 1816 31944 1828
rect 18564 1788 31944 1816
rect 18564 1776 18570 1788
rect 31938 1776 31944 1788
rect 31996 1776 32002 1828
rect 33152 1816 33180 1856
rect 33226 1844 33232 1896
rect 33284 1884 33290 1896
rect 38286 1884 38292 1896
rect 33284 1856 38292 1884
rect 33284 1844 33290 1856
rect 38286 1844 38292 1856
rect 38344 1844 38350 1896
rect 38194 1816 38200 1828
rect 33152 1788 38200 1816
rect 38194 1776 38200 1788
rect 38252 1776 38258 1828
rect 23934 1708 23940 1760
rect 23992 1748 23998 1760
rect 40770 1748 40776 1760
rect 23992 1720 40776 1748
rect 23992 1708 23998 1720
rect 40770 1708 40776 1720
rect 40828 1708 40834 1760
rect 15654 1640 15660 1692
rect 15712 1680 15718 1692
rect 25590 1680 25596 1692
rect 15712 1652 25596 1680
rect 15712 1640 15718 1652
rect 25590 1640 25596 1652
rect 25648 1640 25654 1692
rect 18874 1572 18880 1624
rect 18932 1612 18938 1624
rect 31478 1612 31484 1624
rect 18932 1584 31484 1612
rect 18932 1572 18938 1584
rect 31478 1572 31484 1584
rect 31536 1572 31542 1624
rect 8018 1368 8024 1420
rect 8076 1408 8082 1420
rect 9674 1408 9680 1420
rect 8076 1380 9680 1408
rect 8076 1368 8082 1380
rect 9674 1368 9680 1380
rect 9732 1368 9738 1420
rect 14274 1368 14280 1420
rect 14332 1408 14338 1420
rect 21266 1408 21272 1420
rect 14332 1380 21272 1408
rect 14332 1368 14338 1380
rect 21266 1368 21272 1380
rect 21324 1368 21330 1420
rect 22186 1368 22192 1420
rect 22244 1408 22250 1420
rect 23198 1408 23204 1420
rect 22244 1380 23204 1408
rect 22244 1368 22250 1380
rect 23198 1368 23204 1380
rect 23256 1368 23262 1420
rect 10042 1300 10048 1352
rect 10100 1340 10106 1352
rect 16114 1340 16120 1352
rect 10100 1312 16120 1340
rect 10100 1300 10106 1312
rect 16114 1300 16120 1312
rect 16172 1300 16178 1352
rect 17034 1300 17040 1352
rect 17092 1340 17098 1352
rect 19334 1340 19340 1352
rect 17092 1312 19340 1340
rect 17092 1300 17098 1312
rect 19334 1300 19340 1312
rect 19392 1300 19398 1352
rect 13262 1232 13268 1284
rect 13320 1272 13326 1284
rect 18046 1272 18052 1284
rect 13320 1244 18052 1272
rect 13320 1232 13326 1244
rect 18046 1232 18052 1244
rect 18104 1232 18110 1284
rect 16942 1164 16948 1216
rect 17000 1204 17006 1216
rect 25774 1204 25780 1216
rect 17000 1176 25780 1204
rect 17000 1164 17006 1176
rect 25774 1164 25780 1176
rect 25832 1164 25838 1216
rect 21174 280 21180 332
rect 21232 320 21238 332
rect 29546 320 29552 332
rect 21232 292 29552 320
rect 21232 280 21238 292
rect 29546 280 29552 292
rect 29604 280 29610 332
rect 10686 212 10692 264
rect 10744 252 10750 264
rect 21818 252 21824 264
rect 10744 224 21824 252
rect 10744 212 10750 224
rect 21818 212 21824 224
rect 21876 212 21882 264
rect 21542 144 21548 196
rect 21600 184 21606 196
rect 33410 184 33416 196
rect 21600 156 33416 184
rect 21600 144 21606 156
rect 33410 144 33416 156
rect 33468 144 33474 196
rect 9582 76 9588 128
rect 9640 116 9646 128
rect 23750 116 23756 128
rect 9640 88 23756 116
rect 9640 76 9646 88
rect 23750 76 23756 88
rect 23808 76 23814 128
<< via1 >>
rect 5134 37510 5186 37562
rect 5198 37510 5250 37562
rect 5262 37510 5314 37562
rect 5326 37510 5378 37562
rect 5390 37510 5442 37562
rect 35854 37510 35906 37562
rect 35918 37510 35970 37562
rect 35982 37510 36034 37562
rect 36046 37510 36098 37562
rect 36110 37510 36162 37562
rect 66574 37510 66626 37562
rect 66638 37510 66690 37562
rect 66702 37510 66754 37562
rect 66766 37510 66818 37562
rect 66830 37510 66882 37562
rect 2228 37272 2280 37324
rect 13268 37272 13320 37324
rect 33508 37272 33560 37324
rect 39028 37272 39080 37324
rect 3516 37247 3568 37256
rect 3516 37213 3525 37247
rect 3525 37213 3559 37247
rect 3559 37213 3568 37247
rect 3516 37204 3568 37213
rect 5908 37247 5960 37256
rect 5908 37213 5917 37247
rect 5917 37213 5951 37247
rect 5951 37213 5960 37247
rect 5908 37204 5960 37213
rect 7104 37247 7156 37256
rect 7104 37213 7113 37247
rect 7113 37213 7147 37247
rect 7147 37213 7156 37247
rect 7104 37204 7156 37213
rect 7748 37204 7800 37256
rect 7932 37204 7984 37256
rect 11428 37204 11480 37256
rect 11888 37204 11940 37256
rect 14556 37247 14608 37256
rect 14556 37213 14565 37247
rect 14565 37213 14599 37247
rect 14599 37213 14608 37247
rect 14556 37204 14608 37213
rect 15108 37204 15160 37256
rect 18696 37247 18748 37256
rect 18696 37213 18705 37247
rect 18705 37213 18739 37247
rect 18739 37213 18748 37247
rect 18696 37204 18748 37213
rect 18788 37204 18840 37256
rect 20628 37204 20680 37256
rect 21916 37247 21968 37256
rect 21916 37213 21925 37247
rect 21925 37213 21959 37247
rect 21959 37213 21968 37247
rect 21916 37204 21968 37213
rect 22468 37204 22520 37256
rect 26056 37204 26108 37256
rect 27988 37204 28040 37256
rect 15016 37136 15068 37188
rect 22560 37136 22612 37188
rect 26148 37136 26200 37188
rect 31668 37204 31720 37256
rect 32680 37247 32732 37256
rect 32680 37213 32689 37247
rect 32689 37213 32723 37247
rect 32723 37213 32732 37247
rect 32680 37204 32732 37213
rect 33784 37247 33836 37256
rect 33784 37213 33793 37247
rect 33793 37213 33827 37247
rect 33827 37213 33836 37247
rect 33784 37204 33836 37213
rect 37004 37204 37056 37256
rect 37188 37204 37240 37256
rect 39120 37247 39172 37256
rect 39120 37213 39129 37247
rect 39129 37213 39163 37247
rect 39163 37213 39172 37247
rect 39120 37204 39172 37213
rect 40868 37204 40920 37256
rect 41052 37204 41104 37256
rect 43352 37247 43404 37256
rect 43352 37213 43361 37247
rect 43361 37213 43395 37247
rect 43395 37213 43404 37247
rect 43352 37204 43404 37213
rect 46480 37247 46532 37256
rect 46480 37213 46489 37247
rect 46489 37213 46523 37247
rect 46523 37213 46532 37247
rect 46480 37204 46532 37213
rect 48228 37204 48280 37256
rect 51908 37204 51960 37256
rect 52092 37204 52144 37256
rect 53840 37247 53892 37256
rect 53840 37213 53849 37247
rect 53849 37213 53883 37247
rect 53883 37213 53892 37247
rect 53840 37204 53892 37213
rect 55588 37204 55640 37256
rect 58808 37247 58860 37256
rect 58808 37213 58817 37247
rect 58817 37213 58851 37247
rect 58851 37213 58860 37247
rect 58808 37204 58860 37213
rect 33048 37136 33100 37188
rect 42708 37136 42760 37188
rect 46388 37136 46440 37188
rect 48136 37136 48188 37188
rect 53748 37136 53800 37188
rect 55680 37136 55732 37188
rect 57428 37136 57480 37188
rect 5794 36966 5846 37018
rect 5858 36966 5910 37018
rect 5922 36966 5974 37018
rect 5986 36966 6038 37018
rect 6050 36966 6102 37018
rect 36514 36966 36566 37018
rect 36578 36966 36630 37018
rect 36642 36966 36694 37018
rect 36706 36966 36758 37018
rect 36770 36966 36822 37018
rect 67234 36966 67286 37018
rect 67298 36966 67350 37018
rect 67362 36966 67414 37018
rect 67426 36966 67478 37018
rect 67490 36966 67542 37018
rect 7748 36907 7800 36916
rect 7748 36873 7757 36907
rect 7757 36873 7791 36907
rect 7791 36873 7800 36907
rect 7748 36864 7800 36873
rect 11888 36907 11940 36916
rect 11888 36873 11897 36907
rect 11897 36873 11931 36907
rect 11931 36873 11940 36907
rect 11888 36864 11940 36873
rect 15108 36907 15160 36916
rect 15108 36873 15117 36907
rect 15117 36873 15151 36907
rect 15151 36873 15160 36907
rect 15108 36864 15160 36873
rect 18696 36864 18748 36916
rect 22468 36907 22520 36916
rect 22468 36873 22477 36907
rect 22477 36873 22511 36907
rect 22511 36873 22520 36907
rect 22468 36864 22520 36873
rect 26056 36864 26108 36916
rect 4068 36796 4120 36848
rect 9588 36796 9640 36848
rect 16948 36796 17000 36848
rect 24308 36796 24360 36848
rect 10968 36771 11020 36780
rect 10968 36737 10977 36771
rect 10977 36737 11011 36771
rect 11011 36737 11020 36771
rect 10968 36728 11020 36737
rect 11796 36771 11848 36780
rect 11796 36737 11805 36771
rect 11805 36737 11839 36771
rect 11839 36737 11848 36771
rect 11796 36728 11848 36737
rect 18788 36771 18840 36780
rect 18788 36737 18797 36771
rect 18797 36737 18831 36771
rect 18831 36737 18840 36771
rect 18788 36728 18840 36737
rect 25780 36771 25832 36780
rect 25780 36737 25789 36771
rect 25789 36737 25823 36771
rect 25823 36737 25832 36771
rect 25780 36728 25832 36737
rect 29828 36796 29880 36848
rect 33784 36907 33836 36916
rect 33784 36873 33793 36907
rect 33793 36873 33827 36907
rect 33827 36873 33836 36907
rect 33784 36864 33836 36873
rect 37004 36907 37056 36916
rect 37004 36873 37013 36907
rect 37013 36873 37047 36907
rect 37047 36873 37056 36907
rect 37004 36864 37056 36873
rect 40868 36907 40920 36916
rect 40868 36873 40877 36907
rect 40877 36873 40911 36907
rect 40911 36873 40920 36907
rect 40868 36864 40920 36873
rect 48228 36907 48280 36916
rect 48228 36873 48237 36907
rect 48237 36873 48271 36907
rect 48271 36873 48280 36907
rect 48228 36864 48280 36873
rect 51908 36907 51960 36916
rect 51908 36873 51917 36907
rect 51917 36873 51951 36907
rect 51951 36873 51960 36907
rect 51908 36864 51960 36873
rect 55588 36907 55640 36916
rect 55588 36873 55597 36907
rect 55597 36873 55631 36907
rect 55631 36873 55640 36907
rect 55588 36864 55640 36873
rect 11796 36592 11848 36644
rect 35440 36771 35492 36780
rect 35440 36737 35449 36771
rect 35449 36737 35483 36771
rect 35483 36737 35492 36771
rect 35440 36728 35492 36737
rect 35348 36660 35400 36712
rect 44732 36660 44784 36712
rect 50160 36771 50212 36780
rect 50160 36737 50169 36771
rect 50169 36737 50203 36771
rect 50203 36737 50212 36771
rect 50160 36728 50212 36737
rect 59268 36796 59320 36848
rect 50068 36660 50120 36712
rect 5134 36422 5186 36474
rect 5198 36422 5250 36474
rect 5262 36422 5314 36474
rect 5326 36422 5378 36474
rect 5390 36422 5442 36474
rect 35854 36422 35906 36474
rect 35918 36422 35970 36474
rect 35982 36422 36034 36474
rect 36046 36422 36098 36474
rect 36110 36422 36162 36474
rect 66574 36422 66626 36474
rect 66638 36422 66690 36474
rect 66702 36422 66754 36474
rect 66766 36422 66818 36474
rect 66830 36422 66882 36474
rect 25780 36320 25832 36372
rect 33232 36320 33284 36372
rect 5794 35878 5846 35930
rect 5858 35878 5910 35930
rect 5922 35878 5974 35930
rect 5986 35878 6038 35930
rect 6050 35878 6102 35930
rect 36514 35878 36566 35930
rect 36578 35878 36630 35930
rect 36642 35878 36694 35930
rect 36706 35878 36758 35930
rect 36770 35878 36822 35930
rect 67234 35878 67286 35930
rect 67298 35878 67350 35930
rect 67362 35878 67414 35930
rect 67426 35878 67478 35930
rect 67490 35878 67542 35930
rect 5134 35334 5186 35386
rect 5198 35334 5250 35386
rect 5262 35334 5314 35386
rect 5326 35334 5378 35386
rect 5390 35334 5442 35386
rect 35854 35334 35906 35386
rect 35918 35334 35970 35386
rect 35982 35334 36034 35386
rect 36046 35334 36098 35386
rect 36110 35334 36162 35386
rect 66574 35334 66626 35386
rect 66638 35334 66690 35386
rect 66702 35334 66754 35386
rect 66766 35334 66818 35386
rect 66830 35334 66882 35386
rect 5794 34790 5846 34842
rect 5858 34790 5910 34842
rect 5922 34790 5974 34842
rect 5986 34790 6038 34842
rect 6050 34790 6102 34842
rect 36514 34790 36566 34842
rect 36578 34790 36630 34842
rect 36642 34790 36694 34842
rect 36706 34790 36758 34842
rect 36770 34790 36822 34842
rect 67234 34790 67286 34842
rect 67298 34790 67350 34842
rect 67362 34790 67414 34842
rect 67426 34790 67478 34842
rect 67490 34790 67542 34842
rect 5134 34246 5186 34298
rect 5198 34246 5250 34298
rect 5262 34246 5314 34298
rect 5326 34246 5378 34298
rect 5390 34246 5442 34298
rect 35854 34246 35906 34298
rect 35918 34246 35970 34298
rect 35982 34246 36034 34298
rect 36046 34246 36098 34298
rect 36110 34246 36162 34298
rect 66574 34246 66626 34298
rect 66638 34246 66690 34298
rect 66702 34246 66754 34298
rect 66766 34246 66818 34298
rect 66830 34246 66882 34298
rect 5794 33702 5846 33754
rect 5858 33702 5910 33754
rect 5922 33702 5974 33754
rect 5986 33702 6038 33754
rect 6050 33702 6102 33754
rect 36514 33702 36566 33754
rect 36578 33702 36630 33754
rect 36642 33702 36694 33754
rect 36706 33702 36758 33754
rect 36770 33702 36822 33754
rect 67234 33702 67286 33754
rect 67298 33702 67350 33754
rect 67362 33702 67414 33754
rect 67426 33702 67478 33754
rect 67490 33702 67542 33754
rect 5134 33158 5186 33210
rect 5198 33158 5250 33210
rect 5262 33158 5314 33210
rect 5326 33158 5378 33210
rect 5390 33158 5442 33210
rect 35854 33158 35906 33210
rect 35918 33158 35970 33210
rect 35982 33158 36034 33210
rect 36046 33158 36098 33210
rect 36110 33158 36162 33210
rect 66574 33158 66626 33210
rect 66638 33158 66690 33210
rect 66702 33158 66754 33210
rect 66766 33158 66818 33210
rect 66830 33158 66882 33210
rect 5794 32614 5846 32666
rect 5858 32614 5910 32666
rect 5922 32614 5974 32666
rect 5986 32614 6038 32666
rect 6050 32614 6102 32666
rect 36514 32614 36566 32666
rect 36578 32614 36630 32666
rect 36642 32614 36694 32666
rect 36706 32614 36758 32666
rect 36770 32614 36822 32666
rect 67234 32614 67286 32666
rect 67298 32614 67350 32666
rect 67362 32614 67414 32666
rect 67426 32614 67478 32666
rect 67490 32614 67542 32666
rect 27252 32376 27304 32428
rect 50160 32376 50212 32428
rect 5134 32070 5186 32122
rect 5198 32070 5250 32122
rect 5262 32070 5314 32122
rect 5326 32070 5378 32122
rect 5390 32070 5442 32122
rect 35854 32070 35906 32122
rect 35918 32070 35970 32122
rect 35982 32070 36034 32122
rect 36046 32070 36098 32122
rect 36110 32070 36162 32122
rect 66574 32070 66626 32122
rect 66638 32070 66690 32122
rect 66702 32070 66754 32122
rect 66766 32070 66818 32122
rect 66830 32070 66882 32122
rect 5794 31526 5846 31578
rect 5858 31526 5910 31578
rect 5922 31526 5974 31578
rect 5986 31526 6038 31578
rect 6050 31526 6102 31578
rect 36514 31526 36566 31578
rect 36578 31526 36630 31578
rect 36642 31526 36694 31578
rect 36706 31526 36758 31578
rect 36770 31526 36822 31578
rect 67234 31526 67286 31578
rect 67298 31526 67350 31578
rect 67362 31526 67414 31578
rect 67426 31526 67478 31578
rect 67490 31526 67542 31578
rect 5134 30982 5186 31034
rect 5198 30982 5250 31034
rect 5262 30982 5314 31034
rect 5326 30982 5378 31034
rect 5390 30982 5442 31034
rect 35854 30982 35906 31034
rect 35918 30982 35970 31034
rect 35982 30982 36034 31034
rect 36046 30982 36098 31034
rect 36110 30982 36162 31034
rect 66574 30982 66626 31034
rect 66638 30982 66690 31034
rect 66702 30982 66754 31034
rect 66766 30982 66818 31034
rect 66830 30982 66882 31034
rect 5794 30438 5846 30490
rect 5858 30438 5910 30490
rect 5922 30438 5974 30490
rect 5986 30438 6038 30490
rect 6050 30438 6102 30490
rect 36514 30438 36566 30490
rect 36578 30438 36630 30490
rect 36642 30438 36694 30490
rect 36706 30438 36758 30490
rect 36770 30438 36822 30490
rect 67234 30438 67286 30490
rect 67298 30438 67350 30490
rect 67362 30438 67414 30490
rect 67426 30438 67478 30490
rect 67490 30438 67542 30490
rect 5134 29894 5186 29946
rect 5198 29894 5250 29946
rect 5262 29894 5314 29946
rect 5326 29894 5378 29946
rect 5390 29894 5442 29946
rect 35854 29894 35906 29946
rect 35918 29894 35970 29946
rect 35982 29894 36034 29946
rect 36046 29894 36098 29946
rect 36110 29894 36162 29946
rect 66574 29894 66626 29946
rect 66638 29894 66690 29946
rect 66702 29894 66754 29946
rect 66766 29894 66818 29946
rect 66830 29894 66882 29946
rect 24952 29588 25004 29640
rect 53840 29588 53892 29640
rect 5794 29350 5846 29402
rect 5858 29350 5910 29402
rect 5922 29350 5974 29402
rect 5986 29350 6038 29402
rect 6050 29350 6102 29402
rect 36514 29350 36566 29402
rect 36578 29350 36630 29402
rect 36642 29350 36694 29402
rect 36706 29350 36758 29402
rect 36770 29350 36822 29402
rect 67234 29350 67286 29402
rect 67298 29350 67350 29402
rect 67362 29350 67414 29402
rect 67426 29350 67478 29402
rect 67490 29350 67542 29402
rect 5134 28806 5186 28858
rect 5198 28806 5250 28858
rect 5262 28806 5314 28858
rect 5326 28806 5378 28858
rect 5390 28806 5442 28858
rect 35854 28806 35906 28858
rect 35918 28806 35970 28858
rect 35982 28806 36034 28858
rect 36046 28806 36098 28858
rect 36110 28806 36162 28858
rect 66574 28806 66626 28858
rect 66638 28806 66690 28858
rect 66702 28806 66754 28858
rect 66766 28806 66818 28858
rect 66830 28806 66882 28858
rect 5794 28262 5846 28314
rect 5858 28262 5910 28314
rect 5922 28262 5974 28314
rect 5986 28262 6038 28314
rect 6050 28262 6102 28314
rect 36514 28262 36566 28314
rect 36578 28262 36630 28314
rect 36642 28262 36694 28314
rect 36706 28262 36758 28314
rect 36770 28262 36822 28314
rect 67234 28262 67286 28314
rect 67298 28262 67350 28314
rect 67362 28262 67414 28314
rect 67426 28262 67478 28314
rect 67490 28262 67542 28314
rect 5134 27718 5186 27770
rect 5198 27718 5250 27770
rect 5262 27718 5314 27770
rect 5326 27718 5378 27770
rect 5390 27718 5442 27770
rect 35854 27718 35906 27770
rect 35918 27718 35970 27770
rect 35982 27718 36034 27770
rect 36046 27718 36098 27770
rect 36110 27718 36162 27770
rect 66574 27718 66626 27770
rect 66638 27718 66690 27770
rect 66702 27718 66754 27770
rect 66766 27718 66818 27770
rect 66830 27718 66882 27770
rect 5794 27174 5846 27226
rect 5858 27174 5910 27226
rect 5922 27174 5974 27226
rect 5986 27174 6038 27226
rect 6050 27174 6102 27226
rect 36514 27174 36566 27226
rect 36578 27174 36630 27226
rect 36642 27174 36694 27226
rect 36706 27174 36758 27226
rect 36770 27174 36822 27226
rect 67234 27174 67286 27226
rect 67298 27174 67350 27226
rect 67362 27174 67414 27226
rect 67426 27174 67478 27226
rect 67490 27174 67542 27226
rect 18788 26936 18840 26988
rect 34796 26936 34848 26988
rect 26240 26868 26292 26920
rect 46480 26868 46532 26920
rect 5134 26630 5186 26682
rect 5198 26630 5250 26682
rect 5262 26630 5314 26682
rect 5326 26630 5378 26682
rect 5390 26630 5442 26682
rect 35854 26630 35906 26682
rect 35918 26630 35970 26682
rect 35982 26630 36034 26682
rect 36046 26630 36098 26682
rect 36110 26630 36162 26682
rect 66574 26630 66626 26682
rect 66638 26630 66690 26682
rect 66702 26630 66754 26682
rect 66766 26630 66818 26682
rect 66830 26630 66882 26682
rect 5794 26086 5846 26138
rect 5858 26086 5910 26138
rect 5922 26086 5974 26138
rect 5986 26086 6038 26138
rect 6050 26086 6102 26138
rect 36514 26086 36566 26138
rect 36578 26086 36630 26138
rect 36642 26086 36694 26138
rect 36706 26086 36758 26138
rect 36770 26086 36822 26138
rect 67234 26086 67286 26138
rect 67298 26086 67350 26138
rect 67362 26086 67414 26138
rect 67426 26086 67478 26138
rect 67490 26086 67542 26138
rect 5134 25542 5186 25594
rect 5198 25542 5250 25594
rect 5262 25542 5314 25594
rect 5326 25542 5378 25594
rect 5390 25542 5442 25594
rect 35854 25542 35906 25594
rect 35918 25542 35970 25594
rect 35982 25542 36034 25594
rect 36046 25542 36098 25594
rect 36110 25542 36162 25594
rect 66574 25542 66626 25594
rect 66638 25542 66690 25594
rect 66702 25542 66754 25594
rect 66766 25542 66818 25594
rect 66830 25542 66882 25594
rect 5794 24998 5846 25050
rect 5858 24998 5910 25050
rect 5922 24998 5974 25050
rect 5986 24998 6038 25050
rect 6050 24998 6102 25050
rect 36514 24998 36566 25050
rect 36578 24998 36630 25050
rect 36642 24998 36694 25050
rect 36706 24998 36758 25050
rect 36770 24998 36822 25050
rect 67234 24998 67286 25050
rect 67298 24998 67350 25050
rect 67362 24998 67414 25050
rect 67426 24998 67478 25050
rect 67490 24998 67542 25050
rect 5134 24454 5186 24506
rect 5198 24454 5250 24506
rect 5262 24454 5314 24506
rect 5326 24454 5378 24506
rect 5390 24454 5442 24506
rect 35854 24454 35906 24506
rect 35918 24454 35970 24506
rect 35982 24454 36034 24506
rect 36046 24454 36098 24506
rect 36110 24454 36162 24506
rect 66574 24454 66626 24506
rect 66638 24454 66690 24506
rect 66702 24454 66754 24506
rect 66766 24454 66818 24506
rect 66830 24454 66882 24506
rect 21916 24148 21968 24200
rect 33324 24148 33376 24200
rect 3516 24080 3568 24132
rect 35348 24080 35400 24132
rect 5794 23910 5846 23962
rect 5858 23910 5910 23962
rect 5922 23910 5974 23962
rect 5986 23910 6038 23962
rect 6050 23910 6102 23962
rect 36514 23910 36566 23962
rect 36578 23910 36630 23962
rect 36642 23910 36694 23962
rect 36706 23910 36758 23962
rect 36770 23910 36822 23962
rect 67234 23910 67286 23962
rect 67298 23910 67350 23962
rect 67362 23910 67414 23962
rect 67426 23910 67478 23962
rect 67490 23910 67542 23962
rect 5134 23366 5186 23418
rect 5198 23366 5250 23418
rect 5262 23366 5314 23418
rect 5326 23366 5378 23418
rect 5390 23366 5442 23418
rect 35854 23366 35906 23418
rect 35918 23366 35970 23418
rect 35982 23366 36034 23418
rect 36046 23366 36098 23418
rect 36110 23366 36162 23418
rect 66574 23366 66626 23418
rect 66638 23366 66690 23418
rect 66702 23366 66754 23418
rect 66766 23366 66818 23418
rect 66830 23366 66882 23418
rect 5794 22822 5846 22874
rect 5858 22822 5910 22874
rect 5922 22822 5974 22874
rect 5986 22822 6038 22874
rect 6050 22822 6102 22874
rect 36514 22822 36566 22874
rect 36578 22822 36630 22874
rect 36642 22822 36694 22874
rect 36706 22822 36758 22874
rect 36770 22822 36822 22874
rect 67234 22822 67286 22874
rect 67298 22822 67350 22874
rect 67362 22822 67414 22874
rect 67426 22822 67478 22874
rect 67490 22822 67542 22874
rect 5134 22278 5186 22330
rect 5198 22278 5250 22330
rect 5262 22278 5314 22330
rect 5326 22278 5378 22330
rect 5390 22278 5442 22330
rect 35854 22278 35906 22330
rect 35918 22278 35970 22330
rect 35982 22278 36034 22330
rect 36046 22278 36098 22330
rect 36110 22278 36162 22330
rect 66574 22278 66626 22330
rect 66638 22278 66690 22330
rect 66702 22278 66754 22330
rect 66766 22278 66818 22330
rect 66830 22278 66882 22330
rect 5794 21734 5846 21786
rect 5858 21734 5910 21786
rect 5922 21734 5974 21786
rect 5986 21734 6038 21786
rect 6050 21734 6102 21786
rect 36514 21734 36566 21786
rect 36578 21734 36630 21786
rect 36642 21734 36694 21786
rect 36706 21734 36758 21786
rect 36770 21734 36822 21786
rect 67234 21734 67286 21786
rect 67298 21734 67350 21786
rect 67362 21734 67414 21786
rect 67426 21734 67478 21786
rect 67490 21734 67542 21786
rect 28724 21360 28776 21412
rect 39120 21360 39172 21412
rect 5134 21190 5186 21242
rect 5198 21190 5250 21242
rect 5262 21190 5314 21242
rect 5326 21190 5378 21242
rect 5390 21190 5442 21242
rect 35854 21190 35906 21242
rect 35918 21190 35970 21242
rect 35982 21190 36034 21242
rect 36046 21190 36098 21242
rect 36110 21190 36162 21242
rect 66574 21190 66626 21242
rect 66638 21190 66690 21242
rect 66702 21190 66754 21242
rect 66766 21190 66818 21242
rect 66830 21190 66882 21242
rect 5794 20646 5846 20698
rect 5858 20646 5910 20698
rect 5922 20646 5974 20698
rect 5986 20646 6038 20698
rect 6050 20646 6102 20698
rect 36514 20646 36566 20698
rect 36578 20646 36630 20698
rect 36642 20646 36694 20698
rect 36706 20646 36758 20698
rect 36770 20646 36822 20698
rect 67234 20646 67286 20698
rect 67298 20646 67350 20698
rect 67362 20646 67414 20698
rect 67426 20646 67478 20698
rect 67490 20646 67542 20698
rect 5134 20102 5186 20154
rect 5198 20102 5250 20154
rect 5262 20102 5314 20154
rect 5326 20102 5378 20154
rect 5390 20102 5442 20154
rect 35854 20102 35906 20154
rect 35918 20102 35970 20154
rect 35982 20102 36034 20154
rect 36046 20102 36098 20154
rect 36110 20102 36162 20154
rect 66574 20102 66626 20154
rect 66638 20102 66690 20154
rect 66702 20102 66754 20154
rect 66766 20102 66818 20154
rect 66830 20102 66882 20154
rect 5794 19558 5846 19610
rect 5858 19558 5910 19610
rect 5922 19558 5974 19610
rect 5986 19558 6038 19610
rect 6050 19558 6102 19610
rect 36514 19558 36566 19610
rect 36578 19558 36630 19610
rect 36642 19558 36694 19610
rect 36706 19558 36758 19610
rect 36770 19558 36822 19610
rect 67234 19558 67286 19610
rect 67298 19558 67350 19610
rect 67362 19558 67414 19610
rect 67426 19558 67478 19610
rect 67490 19558 67542 19610
rect 5134 19014 5186 19066
rect 5198 19014 5250 19066
rect 5262 19014 5314 19066
rect 5326 19014 5378 19066
rect 5390 19014 5442 19066
rect 35854 19014 35906 19066
rect 35918 19014 35970 19066
rect 35982 19014 36034 19066
rect 36046 19014 36098 19066
rect 36110 19014 36162 19066
rect 66574 19014 66626 19066
rect 66638 19014 66690 19066
rect 66702 19014 66754 19066
rect 66766 19014 66818 19066
rect 66830 19014 66882 19066
rect 5794 18470 5846 18522
rect 5858 18470 5910 18522
rect 5922 18470 5974 18522
rect 5986 18470 6038 18522
rect 6050 18470 6102 18522
rect 36514 18470 36566 18522
rect 36578 18470 36630 18522
rect 36642 18470 36694 18522
rect 36706 18470 36758 18522
rect 36770 18470 36822 18522
rect 67234 18470 67286 18522
rect 67298 18470 67350 18522
rect 67362 18470 67414 18522
rect 67426 18470 67478 18522
rect 67490 18470 67542 18522
rect 5134 17926 5186 17978
rect 5198 17926 5250 17978
rect 5262 17926 5314 17978
rect 5326 17926 5378 17978
rect 5390 17926 5442 17978
rect 35854 17926 35906 17978
rect 35918 17926 35970 17978
rect 35982 17926 36034 17978
rect 36046 17926 36098 17978
rect 36110 17926 36162 17978
rect 66574 17926 66626 17978
rect 66638 17926 66690 17978
rect 66702 17926 66754 17978
rect 66766 17926 66818 17978
rect 66830 17926 66882 17978
rect 5794 17382 5846 17434
rect 5858 17382 5910 17434
rect 5922 17382 5974 17434
rect 5986 17382 6038 17434
rect 6050 17382 6102 17434
rect 36514 17382 36566 17434
rect 36578 17382 36630 17434
rect 36642 17382 36694 17434
rect 36706 17382 36758 17434
rect 36770 17382 36822 17434
rect 67234 17382 67286 17434
rect 67298 17382 67350 17434
rect 67362 17382 67414 17434
rect 67426 17382 67478 17434
rect 67490 17382 67542 17434
rect 5134 16838 5186 16890
rect 5198 16838 5250 16890
rect 5262 16838 5314 16890
rect 5326 16838 5378 16890
rect 5390 16838 5442 16890
rect 35854 16838 35906 16890
rect 35918 16838 35970 16890
rect 35982 16838 36034 16890
rect 36046 16838 36098 16890
rect 36110 16838 36162 16890
rect 66574 16838 66626 16890
rect 66638 16838 66690 16890
rect 66702 16838 66754 16890
rect 66766 16838 66818 16890
rect 66830 16838 66882 16890
rect 5794 16294 5846 16346
rect 5858 16294 5910 16346
rect 5922 16294 5974 16346
rect 5986 16294 6038 16346
rect 6050 16294 6102 16346
rect 36514 16294 36566 16346
rect 36578 16294 36630 16346
rect 36642 16294 36694 16346
rect 36706 16294 36758 16346
rect 36770 16294 36822 16346
rect 67234 16294 67286 16346
rect 67298 16294 67350 16346
rect 67362 16294 67414 16346
rect 67426 16294 67478 16346
rect 67490 16294 67542 16346
rect 5134 15750 5186 15802
rect 5198 15750 5250 15802
rect 5262 15750 5314 15802
rect 5326 15750 5378 15802
rect 5390 15750 5442 15802
rect 35854 15750 35906 15802
rect 35918 15750 35970 15802
rect 35982 15750 36034 15802
rect 36046 15750 36098 15802
rect 36110 15750 36162 15802
rect 66574 15750 66626 15802
rect 66638 15750 66690 15802
rect 66702 15750 66754 15802
rect 66766 15750 66818 15802
rect 66830 15750 66882 15802
rect 5794 15206 5846 15258
rect 5858 15206 5910 15258
rect 5922 15206 5974 15258
rect 5986 15206 6038 15258
rect 6050 15206 6102 15258
rect 36514 15206 36566 15258
rect 36578 15206 36630 15258
rect 36642 15206 36694 15258
rect 36706 15206 36758 15258
rect 36770 15206 36822 15258
rect 67234 15206 67286 15258
rect 67298 15206 67350 15258
rect 67362 15206 67414 15258
rect 67426 15206 67478 15258
rect 67490 15206 67542 15258
rect 5134 14662 5186 14714
rect 5198 14662 5250 14714
rect 5262 14662 5314 14714
rect 5326 14662 5378 14714
rect 5390 14662 5442 14714
rect 35854 14662 35906 14714
rect 35918 14662 35970 14714
rect 35982 14662 36034 14714
rect 36046 14662 36098 14714
rect 36110 14662 36162 14714
rect 66574 14662 66626 14714
rect 66638 14662 66690 14714
rect 66702 14662 66754 14714
rect 66766 14662 66818 14714
rect 66830 14662 66882 14714
rect 27436 14492 27488 14544
rect 43352 14492 43404 14544
rect 24860 14424 24912 14476
rect 58808 14424 58860 14476
rect 5794 14118 5846 14170
rect 5858 14118 5910 14170
rect 5922 14118 5974 14170
rect 5986 14118 6038 14170
rect 6050 14118 6102 14170
rect 36514 14118 36566 14170
rect 36578 14118 36630 14170
rect 36642 14118 36694 14170
rect 36706 14118 36758 14170
rect 36770 14118 36822 14170
rect 67234 14118 67286 14170
rect 67298 14118 67350 14170
rect 67362 14118 67414 14170
rect 67426 14118 67478 14170
rect 67490 14118 67542 14170
rect 5134 13574 5186 13626
rect 5198 13574 5250 13626
rect 5262 13574 5314 13626
rect 5326 13574 5378 13626
rect 5390 13574 5442 13626
rect 35854 13574 35906 13626
rect 35918 13574 35970 13626
rect 35982 13574 36034 13626
rect 36046 13574 36098 13626
rect 36110 13574 36162 13626
rect 66574 13574 66626 13626
rect 66638 13574 66690 13626
rect 66702 13574 66754 13626
rect 66766 13574 66818 13626
rect 66830 13574 66882 13626
rect 5794 13030 5846 13082
rect 5858 13030 5910 13082
rect 5922 13030 5974 13082
rect 5986 13030 6038 13082
rect 6050 13030 6102 13082
rect 36514 13030 36566 13082
rect 36578 13030 36630 13082
rect 36642 13030 36694 13082
rect 36706 13030 36758 13082
rect 36770 13030 36822 13082
rect 67234 13030 67286 13082
rect 67298 13030 67350 13082
rect 67362 13030 67414 13082
rect 67426 13030 67478 13082
rect 67490 13030 67542 13082
rect 5134 12486 5186 12538
rect 5198 12486 5250 12538
rect 5262 12486 5314 12538
rect 5326 12486 5378 12538
rect 5390 12486 5442 12538
rect 35854 12486 35906 12538
rect 35918 12486 35970 12538
rect 35982 12486 36034 12538
rect 36046 12486 36098 12538
rect 36110 12486 36162 12538
rect 66574 12486 66626 12538
rect 66638 12486 66690 12538
rect 66702 12486 66754 12538
rect 66766 12486 66818 12538
rect 66830 12486 66882 12538
rect 28632 12180 28684 12232
rect 31024 12180 31076 12232
rect 16580 12112 16632 12164
rect 30012 12112 30064 12164
rect 17592 12044 17644 12096
rect 25320 12044 25372 12096
rect 28908 12044 28960 12096
rect 30564 12044 30616 12096
rect 5794 11942 5846 11994
rect 5858 11942 5910 11994
rect 5922 11942 5974 11994
rect 5986 11942 6038 11994
rect 6050 11942 6102 11994
rect 36514 11942 36566 11994
rect 36578 11942 36630 11994
rect 36642 11942 36694 11994
rect 36706 11942 36758 11994
rect 36770 11942 36822 11994
rect 67234 11942 67286 11994
rect 67298 11942 67350 11994
rect 67362 11942 67414 11994
rect 67426 11942 67478 11994
rect 67490 11942 67542 11994
rect 9220 11840 9272 11892
rect 22468 11840 22520 11892
rect 27252 11840 27304 11892
rect 27436 11840 27488 11892
rect 28908 11840 28960 11892
rect 32128 11840 32180 11892
rect 8484 11772 8536 11824
rect 22008 11772 22060 11824
rect 22192 11772 22244 11824
rect 23940 11772 23992 11824
rect 26424 11815 26476 11824
rect 26424 11781 26433 11815
rect 26433 11781 26467 11815
rect 26467 11781 26476 11815
rect 26424 11772 26476 11781
rect 22468 11747 22520 11756
rect 22468 11713 22477 11747
rect 22477 11713 22511 11747
rect 22511 11713 22520 11747
rect 22468 11704 22520 11713
rect 12624 11636 12676 11688
rect 24308 11704 24360 11756
rect 15016 11568 15068 11620
rect 26884 11568 26936 11620
rect 27896 11704 27948 11756
rect 28632 11747 28684 11756
rect 28632 11713 28641 11747
rect 28641 11713 28675 11747
rect 28675 11713 28684 11747
rect 28632 11704 28684 11713
rect 27436 11636 27488 11688
rect 28448 11679 28500 11688
rect 28448 11645 28457 11679
rect 28457 11645 28491 11679
rect 28491 11645 28500 11679
rect 28448 11636 28500 11645
rect 28724 11636 28776 11688
rect 29092 11704 29144 11756
rect 29184 11704 29236 11756
rect 30012 11815 30064 11824
rect 30012 11781 30021 11815
rect 30021 11781 30055 11815
rect 30055 11781 30064 11815
rect 30012 11772 30064 11781
rect 30564 11815 30616 11824
rect 30564 11781 30573 11815
rect 30573 11781 30607 11815
rect 30607 11781 30616 11815
rect 30564 11772 30616 11781
rect 33232 11815 33284 11824
rect 33232 11781 33241 11815
rect 33241 11781 33275 11815
rect 33275 11781 33284 11815
rect 33232 11772 33284 11781
rect 33876 11772 33928 11824
rect 30472 11747 30524 11756
rect 30472 11713 30481 11747
rect 30481 11713 30515 11747
rect 30515 11713 30524 11747
rect 30472 11704 30524 11713
rect 31024 11704 31076 11756
rect 33324 11747 33376 11756
rect 33324 11713 33333 11747
rect 33333 11713 33367 11747
rect 33367 11713 33376 11747
rect 33324 11704 33376 11713
rect 33968 11704 34020 11756
rect 28908 11568 28960 11620
rect 30656 11636 30708 11688
rect 33232 11636 33284 11688
rect 33048 11611 33100 11620
rect 33048 11577 33057 11611
rect 33057 11577 33091 11611
rect 33091 11577 33100 11611
rect 33048 11568 33100 11577
rect 22284 11543 22336 11552
rect 22284 11509 22293 11543
rect 22293 11509 22327 11543
rect 22327 11509 22336 11543
rect 22284 11500 22336 11509
rect 22744 11543 22796 11552
rect 22744 11509 22753 11543
rect 22753 11509 22787 11543
rect 22787 11509 22796 11543
rect 22744 11500 22796 11509
rect 23480 11543 23532 11552
rect 23480 11509 23489 11543
rect 23489 11509 23523 11543
rect 23523 11509 23532 11543
rect 23480 11500 23532 11509
rect 24216 11500 24268 11552
rect 24676 11500 24728 11552
rect 25228 11543 25280 11552
rect 25228 11509 25237 11543
rect 25237 11509 25271 11543
rect 25271 11509 25280 11543
rect 25228 11500 25280 11509
rect 25964 11500 26016 11552
rect 26516 11500 26568 11552
rect 26608 11500 26660 11552
rect 28356 11500 28408 11552
rect 29368 11500 29420 11552
rect 30288 11500 30340 11552
rect 35624 11500 35676 11552
rect 5134 11398 5186 11450
rect 5198 11398 5250 11450
rect 5262 11398 5314 11450
rect 5326 11398 5378 11450
rect 5390 11398 5442 11450
rect 35854 11398 35906 11450
rect 35918 11398 35970 11450
rect 35982 11398 36034 11450
rect 36046 11398 36098 11450
rect 36110 11398 36162 11450
rect 66574 11398 66626 11450
rect 66638 11398 66690 11450
rect 66702 11398 66754 11450
rect 66766 11398 66818 11450
rect 66830 11398 66882 11450
rect 14556 11296 14608 11348
rect 22284 11296 22336 11348
rect 22652 11296 22704 11348
rect 23296 11296 23348 11348
rect 24860 11296 24912 11348
rect 25320 11339 25372 11348
rect 25320 11305 25329 11339
rect 25329 11305 25363 11339
rect 25363 11305 25372 11339
rect 25320 11296 25372 11305
rect 26056 11339 26108 11348
rect 26056 11305 26065 11339
rect 26065 11305 26099 11339
rect 26099 11305 26108 11339
rect 26056 11296 26108 11305
rect 16212 11228 16264 11280
rect 23480 11228 23532 11280
rect 12348 11160 12400 11212
rect 22468 11160 22520 11212
rect 21732 11135 21784 11144
rect 21732 11101 21741 11135
rect 21741 11101 21775 11135
rect 21775 11101 21784 11135
rect 21732 11092 21784 11101
rect 22744 11160 22796 11212
rect 23940 11203 23992 11212
rect 23940 11169 23949 11203
rect 23949 11169 23983 11203
rect 23983 11169 23992 11203
rect 23940 11160 23992 11169
rect 24216 11203 24268 11212
rect 24216 11169 24225 11203
rect 24225 11169 24259 11203
rect 24259 11169 24268 11203
rect 24216 11160 24268 11169
rect 25228 11160 25280 11212
rect 26240 11203 26292 11212
rect 26240 11169 26249 11203
rect 26249 11169 26283 11203
rect 26283 11169 26292 11203
rect 26240 11160 26292 11169
rect 28816 11339 28868 11348
rect 28816 11305 28825 11339
rect 28825 11305 28859 11339
rect 28859 11305 28868 11339
rect 28816 11296 28868 11305
rect 38384 11296 38436 11348
rect 26884 11228 26936 11280
rect 33232 11228 33284 11280
rect 24676 11135 24728 11144
rect 24676 11101 24685 11135
rect 24685 11101 24719 11135
rect 24719 11101 24728 11135
rect 24676 11092 24728 11101
rect 24860 11135 24912 11144
rect 24860 11101 24869 11135
rect 24869 11101 24903 11135
rect 24903 11101 24912 11135
rect 24860 11092 24912 11101
rect 24952 11135 25004 11144
rect 24952 11101 24961 11135
rect 24961 11101 24995 11135
rect 24995 11101 25004 11135
rect 24952 11092 25004 11101
rect 25044 11092 25096 11144
rect 26976 11135 27028 11144
rect 26976 11101 26985 11135
rect 26985 11101 27019 11135
rect 27019 11101 27028 11135
rect 26976 11092 27028 11101
rect 28448 11135 28500 11144
rect 28448 11101 28457 11135
rect 28457 11101 28491 11135
rect 28491 11101 28500 11135
rect 28448 11092 28500 11101
rect 29184 11160 29236 11212
rect 30196 11160 30248 11212
rect 32588 11160 32640 11212
rect 31392 11135 31444 11144
rect 31392 11101 31401 11135
rect 31401 11101 31435 11135
rect 31435 11101 31444 11135
rect 31392 11092 31444 11101
rect 33416 11092 33468 11144
rect 21824 11067 21876 11076
rect 21824 11033 21833 11067
rect 21833 11033 21867 11067
rect 21867 11033 21876 11067
rect 21824 11024 21876 11033
rect 22376 11067 22428 11076
rect 22376 11033 22385 11067
rect 22385 11033 22419 11067
rect 22419 11033 22428 11067
rect 22376 11024 22428 11033
rect 17684 10956 17736 11008
rect 22744 10999 22796 11008
rect 22744 10965 22753 10999
rect 22753 10965 22787 10999
rect 22787 10965 22796 10999
rect 22744 10956 22796 10965
rect 23204 11067 23256 11076
rect 23204 11033 23213 11067
rect 23213 11033 23247 11067
rect 23247 11033 23256 11067
rect 23204 11024 23256 11033
rect 23388 11067 23440 11076
rect 23388 11033 23397 11067
rect 23397 11033 23431 11067
rect 23431 11033 23440 11067
rect 23388 11024 23440 11033
rect 23480 11024 23532 11076
rect 26884 11024 26936 11076
rect 29552 11067 29604 11076
rect 29552 11033 29561 11067
rect 29561 11033 29595 11067
rect 29595 11033 29604 11067
rect 29552 11024 29604 11033
rect 30748 11067 30800 11076
rect 30748 11033 30757 11067
rect 30757 11033 30791 11067
rect 30791 11033 30800 11067
rect 30748 11024 30800 11033
rect 33048 11024 33100 11076
rect 33968 11135 34020 11144
rect 33968 11101 33977 11135
rect 33977 11101 34011 11135
rect 34011 11101 34020 11135
rect 33968 11092 34020 11101
rect 33876 11024 33928 11076
rect 34520 11092 34572 11144
rect 35716 11160 35768 11212
rect 34796 11135 34848 11144
rect 34796 11101 34805 11135
rect 34805 11101 34839 11135
rect 34839 11101 34848 11135
rect 34796 11092 34848 11101
rect 37832 11092 37884 11144
rect 35256 11024 35308 11076
rect 24032 10956 24084 11008
rect 24124 10956 24176 11008
rect 24952 10956 25004 11008
rect 27436 10956 27488 11008
rect 5794 10854 5846 10906
rect 5858 10854 5910 10906
rect 5922 10854 5974 10906
rect 5986 10854 6038 10906
rect 6050 10854 6102 10906
rect 36514 10854 36566 10906
rect 36578 10854 36630 10906
rect 36642 10854 36694 10906
rect 36706 10854 36758 10906
rect 36770 10854 36822 10906
rect 67234 10854 67286 10906
rect 67298 10854 67350 10906
rect 67362 10854 67414 10906
rect 67426 10854 67478 10906
rect 67490 10854 67542 10906
rect 13176 10752 13228 10804
rect 13728 10684 13780 10736
rect 19340 10616 19392 10668
rect 20996 10659 21048 10668
rect 20996 10625 21005 10659
rect 21005 10625 21039 10659
rect 21039 10625 21048 10659
rect 20996 10616 21048 10625
rect 22560 10684 22612 10736
rect 15476 10548 15528 10600
rect 22928 10659 22980 10668
rect 22928 10625 22937 10659
rect 22937 10625 22971 10659
rect 22971 10625 22980 10659
rect 22928 10616 22980 10625
rect 23020 10616 23072 10668
rect 17868 10480 17920 10532
rect 21640 10523 21692 10532
rect 21640 10489 21649 10523
rect 21649 10489 21683 10523
rect 21683 10489 21692 10523
rect 21640 10480 21692 10489
rect 22192 10548 22244 10600
rect 23296 10548 23348 10600
rect 23572 10548 23624 10600
rect 24124 10591 24176 10600
rect 24124 10557 24133 10591
rect 24133 10557 24167 10591
rect 24167 10557 24176 10591
rect 24124 10548 24176 10557
rect 24400 10659 24452 10668
rect 24400 10625 24409 10659
rect 24409 10625 24443 10659
rect 24443 10625 24452 10659
rect 24400 10616 24452 10625
rect 28448 10752 28500 10804
rect 33324 10795 33376 10804
rect 33324 10761 33333 10795
rect 33333 10761 33367 10795
rect 33367 10761 33376 10795
rect 33324 10752 33376 10761
rect 26792 10684 26844 10736
rect 26056 10659 26108 10668
rect 26056 10625 26065 10659
rect 26065 10625 26099 10659
rect 26099 10625 26108 10659
rect 26056 10616 26108 10625
rect 26516 10616 26568 10668
rect 28080 10659 28132 10668
rect 28080 10625 28089 10659
rect 28089 10625 28123 10659
rect 28123 10625 28132 10659
rect 28080 10616 28132 10625
rect 26424 10591 26476 10600
rect 26424 10557 26433 10591
rect 26433 10557 26467 10591
rect 26467 10557 26476 10591
rect 26424 10548 26476 10557
rect 27068 10591 27120 10600
rect 27068 10557 27077 10591
rect 27077 10557 27111 10591
rect 27111 10557 27120 10591
rect 27068 10548 27120 10557
rect 18972 10412 19024 10464
rect 20904 10412 20956 10464
rect 21180 10455 21232 10464
rect 21180 10421 21189 10455
rect 21189 10421 21223 10455
rect 21223 10421 21232 10455
rect 21180 10412 21232 10421
rect 21456 10412 21508 10464
rect 22836 10480 22888 10532
rect 21824 10455 21876 10464
rect 21824 10421 21833 10455
rect 21833 10421 21867 10455
rect 21867 10421 21876 10455
rect 21824 10412 21876 10421
rect 23112 10455 23164 10464
rect 23112 10421 23121 10455
rect 23121 10421 23155 10455
rect 23155 10421 23164 10455
rect 23112 10412 23164 10421
rect 24768 10480 24820 10532
rect 26516 10480 26568 10532
rect 28816 10591 28868 10600
rect 28816 10557 28825 10591
rect 28825 10557 28859 10591
rect 28859 10557 28868 10591
rect 28816 10548 28868 10557
rect 30472 10591 30524 10600
rect 30472 10557 30481 10591
rect 30481 10557 30515 10591
rect 30515 10557 30524 10591
rect 30472 10548 30524 10557
rect 31392 10480 31444 10532
rect 32772 10591 32824 10600
rect 32772 10557 32781 10591
rect 32781 10557 32815 10591
rect 32815 10557 32824 10591
rect 32772 10548 32824 10557
rect 33324 10548 33376 10600
rect 34796 10591 34848 10600
rect 34796 10557 34805 10591
rect 34805 10557 34839 10591
rect 34839 10557 34848 10591
rect 34796 10548 34848 10557
rect 35532 10591 35584 10600
rect 35532 10557 35541 10591
rect 35541 10557 35575 10591
rect 35575 10557 35584 10591
rect 35532 10548 35584 10557
rect 34980 10523 35032 10532
rect 34980 10489 34989 10523
rect 34989 10489 35023 10523
rect 35023 10489 35032 10523
rect 34980 10480 35032 10489
rect 24124 10412 24176 10464
rect 25228 10412 25280 10464
rect 27528 10412 27580 10464
rect 27620 10412 27672 10464
rect 28264 10455 28316 10464
rect 28264 10421 28273 10455
rect 28273 10421 28307 10455
rect 28307 10421 28316 10455
rect 28264 10412 28316 10421
rect 29000 10455 29052 10464
rect 29000 10421 29009 10455
rect 29009 10421 29043 10455
rect 29043 10421 29052 10455
rect 29000 10412 29052 10421
rect 29276 10412 29328 10464
rect 29552 10412 29604 10464
rect 31484 10455 31536 10464
rect 31484 10421 31493 10455
rect 31493 10421 31527 10455
rect 31527 10421 31536 10455
rect 31484 10412 31536 10421
rect 31576 10412 31628 10464
rect 33140 10412 33192 10464
rect 5134 10310 5186 10362
rect 5198 10310 5250 10362
rect 5262 10310 5314 10362
rect 5326 10310 5378 10362
rect 5390 10310 5442 10362
rect 35854 10310 35906 10362
rect 35918 10310 35970 10362
rect 35982 10310 36034 10362
rect 36046 10310 36098 10362
rect 36110 10310 36162 10362
rect 66574 10310 66626 10362
rect 66638 10310 66690 10362
rect 66702 10310 66754 10362
rect 66766 10310 66818 10362
rect 66830 10310 66882 10362
rect 14924 10208 14976 10260
rect 23112 10208 23164 10260
rect 24032 10208 24084 10260
rect 27068 10208 27120 10260
rect 30380 10208 30432 10260
rect 17408 10140 17460 10192
rect 20628 10140 20680 10192
rect 31484 10140 31536 10192
rect 19156 10072 19208 10124
rect 19616 10047 19668 10056
rect 19616 10013 19625 10047
rect 19625 10013 19659 10047
rect 19659 10013 19668 10047
rect 19616 10004 19668 10013
rect 19708 10004 19760 10056
rect 20444 10047 20496 10056
rect 20444 10013 20453 10047
rect 20453 10013 20487 10047
rect 20487 10013 20496 10047
rect 20444 10004 20496 10013
rect 19800 9936 19852 9988
rect 22744 10072 22796 10124
rect 23204 10072 23256 10124
rect 26332 10072 26384 10124
rect 27712 10072 27764 10124
rect 29552 10115 29604 10124
rect 29552 10081 29561 10115
rect 29561 10081 29595 10115
rect 29595 10081 29604 10115
rect 29552 10072 29604 10081
rect 21640 10004 21692 10056
rect 23296 10047 23348 10056
rect 23296 10013 23305 10047
rect 23305 10013 23339 10047
rect 23339 10013 23348 10047
rect 23296 10004 23348 10013
rect 24492 10047 24544 10056
rect 24492 10013 24501 10047
rect 24501 10013 24535 10047
rect 24535 10013 24544 10047
rect 24492 10004 24544 10013
rect 27436 10004 27488 10056
rect 27988 10047 28040 10056
rect 27988 10013 27997 10047
rect 27997 10013 28031 10047
rect 28031 10013 28040 10047
rect 27988 10004 28040 10013
rect 23756 9936 23808 9988
rect 27620 9936 27672 9988
rect 29828 10004 29880 10056
rect 31116 10047 31168 10056
rect 31116 10013 31125 10047
rect 31125 10013 31159 10047
rect 31159 10013 31168 10047
rect 31116 10004 31168 10013
rect 32956 10140 33008 10192
rect 33600 10183 33652 10192
rect 33600 10149 33609 10183
rect 33609 10149 33643 10183
rect 33643 10149 33652 10183
rect 33600 10140 33652 10149
rect 31944 10047 31996 10056
rect 31944 10013 31953 10047
rect 31953 10013 31987 10047
rect 31987 10013 31996 10047
rect 31944 10004 31996 10013
rect 33416 10047 33468 10056
rect 33416 10013 33425 10047
rect 33425 10013 33459 10047
rect 33459 10013 33468 10047
rect 33416 10004 33468 10013
rect 34244 10047 34296 10056
rect 34244 10013 34253 10047
rect 34253 10013 34287 10047
rect 34287 10013 34296 10047
rect 34244 10004 34296 10013
rect 34888 10047 34940 10056
rect 34888 10013 34897 10047
rect 34897 10013 34931 10047
rect 34931 10013 34940 10047
rect 34888 10004 34940 10013
rect 36360 10004 36412 10056
rect 36636 10047 36688 10056
rect 36636 10013 36645 10047
rect 36645 10013 36679 10047
rect 36679 10013 36688 10047
rect 36636 10004 36688 10013
rect 37648 10004 37700 10056
rect 19432 9911 19484 9920
rect 19432 9877 19441 9911
rect 19441 9877 19475 9911
rect 19475 9877 19484 9911
rect 19432 9868 19484 9877
rect 19524 9868 19576 9920
rect 20812 9911 20864 9920
rect 20812 9877 20821 9911
rect 20821 9877 20855 9911
rect 20855 9877 20864 9911
rect 20812 9868 20864 9877
rect 21548 9911 21600 9920
rect 21548 9877 21557 9911
rect 21557 9877 21591 9911
rect 21591 9877 21600 9911
rect 21548 9868 21600 9877
rect 22100 9868 22152 9920
rect 23020 9868 23072 9920
rect 23296 9911 23348 9920
rect 23296 9877 23305 9911
rect 23305 9877 23339 9911
rect 23339 9877 23348 9911
rect 23296 9868 23348 9877
rect 23480 9868 23532 9920
rect 24584 9868 24636 9920
rect 24676 9868 24728 9920
rect 25136 9868 25188 9920
rect 27252 9868 27304 9920
rect 27528 9868 27580 9920
rect 28724 9868 28776 9920
rect 30012 9868 30064 9920
rect 30564 9911 30616 9920
rect 30564 9877 30573 9911
rect 30573 9877 30607 9911
rect 30607 9877 30616 9911
rect 30564 9868 30616 9877
rect 31852 9868 31904 9920
rect 32864 9911 32916 9920
rect 32864 9877 32873 9911
rect 32873 9877 32907 9911
rect 32907 9877 32916 9911
rect 32864 9868 32916 9877
rect 34336 9911 34388 9920
rect 34336 9877 34345 9911
rect 34345 9877 34379 9911
rect 34379 9877 34388 9911
rect 34336 9868 34388 9877
rect 35900 9911 35952 9920
rect 35900 9877 35909 9911
rect 35909 9877 35943 9911
rect 35943 9877 35952 9911
rect 35900 9868 35952 9877
rect 5794 9766 5846 9818
rect 5858 9766 5910 9818
rect 5922 9766 5974 9818
rect 5986 9766 6038 9818
rect 6050 9766 6102 9818
rect 36514 9766 36566 9818
rect 36578 9766 36630 9818
rect 36642 9766 36694 9818
rect 36706 9766 36758 9818
rect 36770 9766 36822 9818
rect 67234 9766 67286 9818
rect 67298 9766 67350 9818
rect 67362 9766 67414 9818
rect 67426 9766 67478 9818
rect 67490 9766 67542 9818
rect 13268 9664 13320 9716
rect 16580 9664 16632 9716
rect 21732 9664 21784 9716
rect 26424 9664 26476 9716
rect 18788 9596 18840 9648
rect 21088 9596 21140 9648
rect 19432 9528 19484 9580
rect 18512 9460 18564 9512
rect 22560 9571 22612 9580
rect 22560 9537 22569 9571
rect 22569 9537 22603 9571
rect 22603 9537 22612 9571
rect 22560 9528 22612 9537
rect 23388 9528 23440 9580
rect 25596 9596 25648 9648
rect 31944 9664 31996 9716
rect 34888 9664 34940 9716
rect 28080 9596 28132 9648
rect 25136 9571 25188 9580
rect 25136 9537 25145 9571
rect 25145 9537 25179 9571
rect 25179 9537 25188 9571
rect 25136 9528 25188 9537
rect 25320 9571 25372 9580
rect 25320 9537 25329 9571
rect 25329 9537 25363 9571
rect 25363 9537 25372 9571
rect 25320 9528 25372 9537
rect 26608 9571 26660 9580
rect 26608 9537 26617 9571
rect 26617 9537 26651 9571
rect 26651 9537 26660 9571
rect 26608 9528 26660 9537
rect 26884 9528 26936 9580
rect 19892 9503 19944 9512
rect 19892 9469 19901 9503
rect 19901 9469 19935 9503
rect 19935 9469 19944 9503
rect 19892 9460 19944 9469
rect 20720 9503 20772 9512
rect 20720 9469 20729 9503
rect 20729 9469 20763 9503
rect 20763 9469 20772 9503
rect 20720 9460 20772 9469
rect 21732 9460 21784 9512
rect 22744 9460 22796 9512
rect 19248 9392 19300 9444
rect 20260 9392 20312 9444
rect 22008 9392 22060 9444
rect 25964 9503 26016 9512
rect 25964 9469 25973 9503
rect 25973 9469 26007 9503
rect 26007 9469 26016 9503
rect 25964 9460 26016 9469
rect 27896 9528 27948 9580
rect 31668 9596 31720 9648
rect 35624 9596 35676 9648
rect 28448 9528 28500 9580
rect 30748 9528 30800 9580
rect 18604 9367 18656 9376
rect 18604 9333 18613 9367
rect 18613 9333 18647 9367
rect 18647 9333 18656 9367
rect 18604 9324 18656 9333
rect 18696 9324 18748 9376
rect 20812 9324 20864 9376
rect 23480 9324 23532 9376
rect 23756 9392 23808 9444
rect 24216 9392 24268 9444
rect 24768 9392 24820 9444
rect 28632 9503 28684 9512
rect 28632 9469 28641 9503
rect 28641 9469 28675 9503
rect 28675 9469 28684 9503
rect 28632 9460 28684 9469
rect 30104 9503 30156 9512
rect 30104 9469 30113 9503
rect 30113 9469 30147 9503
rect 30147 9469 30156 9503
rect 30104 9460 30156 9469
rect 30196 9460 30248 9512
rect 27896 9392 27948 9444
rect 32404 9528 32456 9580
rect 34336 9528 34388 9580
rect 34704 9528 34756 9580
rect 37372 9528 37424 9580
rect 37832 9571 37884 9580
rect 37832 9537 37841 9571
rect 37841 9537 37875 9571
rect 37875 9537 37884 9571
rect 37832 9528 37884 9537
rect 31208 9503 31260 9512
rect 31208 9469 31217 9503
rect 31217 9469 31251 9503
rect 31251 9469 31260 9503
rect 31208 9460 31260 9469
rect 31576 9460 31628 9512
rect 34888 9460 34940 9512
rect 23664 9367 23716 9376
rect 23664 9333 23673 9367
rect 23673 9333 23707 9367
rect 23707 9333 23716 9367
rect 23664 9324 23716 9333
rect 23848 9324 23900 9376
rect 25872 9367 25924 9376
rect 25872 9333 25881 9367
rect 25881 9333 25915 9367
rect 25915 9333 25924 9367
rect 25872 9324 25924 9333
rect 27344 9324 27396 9376
rect 27804 9324 27856 9376
rect 29460 9324 29512 9376
rect 30196 9367 30248 9376
rect 30196 9333 30205 9367
rect 30205 9333 30239 9367
rect 30239 9333 30248 9367
rect 30196 9324 30248 9333
rect 30840 9324 30892 9376
rect 34336 9392 34388 9444
rect 40040 9460 40092 9512
rect 37740 9435 37792 9444
rect 37740 9401 37749 9435
rect 37749 9401 37783 9435
rect 37783 9401 37792 9435
rect 37740 9392 37792 9401
rect 31484 9324 31536 9376
rect 32312 9324 32364 9376
rect 32680 9324 32732 9376
rect 34060 9367 34112 9376
rect 34060 9333 34069 9367
rect 34069 9333 34103 9367
rect 34103 9333 34112 9367
rect 34060 9324 34112 9333
rect 34888 9367 34940 9376
rect 34888 9333 34897 9367
rect 34897 9333 34931 9367
rect 34931 9333 34940 9367
rect 34888 9324 34940 9333
rect 37188 9324 37240 9376
rect 38016 9367 38068 9376
rect 38016 9333 38025 9367
rect 38025 9333 38059 9367
rect 38059 9333 38068 9367
rect 38016 9324 38068 9333
rect 38200 9367 38252 9376
rect 38200 9333 38209 9367
rect 38209 9333 38243 9367
rect 38243 9333 38252 9367
rect 38200 9324 38252 9333
rect 5134 9222 5186 9274
rect 5198 9222 5250 9274
rect 5262 9222 5314 9274
rect 5326 9222 5378 9274
rect 5390 9222 5442 9274
rect 35854 9222 35906 9274
rect 35918 9222 35970 9274
rect 35982 9222 36034 9274
rect 36046 9222 36098 9274
rect 36110 9222 36162 9274
rect 66574 9222 66626 9274
rect 66638 9222 66690 9274
rect 66702 9222 66754 9274
rect 66766 9222 66818 9274
rect 66830 9222 66882 9274
rect 11704 9163 11756 9172
rect 11704 9129 11713 9163
rect 11713 9129 11747 9163
rect 11747 9129 11756 9163
rect 11704 9120 11756 9129
rect 15568 9120 15620 9172
rect 10600 9052 10652 9104
rect 19156 9120 19208 9172
rect 20996 9120 21048 9172
rect 24676 9120 24728 9172
rect 27436 9120 27488 9172
rect 19340 9052 19392 9104
rect 21640 9052 21692 9104
rect 24400 9052 24452 9104
rect 28632 9163 28684 9172
rect 28632 9129 28641 9163
rect 28641 9129 28675 9163
rect 28675 9129 28684 9163
rect 28632 9120 28684 9129
rect 28816 9120 28868 9172
rect 29920 9120 29972 9172
rect 32404 9120 32456 9172
rect 32772 9120 32824 9172
rect 34520 9120 34572 9172
rect 15936 8984 15988 9036
rect 18328 8984 18380 9036
rect 19156 8984 19208 9036
rect 21272 8984 21324 9036
rect 11244 8916 11296 8968
rect 8852 8848 8904 8900
rect 18420 8916 18472 8968
rect 18880 8916 18932 8968
rect 19616 8916 19668 8968
rect 19800 8916 19852 8968
rect 20168 8916 20220 8968
rect 20444 8959 20496 8968
rect 20444 8925 20453 8959
rect 20453 8925 20487 8959
rect 20487 8925 20496 8959
rect 20444 8916 20496 8925
rect 21456 8916 21508 8968
rect 21824 8959 21876 8968
rect 21824 8925 21833 8959
rect 21833 8925 21867 8959
rect 21867 8925 21876 8959
rect 21824 8916 21876 8925
rect 16672 8848 16724 8900
rect 3240 8780 3292 8832
rect 18236 8780 18288 8832
rect 19800 8780 19852 8832
rect 21364 8780 21416 8832
rect 22008 8780 22060 8832
rect 22560 8959 22612 8968
rect 22560 8925 22569 8959
rect 22569 8925 22603 8959
rect 22603 8925 22612 8959
rect 22560 8916 22612 8925
rect 22652 8959 22704 8968
rect 22652 8925 22661 8959
rect 22661 8925 22695 8959
rect 22695 8925 22704 8959
rect 22652 8916 22704 8925
rect 22836 8916 22888 8968
rect 23296 8916 23348 8968
rect 23756 8959 23808 8968
rect 23756 8925 23765 8959
rect 23765 8925 23799 8959
rect 23799 8925 23808 8959
rect 23756 8916 23808 8925
rect 23020 8891 23072 8900
rect 23020 8857 23029 8891
rect 23029 8857 23063 8891
rect 23063 8857 23072 8891
rect 23020 8848 23072 8857
rect 23112 8848 23164 8900
rect 24216 8916 24268 8968
rect 24768 8959 24820 8968
rect 24768 8925 24777 8959
rect 24777 8925 24811 8959
rect 24811 8925 24820 8959
rect 24768 8916 24820 8925
rect 25320 8959 25372 8968
rect 25320 8925 25329 8959
rect 25329 8925 25363 8959
rect 25363 8925 25372 8959
rect 25320 8916 25372 8925
rect 31576 9052 31628 9104
rect 31668 9052 31720 9104
rect 34428 9052 34480 9104
rect 27804 8984 27856 9036
rect 30288 8984 30340 9036
rect 23940 8848 23992 8900
rect 28080 8916 28132 8968
rect 29552 8916 29604 8968
rect 30564 8916 30616 8968
rect 33048 8984 33100 9036
rect 34612 9027 34664 9036
rect 34612 8993 34621 9027
rect 34621 8993 34655 9027
rect 34655 8993 34664 9027
rect 34612 8984 34664 8993
rect 31576 8916 31628 8968
rect 33968 8959 34020 8968
rect 33968 8925 33977 8959
rect 33977 8925 34011 8959
rect 34011 8925 34020 8959
rect 33968 8916 34020 8925
rect 35808 9120 35860 9172
rect 37740 9120 37792 9172
rect 34980 9052 35032 9104
rect 36176 9052 36228 9104
rect 22192 8780 22244 8832
rect 22284 8823 22336 8832
rect 22284 8789 22293 8823
rect 22293 8789 22327 8823
rect 22327 8789 22336 8823
rect 22284 8780 22336 8789
rect 22836 8780 22888 8832
rect 24216 8780 24268 8832
rect 25136 8823 25188 8832
rect 25136 8789 25145 8823
rect 25145 8789 25179 8823
rect 25179 8789 25188 8823
rect 25136 8780 25188 8789
rect 25872 8780 25924 8832
rect 26240 8823 26292 8832
rect 26240 8789 26249 8823
rect 26249 8789 26283 8823
rect 26283 8789 26292 8823
rect 26240 8780 26292 8789
rect 28264 8848 28316 8900
rect 30932 8891 30984 8900
rect 30932 8857 30941 8891
rect 30941 8857 30975 8891
rect 30975 8857 30984 8891
rect 30932 8848 30984 8857
rect 31668 8891 31720 8900
rect 31668 8857 31677 8891
rect 31677 8857 31711 8891
rect 31711 8857 31720 8891
rect 31668 8848 31720 8857
rect 32404 8848 32456 8900
rect 33048 8848 33100 8900
rect 38752 8984 38804 9036
rect 35164 8959 35216 8968
rect 35164 8925 35173 8959
rect 35173 8925 35207 8959
rect 35207 8925 35216 8959
rect 35164 8916 35216 8925
rect 35256 8959 35308 8968
rect 35256 8925 35265 8959
rect 35265 8925 35299 8959
rect 35299 8925 35308 8959
rect 35256 8916 35308 8925
rect 35808 8959 35860 8968
rect 35808 8925 35817 8959
rect 35817 8925 35851 8959
rect 35851 8925 35860 8959
rect 35808 8916 35860 8925
rect 35072 8891 35124 8900
rect 35072 8857 35081 8891
rect 35081 8857 35115 8891
rect 35115 8857 35124 8891
rect 35072 8848 35124 8857
rect 36360 8916 36412 8968
rect 37004 8916 37056 8968
rect 38200 8959 38252 8968
rect 38200 8925 38209 8959
rect 38209 8925 38243 8959
rect 38243 8925 38252 8959
rect 38200 8916 38252 8925
rect 38660 8848 38712 8900
rect 26608 8780 26660 8832
rect 28172 8780 28224 8832
rect 31116 8823 31168 8832
rect 31116 8789 31125 8823
rect 31125 8789 31159 8823
rect 31159 8789 31168 8823
rect 31116 8780 31168 8789
rect 33232 8780 33284 8832
rect 33508 8780 33560 8832
rect 34152 8780 34204 8832
rect 36912 8780 36964 8832
rect 37464 8780 37516 8832
rect 39764 8780 39816 8832
rect 5794 8678 5846 8730
rect 5858 8678 5910 8730
rect 5922 8678 5974 8730
rect 5986 8678 6038 8730
rect 6050 8678 6102 8730
rect 36514 8678 36566 8730
rect 36578 8678 36630 8730
rect 36642 8678 36694 8730
rect 36706 8678 36758 8730
rect 36770 8678 36822 8730
rect 67234 8678 67286 8730
rect 67298 8678 67350 8730
rect 67362 8678 67414 8730
rect 67426 8678 67478 8730
rect 67490 8678 67542 8730
rect 11704 8576 11756 8628
rect 18696 8576 18748 8628
rect 18880 8619 18932 8628
rect 18880 8585 18889 8619
rect 18889 8585 18923 8619
rect 18923 8585 18932 8619
rect 18880 8576 18932 8585
rect 18144 8551 18196 8560
rect 18144 8517 18153 8551
rect 18153 8517 18187 8551
rect 18187 8517 18196 8551
rect 18144 8508 18196 8517
rect 14004 8440 14056 8492
rect 14648 8372 14700 8424
rect 16856 8372 16908 8424
rect 3976 8304 4028 8356
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 18052 8440 18104 8492
rect 21364 8576 21416 8628
rect 22560 8576 22612 8628
rect 22836 8576 22888 8628
rect 23388 8576 23440 8628
rect 24308 8576 24360 8628
rect 29920 8576 29972 8628
rect 30104 8576 30156 8628
rect 21548 8508 21600 8560
rect 21732 8508 21784 8560
rect 22652 8508 22704 8560
rect 23848 8508 23900 8560
rect 24216 8551 24268 8560
rect 24216 8517 24225 8551
rect 24225 8517 24259 8551
rect 24259 8517 24268 8551
rect 24216 8508 24268 8517
rect 25872 8508 25924 8560
rect 26240 8508 26292 8560
rect 19984 8440 20036 8492
rect 22284 8440 22336 8492
rect 22560 8483 22612 8492
rect 22560 8449 22569 8483
rect 22569 8449 22603 8483
rect 22603 8449 22612 8483
rect 22560 8440 22612 8449
rect 22836 8483 22888 8492
rect 22836 8449 22845 8483
rect 22845 8449 22879 8483
rect 22879 8449 22888 8483
rect 22836 8440 22888 8449
rect 26424 8440 26476 8492
rect 27528 8508 27580 8560
rect 17040 8372 17092 8424
rect 15200 8236 15252 8288
rect 17868 8236 17920 8288
rect 18144 8304 18196 8356
rect 20260 8415 20312 8424
rect 20260 8381 20269 8415
rect 20269 8381 20303 8415
rect 20303 8381 20312 8415
rect 20260 8372 20312 8381
rect 20352 8372 20404 8424
rect 18880 8304 18932 8356
rect 22376 8304 22428 8356
rect 25964 8372 26016 8424
rect 26608 8415 26660 8424
rect 26608 8381 26617 8415
rect 26617 8381 26651 8415
rect 26651 8381 26660 8415
rect 26608 8372 26660 8381
rect 27804 8440 27856 8492
rect 28540 8440 28592 8492
rect 29460 8483 29512 8492
rect 29460 8449 29469 8483
rect 29469 8449 29503 8483
rect 29503 8449 29512 8483
rect 29460 8440 29512 8449
rect 27160 8372 27212 8424
rect 27712 8415 27764 8424
rect 27712 8381 27721 8415
rect 27721 8381 27755 8415
rect 27755 8381 27764 8415
rect 27712 8372 27764 8381
rect 28448 8372 28500 8424
rect 25780 8304 25832 8356
rect 26884 8304 26936 8356
rect 29460 8304 29512 8356
rect 30196 8508 30248 8560
rect 30656 8576 30708 8628
rect 32220 8576 32272 8628
rect 35256 8576 35308 8628
rect 35900 8576 35952 8628
rect 31300 8508 31352 8560
rect 29920 8415 29972 8424
rect 29920 8381 29929 8415
rect 29929 8381 29963 8415
rect 29963 8381 29972 8415
rect 29920 8372 29972 8381
rect 32036 8508 32088 8560
rect 33692 8508 33744 8560
rect 35072 8508 35124 8560
rect 35440 8508 35492 8560
rect 37556 8508 37608 8560
rect 32220 8440 32272 8492
rect 33784 8440 33836 8492
rect 36268 8440 36320 8492
rect 36728 8440 36780 8492
rect 39764 8483 39816 8492
rect 39764 8449 39773 8483
rect 39773 8449 39807 8483
rect 39807 8449 39816 8483
rect 39764 8440 39816 8449
rect 32404 8372 32456 8424
rect 33232 8372 33284 8424
rect 34612 8415 34664 8424
rect 34612 8381 34621 8415
rect 34621 8381 34655 8415
rect 34655 8381 34664 8415
rect 34612 8372 34664 8381
rect 35164 8415 35216 8424
rect 35164 8381 35173 8415
rect 35173 8381 35207 8415
rect 35207 8381 35216 8415
rect 35164 8372 35216 8381
rect 35716 8372 35768 8424
rect 30932 8304 30984 8356
rect 19340 8236 19392 8288
rect 22008 8236 22060 8288
rect 22284 8236 22336 8288
rect 23112 8236 23164 8288
rect 23848 8236 23900 8288
rect 26056 8279 26108 8288
rect 26056 8245 26065 8279
rect 26065 8245 26099 8279
rect 26099 8245 26108 8279
rect 26056 8236 26108 8245
rect 26332 8236 26384 8288
rect 28080 8236 28132 8288
rect 28264 8236 28316 8288
rect 29644 8236 29696 8288
rect 37280 8304 37332 8356
rect 39212 8347 39264 8356
rect 39212 8313 39221 8347
rect 39221 8313 39255 8347
rect 39255 8313 39264 8347
rect 39212 8304 39264 8313
rect 39396 8372 39448 8424
rect 39856 8304 39908 8356
rect 41420 8304 41472 8356
rect 31024 8236 31076 8288
rect 31300 8236 31352 8288
rect 31760 8279 31812 8288
rect 31760 8245 31769 8279
rect 31769 8245 31803 8279
rect 31803 8245 31812 8279
rect 31760 8236 31812 8245
rect 32496 8279 32548 8288
rect 32496 8245 32505 8279
rect 32505 8245 32539 8279
rect 32539 8245 32548 8279
rect 32496 8236 32548 8245
rect 32680 8279 32732 8288
rect 32680 8245 32689 8279
rect 32689 8245 32723 8279
rect 32723 8245 32732 8279
rect 32680 8236 32732 8245
rect 32956 8236 33008 8288
rect 33140 8236 33192 8288
rect 35532 8236 35584 8288
rect 36728 8236 36780 8288
rect 39028 8236 39080 8288
rect 5134 8134 5186 8186
rect 5198 8134 5250 8186
rect 5262 8134 5314 8186
rect 5326 8134 5378 8186
rect 5390 8134 5442 8186
rect 35854 8134 35906 8186
rect 35918 8134 35970 8186
rect 35982 8134 36034 8186
rect 36046 8134 36098 8186
rect 36110 8134 36162 8186
rect 66574 8134 66626 8186
rect 66638 8134 66690 8186
rect 66702 8134 66754 8186
rect 66766 8134 66818 8186
rect 66830 8134 66882 8186
rect 10508 8032 10560 8084
rect 16580 8032 16632 8084
rect 12716 7964 12768 8016
rect 15660 8007 15712 8016
rect 15660 7973 15669 8007
rect 15669 7973 15703 8007
rect 15703 7973 15712 8007
rect 15660 7964 15712 7973
rect 19708 7964 19760 8016
rect 19984 8075 20036 8084
rect 19984 8041 19993 8075
rect 19993 8041 20027 8075
rect 20027 8041 20036 8075
rect 19984 8032 20036 8041
rect 21088 8032 21140 8084
rect 21272 8075 21324 8084
rect 21272 8041 21281 8075
rect 21281 8041 21315 8075
rect 21315 8041 21324 8075
rect 21272 8032 21324 8041
rect 20260 7964 20312 8016
rect 25136 8032 25188 8084
rect 25412 8032 25464 8084
rect 25688 8032 25740 8084
rect 27160 8032 27212 8084
rect 27344 8075 27396 8084
rect 27344 8041 27353 8075
rect 27353 8041 27387 8075
rect 27387 8041 27396 8075
rect 27344 8032 27396 8041
rect 29920 8032 29972 8084
rect 23480 7964 23532 8016
rect 16304 7896 16356 7948
rect 16488 7896 16540 7948
rect 18788 7896 18840 7948
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 14372 7760 14424 7812
rect 15200 7871 15252 7880
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 15844 7760 15896 7812
rect 14464 7692 14516 7744
rect 15016 7692 15068 7744
rect 17132 7871 17184 7880
rect 17132 7837 17141 7871
rect 17141 7837 17175 7871
rect 17175 7837 17184 7871
rect 17132 7828 17184 7837
rect 22008 7939 22060 7948
rect 22008 7905 22017 7939
rect 22017 7905 22051 7939
rect 22051 7905 22060 7939
rect 22008 7896 22060 7905
rect 22376 7896 22428 7948
rect 23572 7896 23624 7948
rect 25872 7964 25924 8016
rect 16488 7760 16540 7812
rect 19156 7828 19208 7880
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 20168 7871 20220 7880
rect 20168 7837 20177 7871
rect 20177 7837 20211 7871
rect 20211 7837 20220 7871
rect 20168 7828 20220 7837
rect 20260 7871 20312 7880
rect 20260 7837 20269 7871
rect 20269 7837 20303 7871
rect 20303 7837 20312 7871
rect 20260 7828 20312 7837
rect 21180 7828 21232 7880
rect 24768 7896 24820 7948
rect 26056 7896 26108 7948
rect 26884 7896 26936 7948
rect 31116 8032 31168 8084
rect 33692 8032 33744 8084
rect 31760 7964 31812 8016
rect 33416 7964 33468 8016
rect 35164 8032 35216 8084
rect 19708 7760 19760 7812
rect 21364 7760 21416 7812
rect 18512 7735 18564 7744
rect 18512 7701 18521 7735
rect 18521 7701 18555 7735
rect 18555 7701 18564 7735
rect 18512 7692 18564 7701
rect 18696 7692 18748 7744
rect 21548 7692 21600 7744
rect 22468 7760 22520 7812
rect 23848 7760 23900 7812
rect 25320 7828 25372 7880
rect 25688 7828 25740 7880
rect 25780 7871 25832 7880
rect 25780 7837 25789 7871
rect 25789 7837 25823 7871
rect 25823 7837 25832 7871
rect 25780 7828 25832 7837
rect 26700 7828 26752 7880
rect 27068 7828 27120 7880
rect 28908 7871 28960 7880
rect 28908 7837 28917 7871
rect 28917 7837 28951 7871
rect 28951 7837 28960 7871
rect 28908 7828 28960 7837
rect 31668 7896 31720 7948
rect 32956 7896 33008 7948
rect 33600 7896 33652 7948
rect 35256 7896 35308 7948
rect 30472 7871 30524 7880
rect 30472 7837 30481 7871
rect 30481 7837 30515 7871
rect 30515 7837 30524 7871
rect 30472 7828 30524 7837
rect 30656 7871 30708 7880
rect 30656 7837 30665 7871
rect 30665 7837 30699 7871
rect 30699 7837 30708 7871
rect 30656 7828 30708 7837
rect 31116 7828 31168 7880
rect 30288 7760 30340 7812
rect 34244 7828 34296 7880
rect 35164 7828 35216 7880
rect 35624 7871 35676 7880
rect 35624 7837 35633 7871
rect 35633 7837 35667 7871
rect 35667 7837 35676 7871
rect 35624 7828 35676 7837
rect 37832 7896 37884 7948
rect 37924 7896 37976 7948
rect 41420 7939 41472 7948
rect 41420 7905 41429 7939
rect 41429 7905 41463 7939
rect 41463 7905 41472 7939
rect 41420 7896 41472 7905
rect 38844 7871 38896 7880
rect 38844 7837 38853 7871
rect 38853 7837 38887 7871
rect 38887 7837 38896 7871
rect 38844 7828 38896 7837
rect 46480 7828 46532 7880
rect 32404 7803 32456 7812
rect 32404 7769 32413 7803
rect 32413 7769 32447 7803
rect 32447 7769 32456 7803
rect 32404 7760 32456 7769
rect 24032 7692 24084 7744
rect 25320 7692 25372 7744
rect 25780 7692 25832 7744
rect 25964 7692 26016 7744
rect 26608 7735 26660 7744
rect 26608 7701 26617 7735
rect 26617 7701 26651 7735
rect 26651 7701 26660 7735
rect 26608 7692 26660 7701
rect 26884 7692 26936 7744
rect 27160 7692 27212 7744
rect 29092 7692 29144 7744
rect 29736 7692 29788 7744
rect 31024 7692 31076 7744
rect 33876 7760 33928 7812
rect 34336 7760 34388 7812
rect 35900 7760 35952 7812
rect 36728 7760 36780 7812
rect 37924 7760 37976 7812
rect 41236 7760 41288 7812
rect 41604 7803 41656 7812
rect 41604 7769 41613 7803
rect 41613 7769 41647 7803
rect 41647 7769 41656 7803
rect 41604 7760 41656 7769
rect 34520 7692 34572 7744
rect 38292 7692 38344 7744
rect 39120 7692 39172 7744
rect 40132 7692 40184 7744
rect 41788 7692 41840 7744
rect 5794 7590 5846 7642
rect 5858 7590 5910 7642
rect 5922 7590 5974 7642
rect 5986 7590 6038 7642
rect 6050 7590 6102 7642
rect 36514 7590 36566 7642
rect 36578 7590 36630 7642
rect 36642 7590 36694 7642
rect 36706 7590 36758 7642
rect 36770 7590 36822 7642
rect 67234 7590 67286 7642
rect 67298 7590 67350 7642
rect 67362 7590 67414 7642
rect 67426 7590 67478 7642
rect 67490 7590 67542 7642
rect 15292 7488 15344 7540
rect 15936 7531 15988 7540
rect 15936 7497 15945 7531
rect 15945 7497 15979 7531
rect 15979 7497 15988 7531
rect 15936 7488 15988 7497
rect 16120 7488 16172 7540
rect 18604 7488 18656 7540
rect 20996 7488 21048 7540
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 8944 7420 8996 7472
rect 6736 7352 6788 7404
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 9128 7284 9180 7336
rect 13360 7327 13412 7336
rect 13360 7293 13369 7327
rect 13369 7293 13403 7327
rect 13403 7293 13412 7327
rect 13360 7284 13412 7293
rect 7564 7216 7616 7268
rect 12072 7216 12124 7268
rect 12164 7216 12216 7268
rect 14372 7395 14424 7404
rect 14372 7361 14381 7395
rect 14381 7361 14415 7395
rect 14415 7361 14424 7395
rect 14372 7352 14424 7361
rect 15384 7420 15436 7472
rect 19524 7420 19576 7472
rect 15108 7352 15160 7404
rect 16488 7352 16540 7404
rect 16580 7395 16632 7404
rect 16580 7361 16589 7395
rect 16589 7361 16623 7395
rect 16623 7361 16632 7395
rect 16580 7352 16632 7361
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 15200 7284 15252 7336
rect 15292 7327 15344 7336
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 15384 7284 15436 7336
rect 17868 7395 17920 7404
rect 17868 7361 17877 7395
rect 17877 7361 17911 7395
rect 17911 7361 17920 7395
rect 17868 7352 17920 7361
rect 19340 7352 19392 7404
rect 20168 7352 20220 7404
rect 21456 7420 21508 7472
rect 18788 7284 18840 7336
rect 18972 7327 19024 7336
rect 18972 7293 18981 7327
rect 18981 7293 19015 7327
rect 19015 7293 19024 7327
rect 18972 7284 19024 7293
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 22284 7488 22336 7540
rect 24308 7488 24360 7540
rect 27620 7488 27672 7540
rect 28908 7488 28960 7540
rect 30104 7488 30156 7540
rect 22468 7420 22520 7472
rect 24768 7420 24820 7472
rect 26884 7420 26936 7472
rect 28264 7420 28316 7472
rect 30932 7488 30984 7540
rect 31024 7488 31076 7540
rect 31760 7463 31812 7472
rect 31760 7429 31769 7463
rect 31769 7429 31803 7463
rect 31803 7429 31812 7463
rect 31760 7420 31812 7429
rect 32220 7531 32272 7540
rect 32220 7497 32229 7531
rect 32229 7497 32263 7531
rect 32263 7497 32272 7531
rect 32220 7488 32272 7497
rect 32404 7420 32456 7472
rect 32680 7420 32732 7472
rect 32864 7420 32916 7472
rect 14832 7216 14884 7268
rect 16120 7216 16172 7268
rect 16488 7216 16540 7268
rect 16764 7259 16816 7268
rect 16764 7225 16773 7259
rect 16773 7225 16807 7259
rect 16807 7225 16816 7259
rect 16764 7216 16816 7225
rect 17684 7216 17736 7268
rect 21180 7284 21232 7336
rect 22376 7352 22428 7404
rect 23480 7352 23532 7404
rect 23572 7284 23624 7336
rect 23756 7327 23808 7336
rect 23756 7293 23765 7327
rect 23765 7293 23799 7327
rect 23799 7293 23808 7327
rect 23756 7284 23808 7293
rect 26424 7352 26476 7404
rect 27160 7395 27212 7404
rect 27160 7361 27169 7395
rect 27169 7361 27203 7395
rect 27203 7361 27212 7395
rect 27160 7352 27212 7361
rect 9680 7148 9732 7200
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 15936 7148 15988 7200
rect 18604 7148 18656 7200
rect 20996 7216 21048 7268
rect 21548 7216 21600 7268
rect 25964 7284 26016 7336
rect 26516 7284 26568 7336
rect 20812 7148 20864 7200
rect 27896 7352 27948 7404
rect 29644 7352 29696 7404
rect 31668 7352 31720 7404
rect 31944 7395 31996 7404
rect 31944 7361 31953 7395
rect 31953 7361 31987 7395
rect 31987 7361 31996 7395
rect 31944 7352 31996 7361
rect 32220 7352 32272 7404
rect 28356 7284 28408 7336
rect 28816 7284 28868 7336
rect 30472 7284 30524 7336
rect 31024 7284 31076 7336
rect 31576 7284 31628 7336
rect 32588 7352 32640 7404
rect 34612 7488 34664 7540
rect 34980 7488 35032 7540
rect 35256 7488 35308 7540
rect 35532 7488 35584 7540
rect 35900 7531 35952 7540
rect 35900 7497 35909 7531
rect 35909 7497 35943 7531
rect 35943 7497 35952 7531
rect 35900 7488 35952 7497
rect 36452 7488 36504 7540
rect 34428 7420 34480 7472
rect 33140 7352 33192 7404
rect 33876 7352 33928 7404
rect 34796 7395 34848 7404
rect 34796 7361 34805 7395
rect 34805 7361 34839 7395
rect 34839 7361 34848 7395
rect 34796 7352 34848 7361
rect 35348 7352 35400 7404
rect 35716 7352 35768 7404
rect 38016 7420 38068 7472
rect 40040 7488 40092 7540
rect 37280 7395 37332 7404
rect 37280 7361 37289 7395
rect 37289 7361 37323 7395
rect 37323 7361 37332 7395
rect 37280 7352 37332 7361
rect 38292 7395 38344 7404
rect 38292 7361 38301 7395
rect 38301 7361 38335 7395
rect 38335 7361 38344 7395
rect 38292 7352 38344 7361
rect 41236 7420 41288 7472
rect 29000 7216 29052 7268
rect 32772 7327 32824 7336
rect 32772 7293 32781 7327
rect 32781 7293 32815 7327
rect 32815 7293 32824 7327
rect 32772 7284 32824 7293
rect 34980 7284 35032 7336
rect 23388 7148 23440 7200
rect 23572 7148 23624 7200
rect 26056 7148 26108 7200
rect 30656 7148 30708 7200
rect 33048 7216 33100 7268
rect 37096 7216 37148 7268
rect 41604 7284 41656 7336
rect 38108 7216 38160 7268
rect 32404 7148 32456 7200
rect 35072 7191 35124 7200
rect 35072 7157 35081 7191
rect 35081 7157 35115 7191
rect 35115 7157 35124 7191
rect 35072 7148 35124 7157
rect 35440 7148 35492 7200
rect 36544 7148 36596 7200
rect 37924 7148 37976 7200
rect 38936 7191 38988 7200
rect 38936 7157 38945 7191
rect 38945 7157 38979 7191
rect 38979 7157 38988 7191
rect 38936 7148 38988 7157
rect 40592 7191 40644 7200
rect 40592 7157 40601 7191
rect 40601 7157 40635 7191
rect 40635 7157 40644 7191
rect 40592 7148 40644 7157
rect 42156 7148 42208 7200
rect 5134 7046 5186 7098
rect 5198 7046 5250 7098
rect 5262 7046 5314 7098
rect 5326 7046 5378 7098
rect 5390 7046 5442 7098
rect 35854 7046 35906 7098
rect 35918 7046 35970 7098
rect 35982 7046 36034 7098
rect 36046 7046 36098 7098
rect 36110 7046 36162 7098
rect 66574 7046 66626 7098
rect 66638 7046 66690 7098
rect 66702 7046 66754 7098
rect 66766 7046 66818 7098
rect 66830 7046 66882 7098
rect 10048 6944 10100 6996
rect 13544 6944 13596 6996
rect 17868 6944 17920 6996
rect 18972 6987 19024 6996
rect 18972 6953 18981 6987
rect 18981 6953 19015 6987
rect 19015 6953 19024 6987
rect 18972 6944 19024 6953
rect 20904 6944 20956 6996
rect 22928 6944 22980 6996
rect 23756 6944 23808 6996
rect 24032 6944 24084 6996
rect 26056 6944 26108 6996
rect 26608 6944 26660 6996
rect 29000 6944 29052 6996
rect 35072 6944 35124 6996
rect 37924 6944 37976 6996
rect 13636 6876 13688 6928
rect 6368 6808 6420 6860
rect 14740 6808 14792 6860
rect 14832 6851 14884 6860
rect 14832 6817 14841 6851
rect 14841 6817 14875 6851
rect 14875 6817 14884 6851
rect 14832 6808 14884 6817
rect 15844 6876 15896 6928
rect 19064 6876 19116 6928
rect 6644 6740 6696 6792
rect 8668 6672 8720 6724
rect 14648 6740 14700 6792
rect 15292 6808 15344 6860
rect 19432 6808 19484 6860
rect 15476 6740 15528 6792
rect 15752 6740 15804 6792
rect 11520 6672 11572 6724
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 18144 6740 18196 6792
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 20444 6808 20496 6860
rect 22376 6808 22428 6860
rect 23388 6876 23440 6928
rect 25412 6876 25464 6928
rect 25964 6876 26016 6928
rect 22560 6740 22612 6792
rect 21364 6672 21416 6724
rect 23940 6808 23992 6860
rect 24860 6808 24912 6860
rect 25504 6783 25556 6792
rect 25504 6749 25513 6783
rect 25513 6749 25547 6783
rect 25547 6749 25556 6783
rect 25504 6740 25556 6749
rect 25688 6783 25740 6792
rect 25688 6749 25697 6783
rect 25697 6749 25731 6783
rect 25731 6749 25740 6783
rect 25688 6740 25740 6749
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 30288 6919 30340 6928
rect 30288 6885 30297 6919
rect 30297 6885 30331 6919
rect 30331 6885 30340 6919
rect 30288 6876 30340 6885
rect 30380 6876 30432 6928
rect 31668 6876 31720 6928
rect 33876 6876 33928 6928
rect 34612 6876 34664 6928
rect 35164 6876 35216 6928
rect 35716 6876 35768 6928
rect 28540 6808 28592 6860
rect 29092 6808 29144 6860
rect 29552 6851 29604 6860
rect 29552 6817 29561 6851
rect 29561 6817 29595 6851
rect 29595 6817 29604 6851
rect 29552 6808 29604 6817
rect 31760 6808 31812 6860
rect 32036 6808 32088 6860
rect 32496 6808 32548 6860
rect 33140 6808 33192 6860
rect 36360 6808 36412 6860
rect 36544 6851 36596 6860
rect 36544 6817 36553 6851
rect 36553 6817 36587 6851
rect 36587 6817 36596 6851
rect 36544 6808 36596 6817
rect 37372 6808 37424 6860
rect 37832 6808 37884 6860
rect 39580 6808 39632 6860
rect 39672 6808 39724 6860
rect 22652 6715 22704 6724
rect 22652 6681 22661 6715
rect 22661 6681 22695 6715
rect 22695 6681 22704 6715
rect 22652 6672 22704 6681
rect 24768 6672 24820 6724
rect 10324 6604 10376 6656
rect 11796 6647 11848 6656
rect 11796 6613 11805 6647
rect 11805 6613 11839 6647
rect 11839 6613 11848 6647
rect 11796 6604 11848 6613
rect 12440 6604 12492 6656
rect 13452 6647 13504 6656
rect 13452 6613 13461 6647
rect 13461 6613 13495 6647
rect 13495 6613 13504 6647
rect 13452 6604 13504 6613
rect 14188 6647 14240 6656
rect 14188 6613 14197 6647
rect 14197 6613 14231 6647
rect 14231 6613 14240 6647
rect 14188 6604 14240 6613
rect 14648 6604 14700 6656
rect 15384 6604 15436 6656
rect 18052 6604 18104 6656
rect 21548 6604 21600 6656
rect 22008 6604 22060 6656
rect 22284 6647 22336 6656
rect 22284 6613 22293 6647
rect 22293 6613 22327 6647
rect 22327 6613 22336 6647
rect 22284 6604 22336 6613
rect 22560 6604 22612 6656
rect 26608 6604 26660 6656
rect 30932 6672 30984 6724
rect 29368 6604 29420 6656
rect 29552 6604 29604 6656
rect 30380 6604 30432 6656
rect 30656 6647 30708 6656
rect 30656 6613 30665 6647
rect 30665 6613 30699 6647
rect 30699 6613 30708 6647
rect 30656 6604 30708 6613
rect 31300 6604 31352 6656
rect 32588 6783 32640 6792
rect 32588 6749 32597 6783
rect 32597 6749 32631 6783
rect 32631 6749 32640 6783
rect 32588 6740 32640 6749
rect 33324 6783 33376 6792
rect 33324 6749 33333 6783
rect 33333 6749 33367 6783
rect 33367 6749 33376 6783
rect 33324 6740 33376 6749
rect 34244 6740 34296 6792
rect 34888 6740 34940 6792
rect 35256 6740 35308 6792
rect 35348 6783 35400 6792
rect 35348 6749 35357 6783
rect 35357 6749 35391 6783
rect 35391 6749 35400 6783
rect 35348 6740 35400 6749
rect 35624 6740 35676 6792
rect 32036 6672 32088 6724
rect 35532 6672 35584 6724
rect 33232 6604 33284 6656
rect 34796 6647 34848 6656
rect 34796 6613 34805 6647
rect 34805 6613 34839 6647
rect 34839 6613 34848 6647
rect 34796 6604 34848 6613
rect 35072 6604 35124 6656
rect 39028 6740 39080 6792
rect 40224 6740 40276 6792
rect 39488 6715 39540 6724
rect 39488 6681 39497 6715
rect 39497 6681 39531 6715
rect 39531 6681 39540 6715
rect 39488 6672 39540 6681
rect 40408 6672 40460 6724
rect 39028 6604 39080 6656
rect 39304 6604 39356 6656
rect 41420 6647 41472 6656
rect 41420 6613 41429 6647
rect 41429 6613 41463 6647
rect 41463 6613 41472 6647
rect 41420 6604 41472 6613
rect 41512 6647 41564 6656
rect 41512 6613 41521 6647
rect 41521 6613 41555 6647
rect 41555 6613 41564 6647
rect 41512 6604 41564 6613
rect 46848 6604 46900 6656
rect 5794 6502 5846 6554
rect 5858 6502 5910 6554
rect 5922 6502 5974 6554
rect 5986 6502 6038 6554
rect 6050 6502 6102 6554
rect 36514 6502 36566 6554
rect 36578 6502 36630 6554
rect 36642 6502 36694 6554
rect 36706 6502 36758 6554
rect 36770 6502 36822 6554
rect 67234 6502 67286 6554
rect 67298 6502 67350 6554
rect 67362 6502 67414 6554
rect 67426 6502 67478 6554
rect 67490 6502 67542 6554
rect 8760 6332 8812 6384
rect 11060 6400 11112 6452
rect 13452 6400 13504 6452
rect 16396 6400 16448 6452
rect 17684 6400 17736 6452
rect 18512 6400 18564 6452
rect 18788 6400 18840 6452
rect 19156 6400 19208 6452
rect 21364 6400 21416 6452
rect 22008 6400 22060 6452
rect 10968 6332 11020 6384
rect 11428 6332 11480 6384
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 8576 6196 8628 6248
rect 5632 6128 5684 6180
rect 11152 6196 11204 6248
rect 12072 6264 12124 6316
rect 14096 6332 14148 6384
rect 15660 6332 15712 6384
rect 17592 6332 17644 6384
rect 17868 6332 17920 6384
rect 19248 6332 19300 6384
rect 11796 6196 11848 6248
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 14740 6264 14792 6316
rect 15476 6264 15528 6316
rect 16212 6264 16264 6316
rect 16672 6307 16724 6316
rect 16672 6273 16681 6307
rect 16681 6273 16715 6307
rect 16715 6273 16724 6307
rect 16672 6264 16724 6273
rect 19616 6264 19668 6316
rect 20076 6264 20128 6316
rect 21088 6332 21140 6384
rect 21364 6264 21416 6316
rect 22376 6375 22428 6384
rect 23296 6400 23348 6452
rect 24032 6400 24084 6452
rect 24400 6443 24452 6452
rect 24400 6409 24409 6443
rect 24409 6409 24443 6443
rect 24443 6409 24452 6443
rect 24400 6400 24452 6409
rect 26700 6400 26752 6452
rect 27712 6400 27764 6452
rect 22376 6341 22401 6375
rect 22401 6341 22428 6375
rect 22376 6332 22428 6341
rect 26792 6332 26844 6384
rect 27528 6332 27580 6384
rect 27620 6332 27672 6384
rect 29460 6332 29512 6384
rect 29736 6332 29788 6384
rect 23296 6307 23348 6316
rect 23296 6273 23305 6307
rect 23305 6273 23339 6307
rect 23339 6273 23348 6307
rect 23296 6264 23348 6273
rect 23388 6264 23440 6316
rect 13268 6196 13320 6248
rect 13912 6196 13964 6248
rect 14372 6239 14424 6248
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 15568 6196 15620 6248
rect 17408 6196 17460 6248
rect 17868 6196 17920 6248
rect 19432 6196 19484 6248
rect 19892 6239 19944 6248
rect 19892 6205 19901 6239
rect 19901 6205 19935 6239
rect 19935 6205 19944 6239
rect 19892 6196 19944 6205
rect 19984 6196 20036 6248
rect 21640 6196 21692 6248
rect 6920 6060 6972 6112
rect 9588 6060 9640 6112
rect 13636 6060 13688 6112
rect 14096 6060 14148 6112
rect 16028 6103 16080 6112
rect 16028 6069 16037 6103
rect 16037 6069 16071 6103
rect 16071 6069 16080 6103
rect 16028 6060 16080 6069
rect 16580 6060 16632 6112
rect 19156 6171 19208 6180
rect 19156 6137 19165 6171
rect 19165 6137 19199 6171
rect 19199 6137 19208 6171
rect 19156 6128 19208 6137
rect 20352 6128 20404 6180
rect 21732 6128 21784 6180
rect 22744 6196 22796 6248
rect 23756 6264 23808 6316
rect 23848 6307 23900 6316
rect 23848 6273 23857 6307
rect 23857 6273 23891 6307
rect 23891 6273 23900 6307
rect 23848 6264 23900 6273
rect 25044 6264 25096 6316
rect 19248 6060 19300 6112
rect 21824 6060 21876 6112
rect 22192 6060 22244 6112
rect 23940 6196 23992 6248
rect 25320 6239 25372 6248
rect 25320 6205 25329 6239
rect 25329 6205 25363 6239
rect 25363 6205 25372 6239
rect 25320 6196 25372 6205
rect 26148 6264 26200 6316
rect 29000 6264 29052 6316
rect 30104 6400 30156 6452
rect 30380 6400 30432 6452
rect 31300 6400 31352 6452
rect 30288 6332 30340 6384
rect 26792 6196 26844 6248
rect 28908 6196 28960 6248
rect 29644 6239 29696 6248
rect 29644 6205 29653 6239
rect 29653 6205 29687 6239
rect 29687 6205 29696 6239
rect 29644 6196 29696 6205
rect 29920 6239 29972 6248
rect 29920 6205 29929 6239
rect 29929 6205 29963 6239
rect 29963 6205 29972 6239
rect 29920 6196 29972 6205
rect 29552 6128 29604 6180
rect 25044 6060 25096 6112
rect 25136 6103 25188 6112
rect 25136 6069 25145 6103
rect 25145 6069 25179 6103
rect 25179 6069 25188 6103
rect 25136 6060 25188 6069
rect 28540 6060 28592 6112
rect 29736 6060 29788 6112
rect 30932 6307 30984 6316
rect 30932 6273 30941 6307
rect 30941 6273 30975 6307
rect 30975 6273 30984 6307
rect 30932 6264 30984 6273
rect 31760 6332 31812 6384
rect 38844 6400 38896 6452
rect 34888 6332 34940 6384
rect 40224 6375 40276 6384
rect 40224 6341 40233 6375
rect 40233 6341 40267 6375
rect 40267 6341 40276 6375
rect 40224 6332 40276 6341
rect 35164 6307 35216 6316
rect 35164 6273 35173 6307
rect 35173 6273 35207 6307
rect 35207 6273 35216 6307
rect 35164 6264 35216 6273
rect 35256 6307 35308 6316
rect 35256 6273 35265 6307
rect 35265 6273 35299 6307
rect 35299 6273 35308 6307
rect 35256 6264 35308 6273
rect 30380 6103 30432 6112
rect 30380 6069 30389 6103
rect 30389 6069 30423 6103
rect 30423 6069 30432 6103
rect 30380 6060 30432 6069
rect 31760 6239 31812 6248
rect 31760 6205 31769 6239
rect 31769 6205 31803 6239
rect 31803 6205 31812 6239
rect 31760 6196 31812 6205
rect 32128 6196 32180 6248
rect 32956 6196 33008 6248
rect 33416 6196 33468 6248
rect 34888 6196 34940 6248
rect 35716 6264 35768 6316
rect 37004 6264 37056 6316
rect 39580 6264 39632 6316
rect 41420 6264 41472 6316
rect 42708 6307 42760 6316
rect 42708 6273 42717 6307
rect 42717 6273 42751 6307
rect 42751 6273 42760 6307
rect 42708 6264 42760 6273
rect 42800 6307 42852 6316
rect 42800 6273 42809 6307
rect 42809 6273 42843 6307
rect 42843 6273 42852 6307
rect 42800 6264 42852 6273
rect 43352 6332 43404 6384
rect 43260 6264 43312 6316
rect 35624 6196 35676 6248
rect 32588 6128 32640 6180
rect 34336 6128 34388 6180
rect 33140 6060 33192 6112
rect 35256 6060 35308 6112
rect 35624 6060 35676 6112
rect 36452 6060 36504 6112
rect 36912 6060 36964 6112
rect 37924 6196 37976 6248
rect 38936 6196 38988 6248
rect 39488 6060 39540 6112
rect 41144 6103 41196 6112
rect 41144 6069 41153 6103
rect 41153 6069 41187 6103
rect 41187 6069 41196 6103
rect 41144 6060 41196 6069
rect 41972 6103 42024 6112
rect 41972 6069 41981 6103
rect 41981 6069 42015 6103
rect 42015 6069 42024 6103
rect 41972 6060 42024 6069
rect 42616 6060 42668 6112
rect 45468 6128 45520 6180
rect 48872 6060 48924 6112
rect 5134 5958 5186 6010
rect 5198 5958 5250 6010
rect 5262 5958 5314 6010
rect 5326 5958 5378 6010
rect 5390 5958 5442 6010
rect 35854 5958 35906 6010
rect 35918 5958 35970 6010
rect 35982 5958 36034 6010
rect 36046 5958 36098 6010
rect 36110 5958 36162 6010
rect 66574 5958 66626 6010
rect 66638 5958 66690 6010
rect 66702 5958 66754 6010
rect 66766 5958 66818 6010
rect 66830 5958 66882 6010
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 5724 5788 5776 5840
rect 11060 5788 11112 5840
rect 7748 5720 7800 5772
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 9036 5695 9088 5704
rect 9036 5661 9045 5695
rect 9045 5661 9079 5695
rect 9079 5661 9088 5695
rect 9036 5652 9088 5661
rect 9588 5652 9640 5704
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 10600 5763 10652 5772
rect 10600 5729 10609 5763
rect 10609 5729 10643 5763
rect 10643 5729 10652 5763
rect 10600 5720 10652 5729
rect 17500 5856 17552 5908
rect 11888 5763 11940 5772
rect 11888 5729 11897 5763
rect 11897 5729 11931 5763
rect 11931 5729 11940 5763
rect 11888 5720 11940 5729
rect 11980 5695 12032 5704
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 8576 5584 8628 5636
rect 10232 5584 10284 5636
rect 14556 5720 14608 5772
rect 14832 5720 14884 5772
rect 19524 5788 19576 5840
rect 20168 5899 20220 5908
rect 20168 5865 20177 5899
rect 20177 5865 20211 5899
rect 20211 5865 20220 5899
rect 20168 5856 20220 5865
rect 20260 5856 20312 5908
rect 20812 5856 20864 5908
rect 21456 5899 21508 5908
rect 21456 5865 21465 5899
rect 21465 5865 21499 5899
rect 21499 5865 21508 5899
rect 21456 5856 21508 5865
rect 22008 5856 22060 5908
rect 23940 5856 23992 5908
rect 24308 5856 24360 5908
rect 20536 5788 20588 5840
rect 22284 5788 22336 5840
rect 23756 5788 23808 5840
rect 13452 5627 13504 5636
rect 13452 5593 13461 5627
rect 13461 5593 13495 5627
rect 13495 5593 13504 5627
rect 13452 5584 13504 5593
rect 14648 5652 14700 5704
rect 15108 5695 15160 5704
rect 15108 5661 15117 5695
rect 15117 5661 15151 5695
rect 15151 5661 15160 5695
rect 15108 5652 15160 5661
rect 15292 5652 15344 5704
rect 14924 5584 14976 5636
rect 16304 5652 16356 5704
rect 17684 5695 17736 5704
rect 17684 5661 17693 5695
rect 17693 5661 17727 5695
rect 17727 5661 17736 5695
rect 17684 5652 17736 5661
rect 17868 5695 17920 5704
rect 17868 5661 17877 5695
rect 17877 5661 17911 5695
rect 17911 5661 17920 5695
rect 17868 5652 17920 5661
rect 18880 5720 18932 5772
rect 22560 5720 22612 5772
rect 23388 5720 23440 5772
rect 24308 5720 24360 5772
rect 24676 5788 24728 5840
rect 20168 5652 20220 5704
rect 21180 5652 21232 5704
rect 22192 5695 22244 5704
rect 22192 5661 22201 5695
rect 22201 5661 22235 5695
rect 22235 5661 22244 5695
rect 22192 5652 22244 5661
rect 3884 5516 3936 5568
rect 6736 5516 6788 5568
rect 9956 5559 10008 5568
rect 9956 5525 9965 5559
rect 9965 5525 9999 5559
rect 9999 5525 10008 5559
rect 9956 5516 10008 5525
rect 16672 5584 16724 5636
rect 24216 5652 24268 5704
rect 26332 5856 26384 5908
rect 27068 5856 27120 5908
rect 27436 5856 27488 5908
rect 25136 5788 25188 5840
rect 25320 5763 25372 5772
rect 25320 5729 25329 5763
rect 25329 5729 25363 5763
rect 25363 5729 25372 5763
rect 25320 5720 25372 5729
rect 25504 5763 25556 5772
rect 25504 5729 25513 5763
rect 25513 5729 25547 5763
rect 25547 5729 25556 5763
rect 25504 5720 25556 5729
rect 25872 5720 25924 5772
rect 25044 5584 25096 5636
rect 25688 5695 25740 5704
rect 25688 5661 25697 5695
rect 25697 5661 25731 5695
rect 25731 5661 25740 5695
rect 25688 5652 25740 5661
rect 27344 5763 27396 5772
rect 27344 5729 27353 5763
rect 27353 5729 27387 5763
rect 27387 5729 27396 5763
rect 27344 5720 27396 5729
rect 29460 5720 29512 5772
rect 29552 5763 29604 5772
rect 29552 5729 29561 5763
rect 29561 5729 29595 5763
rect 29595 5729 29604 5763
rect 29552 5720 29604 5729
rect 29920 5720 29972 5772
rect 26148 5652 26200 5704
rect 25872 5584 25924 5636
rect 28908 5652 28960 5704
rect 30472 5899 30524 5908
rect 30472 5865 30481 5899
rect 30481 5865 30515 5899
rect 30515 5865 30524 5899
rect 30472 5856 30524 5865
rect 31944 5856 31996 5908
rect 32956 5856 33008 5908
rect 33784 5856 33836 5908
rect 35348 5856 35400 5908
rect 36820 5856 36872 5908
rect 37280 5856 37332 5908
rect 38660 5856 38712 5908
rect 30932 5763 30984 5772
rect 30932 5729 30941 5763
rect 30941 5729 30975 5763
rect 30975 5729 30984 5763
rect 30932 5720 30984 5729
rect 29092 5584 29144 5636
rect 16396 5559 16448 5568
rect 16396 5525 16405 5559
rect 16405 5525 16439 5559
rect 16439 5525 16448 5559
rect 16396 5516 16448 5525
rect 17132 5559 17184 5568
rect 17132 5525 17141 5559
rect 17141 5525 17175 5559
rect 17175 5525 17184 5559
rect 17132 5516 17184 5525
rect 18604 5559 18656 5568
rect 18604 5525 18613 5559
rect 18613 5525 18647 5559
rect 18647 5525 18656 5559
rect 18604 5516 18656 5525
rect 18972 5516 19024 5568
rect 19156 5516 19208 5568
rect 19892 5516 19944 5568
rect 20076 5516 20128 5568
rect 20812 5516 20864 5568
rect 21640 5516 21692 5568
rect 22192 5516 22244 5568
rect 24952 5516 25004 5568
rect 25596 5516 25648 5568
rect 26700 5559 26752 5568
rect 26700 5525 26709 5559
rect 26709 5525 26743 5559
rect 26743 5525 26752 5559
rect 26700 5516 26752 5525
rect 27436 5559 27488 5568
rect 27436 5525 27445 5559
rect 27445 5525 27479 5559
rect 27479 5525 27488 5559
rect 27436 5516 27488 5525
rect 28080 5516 28132 5568
rect 32036 5720 32088 5772
rect 31576 5652 31628 5704
rect 32220 5652 32272 5704
rect 32588 5695 32640 5704
rect 32588 5661 32597 5695
rect 32597 5661 32631 5695
rect 32631 5661 32640 5695
rect 32588 5652 32640 5661
rect 34428 5831 34480 5840
rect 34428 5797 34437 5831
rect 34437 5797 34471 5831
rect 34471 5797 34480 5831
rect 34428 5788 34480 5797
rect 34980 5788 35032 5840
rect 36452 5788 36504 5840
rect 33416 5652 33468 5704
rect 31668 5627 31720 5636
rect 31668 5593 31677 5627
rect 31677 5593 31711 5627
rect 31711 5593 31720 5627
rect 31668 5584 31720 5593
rect 32496 5584 32548 5636
rect 32864 5584 32916 5636
rect 34244 5652 34296 5704
rect 34520 5695 34572 5704
rect 34520 5661 34529 5695
rect 34529 5661 34563 5695
rect 34563 5661 34572 5695
rect 34520 5652 34572 5661
rect 35072 5695 35124 5704
rect 35072 5661 35081 5695
rect 35081 5661 35115 5695
rect 35115 5661 35124 5695
rect 35072 5652 35124 5661
rect 35900 5720 35952 5772
rect 35256 5695 35308 5704
rect 35256 5661 35265 5695
rect 35265 5661 35299 5695
rect 35299 5661 35308 5695
rect 35256 5652 35308 5661
rect 35440 5695 35492 5704
rect 35440 5661 35449 5695
rect 35449 5661 35483 5695
rect 35483 5661 35492 5695
rect 35440 5652 35492 5661
rect 36268 5652 36320 5704
rect 36912 5763 36964 5772
rect 36912 5729 36921 5763
rect 36921 5729 36955 5763
rect 36955 5729 36964 5763
rect 36912 5720 36964 5729
rect 38844 5788 38896 5840
rect 39672 5788 39724 5840
rect 39304 5763 39356 5772
rect 39304 5729 39313 5763
rect 39313 5729 39347 5763
rect 39347 5729 39356 5763
rect 39304 5720 39356 5729
rect 42800 5788 42852 5840
rect 41144 5720 41196 5772
rect 42984 5720 43036 5772
rect 45192 5720 45244 5772
rect 42892 5695 42944 5704
rect 42892 5661 42901 5695
rect 42901 5661 42935 5695
rect 42935 5661 42944 5695
rect 42892 5652 42944 5661
rect 34612 5584 34664 5636
rect 35808 5584 35860 5636
rect 36452 5584 36504 5636
rect 37280 5584 37332 5636
rect 44364 5695 44416 5704
rect 44364 5661 44373 5695
rect 44373 5661 44407 5695
rect 44407 5661 44416 5695
rect 44364 5652 44416 5661
rect 45836 5652 45888 5704
rect 45652 5584 45704 5636
rect 36176 5516 36228 5568
rect 37832 5516 37884 5568
rect 37924 5516 37976 5568
rect 38936 5516 38988 5568
rect 39948 5559 40000 5568
rect 39948 5525 39957 5559
rect 39957 5525 39991 5559
rect 39991 5525 40000 5559
rect 39948 5516 40000 5525
rect 40776 5559 40828 5568
rect 40776 5525 40785 5559
rect 40785 5525 40819 5559
rect 40819 5525 40828 5559
rect 40776 5516 40828 5525
rect 43720 5559 43772 5568
rect 43720 5525 43729 5559
rect 43729 5525 43763 5559
rect 43763 5525 43772 5559
rect 43720 5516 43772 5525
rect 47032 5516 47084 5568
rect 5794 5414 5846 5466
rect 5858 5414 5910 5466
rect 5922 5414 5974 5466
rect 5986 5414 6038 5466
rect 6050 5414 6102 5466
rect 36514 5414 36566 5466
rect 36578 5414 36630 5466
rect 36642 5414 36694 5466
rect 36706 5414 36758 5466
rect 36770 5414 36822 5466
rect 67234 5414 67286 5466
rect 67298 5414 67350 5466
rect 67362 5414 67414 5466
rect 67426 5414 67478 5466
rect 67490 5414 67542 5466
rect 9036 5312 9088 5364
rect 9128 5355 9180 5364
rect 9128 5321 9137 5355
rect 9137 5321 9171 5355
rect 9171 5321 9180 5355
rect 9128 5312 9180 5321
rect 11520 5355 11572 5364
rect 11520 5321 11529 5355
rect 11529 5321 11563 5355
rect 11563 5321 11572 5355
rect 11520 5312 11572 5321
rect 12256 5355 12308 5364
rect 12256 5321 12265 5355
rect 12265 5321 12299 5355
rect 12299 5321 12308 5355
rect 12256 5312 12308 5321
rect 13360 5312 13412 5364
rect 15568 5312 15620 5364
rect 16212 5312 16264 5364
rect 16948 5312 17000 5364
rect 17224 5312 17276 5364
rect 17684 5312 17736 5364
rect 17960 5312 18012 5364
rect 18236 5312 18288 5364
rect 7104 5244 7156 5296
rect 16488 5244 16540 5296
rect 16672 5287 16724 5296
rect 16672 5253 16681 5287
rect 16681 5253 16715 5287
rect 16715 5253 16724 5287
rect 16672 5244 16724 5253
rect 18328 5244 18380 5296
rect 18512 5244 18564 5296
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 8668 5176 8720 5228
rect 10048 5176 10100 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 12440 5219 12492 5228
rect 12440 5185 12449 5219
rect 12449 5185 12483 5219
rect 12483 5185 12492 5219
rect 12440 5176 12492 5185
rect 16028 5176 16080 5228
rect 20260 5312 20312 5364
rect 20720 5312 20772 5364
rect 21364 5312 21416 5364
rect 21916 5312 21968 5364
rect 23020 5312 23072 5364
rect 23480 5312 23532 5364
rect 24216 5312 24268 5364
rect 25504 5355 25556 5364
rect 25504 5321 25513 5355
rect 25513 5321 25547 5355
rect 25547 5321 25556 5355
rect 25504 5312 25556 5321
rect 26148 5312 26200 5364
rect 26424 5312 26476 5364
rect 29736 5312 29788 5364
rect 30288 5355 30340 5364
rect 30288 5321 30297 5355
rect 30297 5321 30331 5355
rect 30331 5321 30340 5355
rect 30288 5312 30340 5321
rect 33324 5312 33376 5364
rect 33600 5355 33652 5364
rect 33600 5321 33609 5355
rect 33609 5321 33643 5355
rect 33643 5321 33652 5355
rect 33600 5312 33652 5321
rect 35164 5355 35216 5364
rect 35164 5321 35173 5355
rect 35173 5321 35207 5355
rect 35207 5321 35216 5355
rect 35164 5312 35216 5321
rect 36176 5312 36228 5364
rect 36452 5312 36504 5364
rect 37004 5312 37056 5364
rect 19248 5287 19300 5296
rect 19248 5253 19257 5287
rect 19257 5253 19291 5287
rect 19291 5253 19300 5287
rect 19248 5244 19300 5253
rect 20536 5244 20588 5296
rect 20812 5176 20864 5228
rect 21088 5176 21140 5228
rect 9680 5108 9732 5160
rect 9864 5108 9916 5160
rect 8392 5040 8444 5092
rect 14004 5108 14056 5160
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 14648 5108 14700 5117
rect 16212 5108 16264 5160
rect 16488 5108 16540 5160
rect 16764 5151 16816 5160
rect 16764 5117 16773 5151
rect 16773 5117 16807 5151
rect 16807 5117 16816 5151
rect 16764 5108 16816 5117
rect 17776 5151 17828 5160
rect 17776 5117 17785 5151
rect 17785 5117 17819 5151
rect 17819 5117 17828 5151
rect 17776 5108 17828 5117
rect 17868 5151 17920 5160
rect 17868 5117 17877 5151
rect 17877 5117 17911 5151
rect 17911 5117 17920 5151
rect 17868 5108 17920 5117
rect 18236 5108 18288 5160
rect 18512 5108 18564 5160
rect 18604 5108 18656 5160
rect 21548 5176 21600 5228
rect 21640 5219 21692 5228
rect 21640 5185 21649 5219
rect 21649 5185 21683 5219
rect 21683 5185 21692 5219
rect 21640 5176 21692 5185
rect 22744 5287 22796 5296
rect 22744 5253 22753 5287
rect 22753 5253 22787 5287
rect 22787 5253 22796 5287
rect 22744 5244 22796 5253
rect 23848 5176 23900 5228
rect 24860 5176 24912 5228
rect 25872 5176 25924 5228
rect 21364 5151 21416 5160
rect 21364 5117 21373 5151
rect 21373 5117 21407 5151
rect 21407 5117 21416 5151
rect 21364 5108 21416 5117
rect 11060 5040 11112 5092
rect 12716 5040 12768 5092
rect 12808 5040 12860 5092
rect 16672 5040 16724 5092
rect 8300 4972 8352 5024
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 10876 4972 10928 5024
rect 13452 4972 13504 5024
rect 14280 5015 14332 5024
rect 14280 4981 14289 5015
rect 14289 4981 14323 5015
rect 14323 4981 14332 5015
rect 14280 4972 14332 4981
rect 16212 5015 16264 5024
rect 16212 4981 16221 5015
rect 16221 4981 16255 5015
rect 16255 4981 16264 5015
rect 16212 4972 16264 4981
rect 17776 4972 17828 5024
rect 18052 4972 18104 5024
rect 18328 4972 18380 5024
rect 18696 4972 18748 5024
rect 18880 5015 18932 5024
rect 18880 4981 18889 5015
rect 18889 4981 18923 5015
rect 18923 4981 18932 5015
rect 18880 4972 18932 4981
rect 23388 5040 23440 5092
rect 23572 5040 23624 5092
rect 24400 5040 24452 5092
rect 23112 4972 23164 5024
rect 27344 5108 27396 5160
rect 27896 5219 27948 5228
rect 27896 5185 27905 5219
rect 27905 5185 27939 5219
rect 27939 5185 27948 5219
rect 27896 5176 27948 5185
rect 29644 5244 29696 5296
rect 28540 5176 28592 5228
rect 31300 5244 31352 5296
rect 32404 5244 32456 5296
rect 32128 5176 32180 5228
rect 33140 5244 33192 5296
rect 34336 5244 34388 5296
rect 35256 5244 35308 5296
rect 36820 5244 36872 5296
rect 38936 5312 38988 5364
rect 42708 5312 42760 5364
rect 37464 5244 37516 5296
rect 27896 5040 27948 5092
rect 28356 5108 28408 5160
rect 28816 5108 28868 5160
rect 29644 5040 29696 5092
rect 32036 5108 32088 5160
rect 33416 5219 33468 5228
rect 33416 5185 33425 5219
rect 33425 5185 33459 5219
rect 33459 5185 33468 5219
rect 33416 5176 33468 5185
rect 34796 5176 34848 5228
rect 35532 5176 35584 5228
rect 35808 5219 35860 5228
rect 35808 5185 35817 5219
rect 35817 5185 35851 5219
rect 35851 5185 35860 5219
rect 35808 5176 35860 5185
rect 33692 5151 33744 5160
rect 33692 5117 33701 5151
rect 33701 5117 33735 5151
rect 33735 5117 33744 5151
rect 33692 5108 33744 5117
rect 34152 5108 34204 5160
rect 36084 5219 36136 5228
rect 36084 5185 36093 5219
rect 36093 5185 36127 5219
rect 36127 5185 36136 5219
rect 36084 5176 36136 5185
rect 36176 5219 36228 5228
rect 36176 5185 36185 5219
rect 36185 5185 36219 5219
rect 36219 5185 36228 5219
rect 36176 5176 36228 5185
rect 36912 5176 36964 5228
rect 26884 4972 26936 5024
rect 26976 5015 27028 5024
rect 26976 4981 26985 5015
rect 26985 4981 27019 5015
rect 27019 4981 27028 5015
rect 26976 4972 27028 4981
rect 27712 5015 27764 5024
rect 27712 4981 27721 5015
rect 27721 4981 27755 5015
rect 27755 4981 27764 5015
rect 27712 4972 27764 4981
rect 28264 4972 28316 5024
rect 30472 4972 30524 5024
rect 32220 5040 32272 5092
rect 36544 5108 36596 5160
rect 37740 5108 37792 5160
rect 38200 5219 38252 5228
rect 38200 5185 38209 5219
rect 38209 5185 38243 5219
rect 38243 5185 38252 5219
rect 38200 5176 38252 5185
rect 32036 4972 32088 5024
rect 32772 4972 32824 5024
rect 33416 4972 33468 5024
rect 37280 4972 37332 5024
rect 37372 5015 37424 5024
rect 37372 4981 37381 5015
rect 37381 4981 37415 5015
rect 37415 4981 37424 5015
rect 37372 4972 37424 4981
rect 39948 5176 40000 5228
rect 40776 5176 40828 5228
rect 41328 5176 41380 5228
rect 44180 5176 44232 5228
rect 46756 5176 46808 5228
rect 47032 5219 47084 5228
rect 47032 5185 47041 5219
rect 47041 5185 47075 5219
rect 47075 5185 47084 5219
rect 47032 5176 47084 5185
rect 41696 5108 41748 5160
rect 42708 5040 42760 5092
rect 45560 5151 45612 5160
rect 45560 5117 45569 5151
rect 45569 5117 45603 5151
rect 45603 5117 45612 5151
rect 45560 5108 45612 5117
rect 46940 5151 46992 5160
rect 46940 5117 46949 5151
rect 46949 5117 46983 5151
rect 46983 5117 46992 5151
rect 46940 5108 46992 5117
rect 76932 5108 76984 5160
rect 44824 5083 44876 5092
rect 44824 5049 44833 5083
rect 44833 5049 44867 5083
rect 44867 5049 44876 5083
rect 44824 5040 44876 5049
rect 47952 5040 48004 5092
rect 42064 4972 42116 5024
rect 43260 4972 43312 5024
rect 43352 5015 43404 5024
rect 43352 4981 43361 5015
rect 43361 4981 43395 5015
rect 43395 4981 43404 5015
rect 43352 4972 43404 4981
rect 45744 4972 45796 5024
rect 47216 4972 47268 5024
rect 49608 4972 49660 5024
rect 76656 4972 76708 5024
rect 5134 4870 5186 4922
rect 5198 4870 5250 4922
rect 5262 4870 5314 4922
rect 5326 4870 5378 4922
rect 5390 4870 5442 4922
rect 35854 4870 35906 4922
rect 35918 4870 35970 4922
rect 35982 4870 36034 4922
rect 36046 4870 36098 4922
rect 36110 4870 36162 4922
rect 66574 4870 66626 4922
rect 66638 4870 66690 4922
rect 66702 4870 66754 4922
rect 66766 4870 66818 4922
rect 66830 4870 66882 4922
rect 9772 4768 9824 4820
rect 11244 4768 11296 4820
rect 15752 4768 15804 4820
rect 16120 4768 16172 4820
rect 19064 4811 19116 4820
rect 19064 4777 19073 4811
rect 19073 4777 19107 4811
rect 19107 4777 19116 4811
rect 19064 4768 19116 4777
rect 19432 4768 19484 4820
rect 21456 4768 21508 4820
rect 23204 4768 23256 4820
rect 24492 4768 24544 4820
rect 27988 4768 28040 4820
rect 29644 4811 29696 4820
rect 29644 4777 29653 4811
rect 29653 4777 29687 4811
rect 29687 4777 29696 4811
rect 29644 4768 29696 4777
rect 30196 4768 30248 4820
rect 30564 4768 30616 4820
rect 31208 4768 31260 4820
rect 32772 4768 32824 4820
rect 32864 4811 32916 4820
rect 32864 4777 32873 4811
rect 32873 4777 32907 4811
rect 32907 4777 32916 4811
rect 32864 4768 32916 4777
rect 33692 4768 33744 4820
rect 36268 4768 36320 4820
rect 37280 4768 37332 4820
rect 11060 4700 11112 4752
rect 12348 4700 12400 4752
rect 12624 4743 12676 4752
rect 12624 4709 12633 4743
rect 12633 4709 12667 4743
rect 12667 4709 12676 4743
rect 12624 4700 12676 4709
rect 16764 4700 16816 4752
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 10600 4607 10652 4616
rect 10600 4573 10609 4607
rect 10609 4573 10643 4607
rect 10643 4573 10652 4607
rect 10600 4564 10652 4573
rect 11336 4607 11388 4616
rect 11336 4573 11345 4607
rect 11345 4573 11379 4607
rect 11379 4573 11388 4607
rect 11336 4564 11388 4573
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 13544 4675 13596 4684
rect 13544 4641 13553 4675
rect 13553 4641 13587 4675
rect 13587 4641 13596 4675
rect 13544 4632 13596 4641
rect 14280 4632 14332 4684
rect 16212 4632 16264 4684
rect 12348 4564 12400 4616
rect 12808 4607 12860 4616
rect 12808 4573 12817 4607
rect 12817 4573 12851 4607
rect 12851 4573 12860 4607
rect 12808 4564 12860 4573
rect 15016 4564 15068 4616
rect 17132 4632 17184 4684
rect 19524 4700 19576 4752
rect 19892 4700 19944 4752
rect 21732 4700 21784 4752
rect 21824 4743 21876 4752
rect 21824 4709 21833 4743
rect 21833 4709 21867 4743
rect 21867 4709 21876 4743
rect 21824 4700 21876 4709
rect 9772 4496 9824 4548
rect 12716 4496 12768 4548
rect 15844 4496 15896 4548
rect 17592 4564 17644 4616
rect 20628 4632 20680 4684
rect 23572 4632 23624 4684
rect 24308 4632 24360 4684
rect 24768 4675 24820 4684
rect 24768 4641 24777 4675
rect 24777 4641 24811 4675
rect 24811 4641 24820 4675
rect 24768 4632 24820 4641
rect 25044 4632 25096 4684
rect 32496 4700 32548 4752
rect 26332 4632 26384 4684
rect 26424 4675 26476 4684
rect 26424 4641 26433 4675
rect 26433 4641 26467 4675
rect 26467 4641 26476 4675
rect 26424 4632 26476 4641
rect 26884 4632 26936 4684
rect 20904 4564 20956 4616
rect 21548 4564 21600 4616
rect 21916 4607 21968 4616
rect 21916 4573 21925 4607
rect 21925 4573 21959 4607
rect 21959 4573 21968 4607
rect 21916 4564 21968 4573
rect 22652 4607 22704 4616
rect 22652 4573 22661 4607
rect 22661 4573 22695 4607
rect 22695 4573 22704 4607
rect 22652 4564 22704 4573
rect 23020 4564 23072 4616
rect 23388 4564 23440 4616
rect 24032 4564 24084 4616
rect 24676 4607 24728 4616
rect 24676 4573 24685 4607
rect 24685 4573 24719 4607
rect 24719 4573 24728 4607
rect 24676 4564 24728 4573
rect 27436 4564 27488 4616
rect 17868 4496 17920 4548
rect 18052 4539 18104 4548
rect 18052 4505 18061 4539
rect 18061 4505 18095 4539
rect 18095 4505 18104 4539
rect 18052 4496 18104 4505
rect 6460 4428 6512 4480
rect 6828 4471 6880 4480
rect 6828 4437 6837 4471
rect 6837 4437 6871 4471
rect 6871 4437 6880 4471
rect 6828 4428 6880 4437
rect 9588 4428 9640 4480
rect 12440 4428 12492 4480
rect 12900 4428 12952 4480
rect 15660 4428 15712 4480
rect 18328 4428 18380 4480
rect 18420 4428 18472 4480
rect 20168 4496 20220 4548
rect 19616 4428 19668 4480
rect 19892 4428 19944 4480
rect 22284 4428 22336 4480
rect 24768 4428 24820 4480
rect 24952 4496 25004 4548
rect 26240 4496 26292 4548
rect 27528 4496 27580 4548
rect 28172 4632 28224 4684
rect 27988 4564 28040 4616
rect 28264 4564 28316 4616
rect 28908 4675 28960 4684
rect 28908 4641 28917 4675
rect 28917 4641 28951 4675
rect 28951 4641 28960 4675
rect 28908 4632 28960 4641
rect 30472 4632 30524 4684
rect 30748 4675 30800 4684
rect 30748 4641 30757 4675
rect 30757 4641 30791 4675
rect 30791 4641 30800 4675
rect 30748 4632 30800 4641
rect 31208 4632 31260 4684
rect 31576 4632 31628 4684
rect 31852 4675 31904 4684
rect 31852 4641 31861 4675
rect 31861 4641 31895 4675
rect 31895 4641 31904 4675
rect 31852 4632 31904 4641
rect 31944 4675 31996 4684
rect 31944 4641 31953 4675
rect 31953 4641 31987 4675
rect 31987 4641 31996 4675
rect 31944 4632 31996 4641
rect 36820 4700 36872 4752
rect 37464 4700 37516 4752
rect 32864 4632 32916 4684
rect 33048 4632 33100 4684
rect 33232 4632 33284 4684
rect 37372 4632 37424 4684
rect 37740 4675 37792 4684
rect 37740 4641 37749 4675
rect 37749 4641 37783 4675
rect 37783 4641 37792 4675
rect 37740 4632 37792 4641
rect 37832 4632 37884 4684
rect 38936 4632 38988 4684
rect 29368 4564 29420 4616
rect 29920 4564 29972 4616
rect 30288 4607 30340 4616
rect 30288 4573 30297 4607
rect 30297 4573 30331 4607
rect 30331 4573 30340 4607
rect 30288 4564 30340 4573
rect 29276 4496 29328 4548
rect 30748 4496 30800 4548
rect 31760 4539 31812 4548
rect 31760 4505 31769 4539
rect 31769 4505 31803 4539
rect 31803 4505 31812 4539
rect 31760 4496 31812 4505
rect 33324 4564 33376 4616
rect 27620 4428 27672 4480
rect 28448 4428 28500 4480
rect 29552 4471 29604 4480
rect 29552 4437 29561 4471
rect 29561 4437 29595 4471
rect 29595 4437 29604 4471
rect 29552 4428 29604 4437
rect 30472 4428 30524 4480
rect 31668 4428 31720 4480
rect 32588 4496 32640 4548
rect 33140 4539 33192 4548
rect 33140 4505 33149 4539
rect 33149 4505 33183 4539
rect 33183 4505 33192 4539
rect 33140 4496 33192 4505
rect 34612 4564 34664 4616
rect 35256 4564 35308 4616
rect 34520 4428 34572 4480
rect 36084 4428 36136 4480
rect 36268 4471 36320 4480
rect 36268 4437 36277 4471
rect 36277 4437 36311 4471
rect 36311 4437 36320 4471
rect 36268 4428 36320 4437
rect 37556 4471 37608 4480
rect 37556 4437 37565 4471
rect 37565 4437 37599 4471
rect 37599 4437 37608 4471
rect 37556 4428 37608 4437
rect 37924 4607 37976 4616
rect 37924 4573 37933 4607
rect 37933 4573 37967 4607
rect 37967 4573 37976 4607
rect 37924 4564 37976 4573
rect 41696 4768 41748 4820
rect 42064 4768 42116 4820
rect 42892 4768 42944 4820
rect 43628 4768 43680 4820
rect 45836 4768 45888 4820
rect 76932 4811 76984 4820
rect 76932 4777 76941 4811
rect 76941 4777 76975 4811
rect 76975 4777 76984 4811
rect 76932 4768 76984 4777
rect 43260 4632 43312 4684
rect 45468 4632 45520 4684
rect 47216 4675 47268 4684
rect 47216 4641 47225 4675
rect 47225 4641 47259 4675
rect 47259 4641 47268 4675
rect 47216 4632 47268 4641
rect 48320 4632 48372 4684
rect 40500 4564 40552 4616
rect 41144 4564 41196 4616
rect 43996 4564 44048 4616
rect 39580 4496 39632 4548
rect 39948 4539 40000 4548
rect 39948 4505 39957 4539
rect 39957 4505 39991 4539
rect 39991 4505 40000 4539
rect 39948 4496 40000 4505
rect 40776 4496 40828 4548
rect 41052 4496 41104 4548
rect 43628 4496 43680 4548
rect 38568 4428 38620 4480
rect 39028 4428 39080 4480
rect 41696 4471 41748 4480
rect 41696 4437 41705 4471
rect 41705 4437 41739 4471
rect 41739 4437 41748 4471
rect 41696 4428 41748 4437
rect 41880 4428 41932 4480
rect 45284 4564 45336 4616
rect 48780 4607 48832 4616
rect 48780 4573 48789 4607
rect 48789 4573 48823 4607
rect 48823 4573 48832 4607
rect 48780 4564 48832 4573
rect 77576 4607 77628 4616
rect 77576 4573 77585 4607
rect 77585 4573 77619 4607
rect 77619 4573 77628 4607
rect 77576 4564 77628 4573
rect 44456 4428 44508 4480
rect 48504 4496 48556 4548
rect 47860 4428 47912 4480
rect 48412 4428 48464 4480
rect 49700 4428 49752 4480
rect 5794 4326 5846 4378
rect 5858 4326 5910 4378
rect 5922 4326 5974 4378
rect 5986 4326 6038 4378
rect 6050 4326 6102 4378
rect 36514 4326 36566 4378
rect 36578 4326 36630 4378
rect 36642 4326 36694 4378
rect 36706 4326 36758 4378
rect 36770 4326 36822 4378
rect 67234 4326 67286 4378
rect 67298 4326 67350 4378
rect 67362 4326 67414 4378
rect 67426 4326 67478 4378
rect 67490 4326 67542 4378
rect 7472 4224 7524 4276
rect 9128 4224 9180 4276
rect 14004 4224 14056 4276
rect 17132 4224 17184 4276
rect 17776 4224 17828 4276
rect 19984 4224 20036 4276
rect 20536 4224 20588 4276
rect 21916 4224 21968 4276
rect 22468 4224 22520 4276
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 6460 4131 6512 4140
rect 6460 4097 6469 4131
rect 6469 4097 6503 4131
rect 6503 4097 6512 4131
rect 6460 4088 6512 4097
rect 8576 4156 8628 4208
rect 9772 4156 9824 4208
rect 12440 4156 12492 4208
rect 12808 4156 12860 4208
rect 13176 4156 13228 4208
rect 14832 4156 14884 4208
rect 16304 4156 16356 4208
rect 16764 4156 16816 4208
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 7840 4088 7892 4097
rect 9956 4088 10008 4140
rect 10508 4088 10560 4140
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 12256 4131 12308 4140
rect 12256 4097 12265 4131
rect 12265 4097 12299 4131
rect 12299 4097 12308 4131
rect 12256 4088 12308 4097
rect 3792 4020 3844 4072
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 9496 4020 9548 4029
rect 9772 4020 9824 4072
rect 10048 4063 10100 4072
rect 10048 4029 10057 4063
rect 10057 4029 10091 4063
rect 10091 4029 10100 4063
rect 10048 4020 10100 4029
rect 10416 4020 10468 4072
rect 14096 4088 14148 4140
rect 14188 4088 14240 4140
rect 14740 4088 14792 4140
rect 17592 4131 17644 4140
rect 17592 4097 17601 4131
rect 17601 4097 17635 4131
rect 17635 4097 17644 4131
rect 17592 4088 17644 4097
rect 18420 4088 18472 4140
rect 13728 4020 13780 4072
rect 14372 4063 14424 4072
rect 14372 4029 14381 4063
rect 14381 4029 14415 4063
rect 14415 4029 14424 4063
rect 14372 4020 14424 4029
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 15936 4063 15988 4072
rect 15936 4029 15945 4063
rect 15945 4029 15979 4063
rect 15979 4029 15988 4063
rect 15936 4020 15988 4029
rect 17500 4020 17552 4072
rect 22744 4156 22796 4208
rect 23204 4224 23256 4276
rect 19892 4131 19944 4140
rect 19892 4097 19901 4131
rect 19901 4097 19935 4131
rect 19935 4097 19944 4131
rect 19892 4088 19944 4097
rect 21088 4088 21140 4140
rect 21640 4088 21692 4140
rect 23388 4131 23440 4140
rect 23388 4097 23397 4131
rect 23397 4097 23431 4131
rect 23431 4097 23440 4131
rect 23388 4088 23440 4097
rect 23848 4156 23900 4208
rect 24308 4224 24360 4276
rect 24032 4156 24084 4208
rect 24952 4156 25004 4208
rect 27712 4224 27764 4276
rect 35624 4224 35676 4276
rect 35900 4224 35952 4276
rect 37372 4224 37424 4276
rect 37556 4224 37608 4276
rect 42340 4224 42392 4276
rect 42524 4224 42576 4276
rect 43996 4224 44048 4276
rect 48320 4267 48372 4276
rect 48320 4233 48329 4267
rect 48329 4233 48363 4267
rect 48363 4233 48372 4267
rect 48320 4224 48372 4233
rect 48780 4224 48832 4276
rect 26976 4156 27028 4208
rect 20260 4063 20312 4072
rect 20260 4029 20269 4063
rect 20269 4029 20303 4063
rect 20303 4029 20312 4063
rect 20260 4020 20312 4029
rect 21364 4063 21416 4072
rect 21364 4029 21373 4063
rect 21373 4029 21407 4063
rect 21407 4029 21416 4063
rect 21364 4020 21416 4029
rect 21732 4020 21784 4072
rect 22284 4020 22336 4072
rect 23664 4020 23716 4072
rect 11980 3952 12032 4004
rect 8484 3884 8536 3936
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 9128 3884 9180 3936
rect 17316 3952 17368 4004
rect 18144 3952 18196 4004
rect 18604 3952 18656 4004
rect 15752 3927 15804 3936
rect 15752 3893 15761 3927
rect 15761 3893 15795 3927
rect 15795 3893 15804 3927
rect 15752 3884 15804 3893
rect 16120 3884 16172 3936
rect 16580 3884 16632 3936
rect 22376 3952 22428 4004
rect 22744 3995 22796 4004
rect 22744 3961 22753 3995
rect 22753 3961 22787 3995
rect 22787 3961 22796 3995
rect 22744 3952 22796 3961
rect 20444 3884 20496 3936
rect 21824 3927 21876 3936
rect 21824 3893 21833 3927
rect 21833 3893 21867 3927
rect 21867 3893 21876 3927
rect 21824 3884 21876 3893
rect 21916 3884 21968 3936
rect 23112 3884 23164 3936
rect 23940 4131 23992 4140
rect 23940 4097 23949 4131
rect 23949 4097 23983 4131
rect 23983 4097 23992 4131
rect 23940 4088 23992 4097
rect 24216 4131 24268 4140
rect 24216 4097 24225 4131
rect 24225 4097 24259 4131
rect 24259 4097 24268 4131
rect 24216 4088 24268 4097
rect 24124 4020 24176 4072
rect 24584 4020 24636 4072
rect 26424 4088 26476 4140
rect 28264 4156 28316 4208
rect 28540 4156 28592 4208
rect 28080 4131 28132 4140
rect 28080 4097 28089 4131
rect 28089 4097 28123 4131
rect 28123 4097 28132 4131
rect 28080 4088 28132 4097
rect 26148 4020 26200 4072
rect 26884 4063 26936 4072
rect 26884 4029 26893 4063
rect 26893 4029 26927 4063
rect 26927 4029 26936 4063
rect 26884 4020 26936 4029
rect 28724 4088 28776 4140
rect 29000 4088 29052 4140
rect 29368 4088 29420 4140
rect 29552 4156 29604 4208
rect 35164 4156 35216 4208
rect 35256 4156 35308 4208
rect 38108 4156 38160 4208
rect 38200 4156 38252 4208
rect 38384 4156 38436 4208
rect 30840 4131 30892 4140
rect 30840 4097 30849 4131
rect 30849 4097 30883 4131
rect 30883 4097 30892 4131
rect 30840 4088 30892 4097
rect 30932 4088 30984 4140
rect 28908 4020 28960 4072
rect 29092 4063 29144 4072
rect 29092 4029 29101 4063
rect 29101 4029 29135 4063
rect 29135 4029 29144 4063
rect 29092 4020 29144 4029
rect 29736 4020 29788 4072
rect 25596 3884 25648 3936
rect 27896 3927 27948 3936
rect 27896 3893 27905 3927
rect 27905 3893 27939 3927
rect 27939 3893 27948 3927
rect 27896 3884 27948 3893
rect 30196 3952 30248 4004
rect 30748 4020 30800 4072
rect 31944 4063 31996 4072
rect 31944 4029 31953 4063
rect 31953 4029 31987 4063
rect 31987 4029 31996 4063
rect 31944 4020 31996 4029
rect 32404 4020 32456 4072
rect 33784 4088 33836 4140
rect 34060 4131 34112 4140
rect 34060 4097 34069 4131
rect 34069 4097 34103 4131
rect 34103 4097 34112 4131
rect 34060 4088 34112 4097
rect 36636 4088 36688 4140
rect 37464 4088 37516 4140
rect 37556 4088 37608 4140
rect 38568 4131 38620 4140
rect 38568 4097 38577 4131
rect 38577 4097 38611 4131
rect 38611 4097 38620 4131
rect 38568 4088 38620 4097
rect 39212 4088 39264 4140
rect 39488 4088 39540 4140
rect 40408 4131 40460 4140
rect 40408 4097 40417 4131
rect 40417 4097 40451 4131
rect 40451 4097 40460 4131
rect 40408 4088 40460 4097
rect 40500 4131 40552 4140
rect 40500 4097 40509 4131
rect 40509 4097 40543 4131
rect 40543 4097 40552 4131
rect 40500 4088 40552 4097
rect 43352 4156 43404 4208
rect 33416 4063 33468 4072
rect 33416 4029 33425 4063
rect 33425 4029 33459 4063
rect 33459 4029 33468 4063
rect 33416 4020 33468 4029
rect 35256 4063 35308 4072
rect 35256 4029 35265 4063
rect 35265 4029 35299 4063
rect 35299 4029 35308 4063
rect 35256 4020 35308 4029
rect 29920 3927 29972 3936
rect 29920 3893 29929 3927
rect 29929 3893 29963 3927
rect 29963 3893 29972 3927
rect 29920 3884 29972 3893
rect 30104 3884 30156 3936
rect 31852 3952 31904 4004
rect 33232 3995 33284 4004
rect 33232 3961 33241 3995
rect 33241 3961 33275 3995
rect 33275 3961 33284 3995
rect 33232 3952 33284 3961
rect 33324 3952 33376 4004
rect 36084 4020 36136 4072
rect 36728 4020 36780 4072
rect 36912 4063 36964 4072
rect 36912 4029 36921 4063
rect 36921 4029 36955 4063
rect 36955 4029 36964 4063
rect 36912 4020 36964 4029
rect 37740 4063 37792 4072
rect 37740 4029 37749 4063
rect 37749 4029 37783 4063
rect 37783 4029 37792 4063
rect 37740 4020 37792 4029
rect 38108 4020 38160 4072
rect 40316 4020 40368 4072
rect 42064 4020 42116 4072
rect 42524 4131 42576 4140
rect 42524 4097 42533 4131
rect 42533 4097 42567 4131
rect 42567 4097 42576 4131
rect 42524 4088 42576 4097
rect 42708 4088 42760 4140
rect 43260 4088 43312 4140
rect 46480 4088 46532 4140
rect 42800 4020 42852 4072
rect 42892 4063 42944 4072
rect 42892 4029 42901 4063
rect 42901 4029 42935 4063
rect 42935 4029 42944 4063
rect 42892 4020 42944 4029
rect 43076 4020 43128 4072
rect 31392 3927 31444 3936
rect 31392 3893 31401 3927
rect 31401 3893 31435 3927
rect 31435 3893 31444 3927
rect 31392 3884 31444 3893
rect 32496 3884 32548 3936
rect 33876 3884 33928 3936
rect 36728 3884 36780 3936
rect 39948 3884 40000 3936
rect 41236 3884 41288 3936
rect 42340 3884 42392 3936
rect 42800 3884 42852 3936
rect 43812 3884 43864 3936
rect 44180 4063 44232 4072
rect 44180 4029 44189 4063
rect 44189 4029 44223 4063
rect 44223 4029 44232 4063
rect 44180 4020 44232 4029
rect 44732 4063 44784 4072
rect 44732 4029 44741 4063
rect 44741 4029 44775 4063
rect 44775 4029 44784 4063
rect 44732 4020 44784 4029
rect 45652 4063 45704 4072
rect 45652 4029 45661 4063
rect 45661 4029 45695 4063
rect 45695 4029 45704 4063
rect 45652 4020 45704 4029
rect 48044 4131 48096 4140
rect 48044 4097 48053 4131
rect 48053 4097 48087 4131
rect 48087 4097 48096 4131
rect 48044 4088 48096 4097
rect 48504 4131 48556 4140
rect 48504 4097 48513 4131
rect 48513 4097 48547 4131
rect 48547 4097 48556 4131
rect 48504 4088 48556 4097
rect 74632 4088 74684 4140
rect 47584 3952 47636 4004
rect 44824 3884 44876 3936
rect 44916 3927 44968 3936
rect 44916 3893 44925 3927
rect 44925 3893 44959 3927
rect 44959 3893 44968 3927
rect 44916 3884 44968 3893
rect 46388 3884 46440 3936
rect 53196 4020 53248 4072
rect 53840 4063 53892 4072
rect 53840 4029 53849 4063
rect 53849 4029 53883 4063
rect 53883 4029 53892 4063
rect 53840 4020 53892 4029
rect 65432 4020 65484 4072
rect 68652 4020 68704 4072
rect 69296 4063 69348 4072
rect 69296 4029 69305 4063
rect 69305 4029 69339 4063
rect 69339 4029 69348 4063
rect 69296 4020 69348 4029
rect 71688 4020 71740 4072
rect 74264 4020 74316 4072
rect 76564 4020 76616 4072
rect 77024 4063 77076 4072
rect 77024 4029 77033 4063
rect 77033 4029 77067 4063
rect 77067 4029 77076 4063
rect 77024 4020 77076 4029
rect 51356 3884 51408 3936
rect 52828 3884 52880 3936
rect 54024 3884 54076 3936
rect 66260 3884 66312 3936
rect 68284 3884 68336 3936
rect 69480 3884 69532 3936
rect 73712 3884 73764 3936
rect 5134 3782 5186 3834
rect 5198 3782 5250 3834
rect 5262 3782 5314 3834
rect 5326 3782 5378 3834
rect 5390 3782 5442 3834
rect 35854 3782 35906 3834
rect 35918 3782 35970 3834
rect 35982 3782 36034 3834
rect 36046 3782 36098 3834
rect 36110 3782 36162 3834
rect 66574 3782 66626 3834
rect 66638 3782 66690 3834
rect 66702 3782 66754 3834
rect 66766 3782 66818 3834
rect 66830 3782 66882 3834
rect 6644 3680 6696 3732
rect 8576 3680 8628 3732
rect 13728 3723 13780 3732
rect 13728 3689 13737 3723
rect 13737 3689 13771 3723
rect 13771 3689 13780 3723
rect 13728 3680 13780 3689
rect 14832 3723 14884 3732
rect 14832 3689 14841 3723
rect 14841 3689 14875 3723
rect 14875 3689 14884 3723
rect 14832 3680 14884 3689
rect 15292 3680 15344 3732
rect 15936 3680 15988 3732
rect 6828 3544 6880 3596
rect 5264 3519 5316 3528
rect 5264 3485 5273 3519
rect 5273 3485 5307 3519
rect 5307 3485 5316 3519
rect 5264 3476 5316 3485
rect 8760 3476 8812 3528
rect 9864 3544 9916 3596
rect 10416 3544 10468 3596
rect 10876 3587 10928 3596
rect 10876 3553 10885 3587
rect 10885 3553 10919 3587
rect 10919 3553 10928 3587
rect 10876 3544 10928 3553
rect 12348 3544 12400 3596
rect 4160 3408 4212 3460
rect 10048 3476 10100 3528
rect 10508 3408 10560 3460
rect 8852 3340 8904 3392
rect 9036 3340 9088 3392
rect 9588 3340 9640 3392
rect 10416 3340 10468 3392
rect 10968 3340 11020 3392
rect 11520 3383 11572 3392
rect 11520 3349 11529 3383
rect 11529 3349 11563 3383
rect 11563 3349 11572 3383
rect 11520 3340 11572 3349
rect 12348 3408 12400 3460
rect 13084 3340 13136 3392
rect 14096 3544 14148 3596
rect 16396 3612 16448 3664
rect 19892 3680 19944 3732
rect 20076 3680 20128 3732
rect 27712 3680 27764 3732
rect 28080 3680 28132 3732
rect 29552 3680 29604 3732
rect 31300 3680 31352 3732
rect 33048 3680 33100 3732
rect 33968 3680 34020 3732
rect 34704 3723 34756 3732
rect 34704 3689 34713 3723
rect 34713 3689 34747 3723
rect 34747 3689 34756 3723
rect 34704 3680 34756 3689
rect 16764 3544 16816 3596
rect 17868 3544 17920 3596
rect 18144 3587 18196 3596
rect 18144 3553 18153 3587
rect 18153 3553 18187 3587
rect 18187 3553 18196 3587
rect 18144 3544 18196 3553
rect 20076 3544 20128 3596
rect 20996 3544 21048 3596
rect 22376 3612 22428 3664
rect 24952 3612 25004 3664
rect 25320 3612 25372 3664
rect 25688 3612 25740 3664
rect 26516 3655 26568 3664
rect 26516 3621 26525 3655
rect 26525 3621 26559 3655
rect 26559 3621 26568 3655
rect 26516 3612 26568 3621
rect 27988 3612 28040 3664
rect 14004 3476 14056 3528
rect 14464 3476 14516 3528
rect 14648 3519 14700 3528
rect 14648 3485 14657 3519
rect 14657 3485 14691 3519
rect 14691 3485 14700 3519
rect 14648 3476 14700 3485
rect 15200 3476 15252 3528
rect 15568 3519 15620 3528
rect 15568 3485 15577 3519
rect 15577 3485 15611 3519
rect 15611 3485 15620 3519
rect 15568 3476 15620 3485
rect 16304 3519 16356 3528
rect 16304 3485 16313 3519
rect 16313 3485 16347 3519
rect 16347 3485 16356 3519
rect 16304 3476 16356 3485
rect 14740 3408 14792 3460
rect 14924 3408 14976 3460
rect 19892 3476 19944 3528
rect 26424 3544 26476 3596
rect 27436 3544 27488 3596
rect 23388 3476 23440 3528
rect 24032 3476 24084 3528
rect 25228 3476 25280 3528
rect 25320 3519 25372 3528
rect 25320 3485 25329 3519
rect 25329 3485 25363 3519
rect 25363 3485 25372 3519
rect 25320 3476 25372 3485
rect 20260 3451 20312 3460
rect 14556 3340 14608 3392
rect 15936 3383 15988 3392
rect 15936 3349 15945 3383
rect 15945 3349 15979 3383
rect 15979 3349 15988 3383
rect 15936 3340 15988 3349
rect 20260 3417 20269 3451
rect 20269 3417 20303 3451
rect 20303 3417 20312 3451
rect 20260 3408 20312 3417
rect 21272 3408 21324 3460
rect 21916 3408 21968 3460
rect 22192 3451 22244 3460
rect 22192 3417 22201 3451
rect 22201 3417 22235 3451
rect 22235 3417 22244 3451
rect 22192 3408 22244 3417
rect 22468 3408 22520 3460
rect 28080 3476 28132 3528
rect 25596 3451 25648 3460
rect 25596 3417 25605 3451
rect 25605 3417 25639 3451
rect 25639 3417 25648 3451
rect 25596 3408 25648 3417
rect 25872 3408 25924 3460
rect 26148 3451 26200 3460
rect 26148 3417 26157 3451
rect 26157 3417 26191 3451
rect 26191 3417 26200 3451
rect 26148 3408 26200 3417
rect 27252 3408 27304 3460
rect 28448 3655 28500 3664
rect 28448 3621 28457 3655
rect 28457 3621 28491 3655
rect 28491 3621 28500 3655
rect 28448 3612 28500 3621
rect 30380 3612 30432 3664
rect 32036 3655 32088 3664
rect 32036 3621 32045 3655
rect 32045 3621 32079 3655
rect 32079 3621 32088 3655
rect 32036 3612 32088 3621
rect 34980 3612 35032 3664
rect 29368 3587 29420 3596
rect 29368 3553 29377 3587
rect 29377 3553 29411 3587
rect 29411 3553 29420 3587
rect 29368 3544 29420 3553
rect 30104 3544 30156 3596
rect 30656 3544 30708 3596
rect 31208 3544 31260 3596
rect 32128 3544 32180 3596
rect 32588 3544 32640 3596
rect 33600 3544 33652 3596
rect 36912 3680 36964 3732
rect 40316 3680 40368 3732
rect 41512 3680 41564 3732
rect 41880 3680 41932 3732
rect 44916 3680 44968 3732
rect 45560 3723 45612 3732
rect 45560 3689 45569 3723
rect 45569 3689 45603 3723
rect 45603 3689 45612 3723
rect 45560 3680 45612 3689
rect 46756 3680 46808 3732
rect 48044 3680 48096 3732
rect 53196 3723 53248 3732
rect 53196 3689 53205 3723
rect 53205 3689 53239 3723
rect 53239 3689 53248 3723
rect 53196 3680 53248 3689
rect 68652 3723 68704 3732
rect 68652 3689 68661 3723
rect 68661 3689 68695 3723
rect 68695 3689 68704 3723
rect 68652 3680 68704 3689
rect 71688 3723 71740 3732
rect 71688 3689 71697 3723
rect 71697 3689 71731 3723
rect 71731 3689 71740 3723
rect 71688 3680 71740 3689
rect 77576 3723 77628 3732
rect 77576 3689 77585 3723
rect 77585 3689 77619 3723
rect 77619 3689 77628 3723
rect 77576 3680 77628 3689
rect 28724 3519 28776 3528
rect 28724 3485 28733 3519
rect 28733 3485 28767 3519
rect 28767 3485 28776 3519
rect 28724 3476 28776 3485
rect 29092 3519 29144 3528
rect 29092 3485 29101 3519
rect 29101 3485 29135 3519
rect 29135 3485 29144 3519
rect 29092 3476 29144 3485
rect 31116 3476 31168 3528
rect 31668 3519 31720 3528
rect 31668 3485 31677 3519
rect 31677 3485 31711 3519
rect 31711 3485 31720 3519
rect 31668 3476 31720 3485
rect 30380 3408 30432 3460
rect 18052 3340 18104 3392
rect 18604 3340 18656 3392
rect 19340 3340 19392 3392
rect 20812 3340 20864 3392
rect 21456 3340 21508 3392
rect 24216 3340 24268 3392
rect 24768 3340 24820 3392
rect 25412 3383 25464 3392
rect 25412 3349 25421 3383
rect 25421 3349 25455 3383
rect 25455 3349 25464 3383
rect 25412 3340 25464 3349
rect 25688 3383 25740 3392
rect 25688 3349 25697 3383
rect 25697 3349 25731 3383
rect 25731 3349 25740 3383
rect 25688 3340 25740 3349
rect 26240 3340 26292 3392
rect 29460 3340 29512 3392
rect 30840 3340 30892 3392
rect 34152 3519 34204 3528
rect 34152 3485 34161 3519
rect 34161 3485 34195 3519
rect 34195 3485 34204 3519
rect 34152 3476 34204 3485
rect 34888 3476 34940 3528
rect 32680 3408 32732 3460
rect 33048 3408 33100 3460
rect 33876 3408 33928 3460
rect 35716 3519 35768 3528
rect 35716 3485 35725 3519
rect 35725 3485 35759 3519
rect 35759 3485 35768 3519
rect 35716 3476 35768 3485
rect 38568 3587 38620 3596
rect 38568 3553 38577 3587
rect 38577 3553 38611 3587
rect 38611 3553 38620 3587
rect 38568 3544 38620 3553
rect 42524 3612 42576 3664
rect 43812 3612 43864 3664
rect 36268 3476 36320 3528
rect 37188 3476 37240 3528
rect 37280 3519 37332 3528
rect 37280 3485 37289 3519
rect 37289 3485 37323 3519
rect 37323 3485 37332 3519
rect 37280 3476 37332 3485
rect 39120 3519 39172 3528
rect 39120 3485 39129 3519
rect 39129 3485 39163 3519
rect 39163 3485 39172 3519
rect 39120 3476 39172 3485
rect 40592 3519 40644 3528
rect 40592 3485 40601 3519
rect 40601 3485 40635 3519
rect 40635 3485 40644 3519
rect 40592 3476 40644 3485
rect 33508 3340 33560 3392
rect 34152 3340 34204 3392
rect 35164 3383 35216 3392
rect 35164 3349 35173 3383
rect 35173 3349 35207 3383
rect 35207 3349 35216 3383
rect 35164 3340 35216 3349
rect 38476 3408 38528 3460
rect 39396 3451 39448 3460
rect 39396 3417 39405 3451
rect 39405 3417 39439 3451
rect 39439 3417 39448 3451
rect 39396 3408 39448 3417
rect 35716 3340 35768 3392
rect 36084 3340 36136 3392
rect 40684 3340 40736 3392
rect 40776 3383 40828 3392
rect 40776 3349 40785 3383
rect 40785 3349 40819 3383
rect 40819 3349 40828 3383
rect 40776 3340 40828 3349
rect 41696 3544 41748 3596
rect 42248 3544 42300 3596
rect 46848 3544 46900 3596
rect 47860 3544 47912 3596
rect 48872 3587 48924 3596
rect 48872 3553 48881 3587
rect 48881 3553 48915 3587
rect 48915 3553 48924 3587
rect 48872 3544 48924 3553
rect 54024 3587 54076 3596
rect 54024 3553 54033 3587
rect 54033 3553 54067 3587
rect 54067 3553 54076 3587
rect 54024 3544 54076 3553
rect 69480 3587 69532 3596
rect 69480 3553 69489 3587
rect 69489 3553 69523 3587
rect 69523 3553 69532 3587
rect 69480 3544 69532 3553
rect 73712 3587 73764 3596
rect 73712 3553 73721 3587
rect 73721 3553 73755 3587
rect 73755 3553 73764 3587
rect 73712 3544 73764 3553
rect 77024 3587 77076 3596
rect 77024 3553 77033 3587
rect 77033 3553 77067 3587
rect 77067 3553 77076 3587
rect 77024 3544 77076 3553
rect 41052 3519 41104 3528
rect 41052 3485 41061 3519
rect 41061 3485 41095 3519
rect 41095 3485 41104 3519
rect 41052 3476 41104 3485
rect 41236 3519 41288 3528
rect 41236 3485 41245 3519
rect 41245 3485 41279 3519
rect 41279 3485 41288 3519
rect 41236 3476 41288 3485
rect 41328 3519 41380 3528
rect 41328 3485 41337 3519
rect 41337 3485 41371 3519
rect 41371 3485 41380 3519
rect 41328 3476 41380 3485
rect 42524 3408 42576 3460
rect 43260 3340 43312 3392
rect 43352 3340 43404 3392
rect 43904 3519 43956 3528
rect 43904 3485 43913 3519
rect 43913 3485 43947 3519
rect 43947 3485 43956 3519
rect 43904 3476 43956 3485
rect 45192 3408 45244 3460
rect 47124 3476 47176 3528
rect 47952 3519 48004 3528
rect 47952 3485 47961 3519
rect 47961 3485 47995 3519
rect 47995 3485 48004 3519
rect 47952 3476 48004 3485
rect 50804 3476 50856 3528
rect 53012 3519 53064 3528
rect 53012 3485 53021 3519
rect 53021 3485 53055 3519
rect 53055 3485 53064 3519
rect 53012 3476 53064 3485
rect 48136 3383 48188 3392
rect 48136 3349 48145 3383
rect 48145 3349 48179 3383
rect 48179 3349 48188 3383
rect 48136 3340 48188 3349
rect 50528 3408 50580 3460
rect 57336 3408 57388 3460
rect 59452 3519 59504 3528
rect 59452 3485 59461 3519
rect 59461 3485 59495 3519
rect 59495 3485 59504 3519
rect 59452 3476 59504 3485
rect 60924 3408 60976 3460
rect 63408 3519 63460 3528
rect 63408 3485 63417 3519
rect 63417 3485 63451 3519
rect 63451 3485 63460 3519
rect 63408 3476 63460 3485
rect 64512 3519 64564 3528
rect 64512 3485 64521 3519
rect 64521 3485 64555 3519
rect 64555 3485 64564 3519
rect 64512 3476 64564 3485
rect 68468 3519 68520 3528
rect 68468 3485 68477 3519
rect 68477 3485 68511 3519
rect 68511 3485 68520 3519
rect 68468 3476 68520 3485
rect 72976 3519 73028 3528
rect 72976 3485 72985 3519
rect 72985 3485 73019 3519
rect 73019 3485 73028 3519
rect 72976 3476 73028 3485
rect 74448 3476 74500 3528
rect 76656 3519 76708 3528
rect 76656 3485 76665 3519
rect 76665 3485 76699 3519
rect 76699 3485 76708 3519
rect 76656 3476 76708 3485
rect 75460 3451 75512 3460
rect 75460 3417 75469 3451
rect 75469 3417 75503 3451
rect 75503 3417 75512 3451
rect 75460 3408 75512 3417
rect 49976 3340 50028 3392
rect 56048 3340 56100 3392
rect 57428 3383 57480 3392
rect 57428 3349 57437 3383
rect 57437 3349 57471 3383
rect 57471 3349 57480 3383
rect 57428 3340 57480 3349
rect 58624 3340 58676 3392
rect 61108 3340 61160 3392
rect 62764 3340 62816 3392
rect 64880 3340 64932 3392
rect 71504 3340 71556 3392
rect 73252 3340 73304 3392
rect 74540 3383 74592 3392
rect 74540 3349 74549 3383
rect 74549 3349 74583 3383
rect 74583 3349 74592 3383
rect 74540 3340 74592 3349
rect 5794 3238 5846 3290
rect 5858 3238 5910 3290
rect 5922 3238 5974 3290
rect 5986 3238 6038 3290
rect 6050 3238 6102 3290
rect 36514 3238 36566 3290
rect 36578 3238 36630 3290
rect 36642 3238 36694 3290
rect 36706 3238 36758 3290
rect 36770 3238 36822 3290
rect 67234 3238 67286 3290
rect 67298 3238 67350 3290
rect 67362 3238 67414 3290
rect 67426 3238 67478 3290
rect 67490 3238 67542 3290
rect 3792 3179 3844 3188
rect 3792 3145 3801 3179
rect 3801 3145 3835 3179
rect 3835 3145 3844 3179
rect 3792 3136 3844 3145
rect 5264 3136 5316 3188
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 9220 3136 9272 3188
rect 9956 3136 10008 3188
rect 10416 3136 10468 3188
rect 10140 3068 10192 3120
rect 10784 3111 10836 3120
rect 10784 3077 10793 3111
rect 10793 3077 10827 3111
rect 10827 3077 10836 3111
rect 10784 3068 10836 3077
rect 11244 3068 11296 3120
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 8484 3000 8536 3052
rect 9956 3000 10008 3052
rect 10508 3043 10560 3052
rect 10508 3009 10517 3043
rect 10517 3009 10551 3043
rect 10551 3009 10560 3043
rect 10508 3000 10560 3009
rect 12164 3136 12216 3188
rect 12348 3136 12400 3188
rect 12624 3111 12676 3120
rect 12624 3077 12633 3111
rect 12633 3077 12667 3111
rect 12667 3077 12676 3111
rect 12624 3068 12676 3077
rect 12992 3136 13044 3188
rect 13084 3136 13136 3188
rect 14924 3136 14976 3188
rect 15936 3136 15988 3188
rect 16856 3136 16908 3188
rect 17316 3136 17368 3188
rect 17592 3179 17644 3188
rect 17592 3145 17601 3179
rect 17601 3145 17635 3179
rect 17635 3145 17644 3179
rect 17592 3136 17644 3145
rect 18604 3136 18656 3188
rect 13820 3068 13872 3120
rect 5540 2932 5592 2984
rect 5632 2975 5684 2984
rect 5632 2941 5641 2975
rect 5641 2941 5675 2975
rect 5675 2941 5684 2975
rect 5632 2932 5684 2941
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 5724 2932 5776 2941
rect 6920 2932 6972 2984
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 7656 2932 7708 2984
rect 9128 2975 9180 2984
rect 9128 2941 9137 2975
rect 9137 2941 9171 2975
rect 9171 2941 9180 2975
rect 9128 2932 9180 2941
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 15108 3068 15160 3120
rect 17960 3068 18012 3120
rect 19340 3068 19392 3120
rect 18052 3043 18104 3052
rect 18052 3009 18061 3043
rect 18061 3009 18095 3043
rect 18095 3009 18104 3043
rect 18052 3000 18104 3009
rect 6460 2839 6512 2848
rect 6460 2805 6469 2839
rect 6469 2805 6503 2839
rect 6503 2805 6512 2839
rect 6460 2796 6512 2805
rect 10140 2796 10192 2848
rect 12256 2796 12308 2848
rect 15568 2932 15620 2984
rect 17316 2932 17368 2984
rect 21088 3136 21140 3188
rect 22652 3136 22704 3188
rect 23020 3179 23072 3188
rect 23020 3145 23029 3179
rect 23029 3145 23063 3179
rect 23063 3145 23072 3179
rect 23020 3136 23072 3145
rect 21824 3000 21876 3052
rect 22008 3000 22060 3052
rect 19708 2932 19760 2984
rect 24492 3111 24544 3120
rect 24492 3077 24501 3111
rect 24501 3077 24535 3111
rect 24535 3077 24544 3111
rect 24492 3068 24544 3077
rect 25964 3136 26016 3188
rect 26976 3179 27028 3188
rect 26976 3145 26985 3179
rect 26985 3145 27019 3179
rect 27019 3145 27028 3179
rect 26976 3136 27028 3145
rect 27436 3179 27488 3188
rect 27436 3145 27445 3179
rect 27445 3145 27479 3179
rect 27479 3145 27488 3179
rect 27436 3136 27488 3145
rect 28448 3136 28500 3188
rect 28540 3179 28592 3188
rect 28540 3145 28549 3179
rect 28549 3145 28583 3179
rect 28583 3145 28592 3179
rect 28540 3136 28592 3145
rect 30748 3136 30800 3188
rect 30840 3136 30892 3188
rect 36084 3136 36136 3188
rect 23388 3000 23440 3052
rect 24768 3043 24820 3052
rect 24768 3009 24777 3043
rect 24777 3009 24811 3043
rect 24811 3009 24820 3043
rect 24768 3000 24820 3009
rect 24860 3043 24912 3052
rect 24860 3009 24869 3043
rect 24869 3009 24903 3043
rect 24903 3009 24912 3043
rect 24860 3000 24912 3009
rect 23756 2932 23808 2984
rect 25228 3043 25280 3052
rect 25228 3009 25237 3043
rect 25237 3009 25271 3043
rect 25271 3009 25280 3043
rect 25228 3000 25280 3009
rect 25504 3068 25556 3120
rect 26056 3068 26108 3120
rect 28724 3068 28776 3120
rect 29552 3068 29604 3120
rect 30012 3111 30064 3120
rect 30012 3077 30021 3111
rect 30021 3077 30055 3111
rect 30055 3077 30064 3111
rect 30012 3068 30064 3077
rect 30104 3068 30156 3120
rect 26700 3000 26752 3052
rect 26884 3043 26936 3052
rect 26884 3009 26893 3043
rect 26893 3009 26927 3043
rect 26927 3009 26936 3043
rect 26884 3000 26936 3009
rect 27344 3043 27396 3052
rect 27344 3009 27353 3043
rect 27353 3009 27387 3043
rect 27387 3009 27396 3043
rect 27344 3000 27396 3009
rect 27988 3043 28040 3052
rect 27988 3009 27997 3043
rect 27997 3009 28031 3043
rect 28031 3009 28040 3043
rect 27988 3000 28040 3009
rect 30564 3068 30616 3120
rect 30932 3068 30984 3120
rect 32312 3068 32364 3120
rect 32772 3068 32824 3120
rect 26424 2975 26476 2984
rect 26424 2941 26433 2975
rect 26433 2941 26467 2975
rect 26467 2941 26476 2975
rect 26424 2932 26476 2941
rect 26792 2932 26844 2984
rect 28632 2932 28684 2984
rect 31024 3000 31076 3052
rect 31300 3000 31352 3052
rect 32680 3043 32732 3052
rect 32680 3009 32689 3043
rect 32689 3009 32723 3043
rect 32723 3009 32732 3043
rect 32680 3000 32732 3009
rect 33968 3068 34020 3120
rect 35532 3068 35584 3120
rect 35624 3111 35676 3120
rect 35624 3077 35633 3111
rect 35633 3077 35667 3111
rect 35667 3077 35676 3111
rect 35624 3068 35676 3077
rect 33876 3043 33928 3052
rect 33876 3009 33885 3043
rect 33885 3009 33919 3043
rect 33919 3009 33928 3043
rect 33876 3000 33928 3009
rect 37924 3136 37976 3188
rect 38660 3111 38712 3120
rect 38660 3077 38669 3111
rect 38669 3077 38703 3111
rect 38703 3077 38712 3111
rect 38660 3068 38712 3077
rect 42064 3179 42116 3188
rect 42064 3145 42073 3179
rect 42073 3145 42107 3179
rect 42107 3145 42116 3179
rect 42064 3136 42116 3145
rect 42984 3136 43036 3188
rect 44364 3136 44416 3188
rect 45284 3136 45336 3188
rect 46940 3136 46992 3188
rect 48320 3136 48372 3188
rect 29920 2932 29972 2984
rect 31208 2932 31260 2984
rect 31852 2932 31904 2984
rect 33600 2975 33652 2984
rect 33600 2941 33609 2975
rect 33609 2941 33643 2975
rect 33643 2941 33652 2975
rect 33600 2932 33652 2941
rect 33784 2932 33836 2984
rect 24860 2864 24912 2916
rect 26516 2864 26568 2916
rect 14740 2796 14792 2848
rect 18420 2796 18472 2848
rect 21824 2839 21876 2848
rect 21824 2805 21833 2839
rect 21833 2805 21867 2839
rect 21867 2805 21876 2839
rect 21824 2796 21876 2805
rect 22836 2796 22888 2848
rect 24400 2796 24452 2848
rect 26976 2796 27028 2848
rect 29000 2864 29052 2916
rect 34152 2907 34204 2916
rect 29276 2796 29328 2848
rect 30288 2796 30340 2848
rect 30472 2796 30524 2848
rect 34152 2873 34161 2907
rect 34161 2873 34195 2907
rect 34195 2873 34204 2907
rect 34152 2864 34204 2873
rect 33048 2839 33100 2848
rect 33048 2805 33057 2839
rect 33057 2805 33091 2839
rect 33091 2805 33100 2839
rect 33048 2796 33100 2805
rect 34520 2796 34572 2848
rect 39764 3000 39816 3052
rect 43720 3068 43772 3120
rect 44180 3068 44232 3120
rect 42248 3043 42300 3052
rect 42248 3009 42257 3043
rect 42257 3009 42291 3043
rect 42291 3009 42300 3043
rect 42248 3000 42300 3009
rect 37464 2864 37516 2916
rect 35900 2796 35952 2848
rect 41144 2932 41196 2984
rect 42156 2932 42208 2984
rect 40408 2864 40460 2916
rect 40316 2796 40368 2848
rect 43076 2932 43128 2984
rect 43352 3043 43404 3052
rect 43352 3009 43361 3043
rect 43361 3009 43395 3043
rect 43395 3009 43404 3043
rect 43352 3000 43404 3009
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 46756 3043 46808 3052
rect 46756 3009 46765 3043
rect 46765 3009 46799 3043
rect 46799 3009 46808 3043
rect 46756 3000 46808 3009
rect 50804 3179 50856 3188
rect 50804 3145 50813 3179
rect 50813 3145 50847 3179
rect 50847 3145 50856 3179
rect 50804 3136 50856 3145
rect 53012 3136 53064 3188
rect 53840 3179 53892 3188
rect 53840 3145 53849 3179
rect 53849 3145 53883 3179
rect 53883 3145 53892 3179
rect 53840 3136 53892 3145
rect 57336 3179 57388 3188
rect 57336 3145 57345 3179
rect 57345 3145 57379 3179
rect 57379 3145 57388 3179
rect 57336 3136 57388 3145
rect 59452 3136 59504 3188
rect 60924 3179 60976 3188
rect 60924 3145 60933 3179
rect 60933 3145 60967 3179
rect 60967 3145 60976 3179
rect 60924 3136 60976 3145
rect 63408 3136 63460 3188
rect 64512 3179 64564 3188
rect 64512 3145 64521 3179
rect 64521 3145 64555 3179
rect 64555 3145 64564 3179
rect 64512 3136 64564 3145
rect 65432 3179 65484 3188
rect 65432 3145 65441 3179
rect 65441 3145 65475 3179
rect 65475 3145 65484 3179
rect 65432 3136 65484 3145
rect 68468 3136 68520 3188
rect 69296 3179 69348 3188
rect 69296 3145 69305 3179
rect 69305 3145 69339 3179
rect 69339 3145 69348 3179
rect 69296 3136 69348 3145
rect 74448 3179 74500 3188
rect 74448 3145 74457 3179
rect 74457 3145 74491 3179
rect 74491 3145 74500 3179
rect 74448 3136 74500 3145
rect 49792 3043 49844 3052
rect 49792 3009 49801 3043
rect 49801 3009 49835 3043
rect 49835 3009 49844 3043
rect 49792 3000 49844 3009
rect 51356 3043 51408 3052
rect 51356 3009 51365 3043
rect 51365 3009 51399 3043
rect 51399 3009 51408 3043
rect 51356 3000 51408 3009
rect 52092 3043 52144 3052
rect 52092 3009 52101 3043
rect 52101 3009 52135 3043
rect 52135 3009 52144 3043
rect 52092 3000 52144 3009
rect 54024 3043 54076 3052
rect 54024 3009 54033 3043
rect 54033 3009 54067 3043
rect 54067 3009 54076 3043
rect 54024 3000 54076 3009
rect 56048 3043 56100 3052
rect 56048 3009 56057 3043
rect 56057 3009 56091 3043
rect 56091 3009 56100 3043
rect 56048 3000 56100 3009
rect 57428 3043 57480 3052
rect 57428 3009 57437 3043
rect 57437 3009 57471 3043
rect 57471 3009 57480 3043
rect 57428 3000 57480 3009
rect 61108 3043 61160 3052
rect 61108 3009 61117 3043
rect 61117 3009 61151 3043
rect 61151 3009 61160 3043
rect 61108 3000 61160 3009
rect 61752 3043 61804 3052
rect 61752 3009 61761 3043
rect 61761 3009 61795 3043
rect 61795 3009 61804 3043
rect 61752 3000 61804 3009
rect 64880 3043 64932 3052
rect 64880 3009 64889 3043
rect 64889 3009 64923 3043
rect 64923 3009 64932 3043
rect 64880 3000 64932 3009
rect 65524 3043 65576 3052
rect 65524 3009 65533 3043
rect 65533 3009 65567 3043
rect 65567 3009 65576 3043
rect 65524 3000 65576 3009
rect 67640 3043 67692 3052
rect 67640 3009 67649 3043
rect 67649 3009 67683 3043
rect 67683 3009 67692 3043
rect 67640 3000 67692 3009
rect 70308 3068 70360 3120
rect 69480 3043 69532 3052
rect 69480 3009 69489 3043
rect 69489 3009 69523 3043
rect 69523 3009 69532 3043
rect 69480 3000 69532 3009
rect 71504 3043 71556 3052
rect 71504 3009 71513 3043
rect 71513 3009 71547 3043
rect 71547 3009 71556 3043
rect 71504 3000 71556 3009
rect 72608 3000 72660 3052
rect 74264 3043 74316 3052
rect 74264 3009 74273 3043
rect 74273 3009 74307 3043
rect 74307 3009 74316 3043
rect 74264 3000 74316 3009
rect 74540 3043 74592 3052
rect 74540 3009 74549 3043
rect 74549 3009 74583 3043
rect 74583 3009 74592 3043
rect 74540 3000 74592 3009
rect 76656 3043 76708 3052
rect 76656 3009 76665 3043
rect 76665 3009 76699 3043
rect 76699 3009 76708 3043
rect 76656 3000 76708 3009
rect 44180 2932 44232 2984
rect 45744 2932 45796 2984
rect 47676 2932 47728 2984
rect 49608 2932 49660 2984
rect 53472 2932 53524 2984
rect 61200 2932 61252 2984
rect 65064 2932 65116 2984
rect 68928 2932 68980 2984
rect 70860 2932 70912 2984
rect 74724 2932 74776 2984
rect 51540 2864 51592 2916
rect 66996 2864 67048 2916
rect 45284 2796 45336 2848
rect 55312 2796 55364 2848
rect 59268 2796 59320 2848
rect 70492 2796 70544 2848
rect 76196 2796 76248 2848
rect 5134 2694 5186 2746
rect 5198 2694 5250 2746
rect 5262 2694 5314 2746
rect 5326 2694 5378 2746
rect 5390 2694 5442 2746
rect 35854 2694 35906 2746
rect 35918 2694 35970 2746
rect 35982 2694 36034 2746
rect 36046 2694 36098 2746
rect 36110 2694 36162 2746
rect 66574 2694 66626 2746
rect 66638 2694 66690 2746
rect 66702 2694 66754 2746
rect 66766 2694 66818 2746
rect 66830 2694 66882 2746
rect 3884 2592 3936 2644
rect 7656 2592 7708 2644
rect 8576 2635 8628 2644
rect 8576 2601 8585 2635
rect 8585 2601 8619 2635
rect 8619 2601 8628 2635
rect 8576 2592 8628 2601
rect 11888 2592 11940 2644
rect 12072 2592 12124 2644
rect 16672 2592 16724 2644
rect 20720 2592 20772 2644
rect 21916 2592 21968 2644
rect 3240 2499 3292 2508
rect 3240 2465 3249 2499
rect 3249 2465 3283 2499
rect 3283 2465 3292 2499
rect 3240 2456 3292 2465
rect 3976 2499 4028 2508
rect 3976 2465 3985 2499
rect 3985 2465 4019 2499
rect 4019 2465 4028 2499
rect 3976 2456 4028 2465
rect 8852 2524 8904 2576
rect 4160 2388 4212 2440
rect 4896 2295 4948 2304
rect 4896 2261 4905 2295
rect 4905 2261 4939 2295
rect 4939 2261 4948 2295
rect 4896 2252 4948 2261
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 8392 2456 8444 2508
rect 14096 2456 14148 2508
rect 9588 2388 9640 2440
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 11612 2388 11664 2440
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 13728 2388 13780 2440
rect 14372 2388 14424 2440
rect 16120 2524 16172 2576
rect 22560 2524 22612 2576
rect 17868 2456 17920 2508
rect 16028 2388 16080 2440
rect 19892 2456 19944 2508
rect 19984 2456 20036 2508
rect 23204 2592 23256 2644
rect 25964 2592 26016 2644
rect 27160 2592 27212 2644
rect 28816 2592 28868 2644
rect 34520 2592 34572 2644
rect 36268 2592 36320 2644
rect 36360 2592 36412 2644
rect 38844 2592 38896 2644
rect 41604 2635 41656 2644
rect 41604 2601 41613 2635
rect 41613 2601 41647 2635
rect 41647 2601 41656 2635
rect 41604 2592 41656 2601
rect 47124 2592 47176 2644
rect 49976 2635 50028 2644
rect 49976 2601 49985 2635
rect 49985 2601 50019 2635
rect 50019 2601 50028 2635
rect 49976 2592 50028 2601
rect 72976 2592 73028 2644
rect 74632 2592 74684 2644
rect 76656 2592 76708 2644
rect 23664 2524 23716 2576
rect 5540 2320 5592 2372
rect 6460 2252 6512 2304
rect 11428 2320 11480 2372
rect 12624 2320 12676 2372
rect 13544 2320 13596 2372
rect 17132 2320 17184 2372
rect 17316 2363 17368 2372
rect 17316 2329 17325 2363
rect 17325 2329 17359 2363
rect 17359 2329 17368 2363
rect 17316 2320 17368 2329
rect 11060 2252 11112 2304
rect 12164 2252 12216 2304
rect 12256 2295 12308 2304
rect 12256 2261 12265 2295
rect 12265 2261 12299 2295
rect 12299 2261 12308 2295
rect 12256 2252 12308 2261
rect 14096 2252 14148 2304
rect 17592 2295 17644 2304
rect 17592 2261 17601 2295
rect 17601 2261 17635 2295
rect 17635 2261 17644 2295
rect 17592 2252 17644 2261
rect 18144 2320 18196 2372
rect 19616 2388 19668 2440
rect 19800 2431 19852 2440
rect 19800 2397 19809 2431
rect 19809 2397 19843 2431
rect 19843 2397 19852 2431
rect 19800 2388 19852 2397
rect 21824 2388 21876 2440
rect 22468 2431 22520 2440
rect 22468 2397 22477 2431
rect 22477 2397 22511 2431
rect 22511 2397 22520 2431
rect 22468 2388 22520 2397
rect 22560 2388 22612 2440
rect 23020 2388 23072 2440
rect 24768 2456 24820 2508
rect 26792 2456 26844 2508
rect 30196 2456 30248 2508
rect 28264 2431 28316 2440
rect 28264 2397 28273 2431
rect 28273 2397 28307 2431
rect 28307 2397 28316 2431
rect 28264 2388 28316 2397
rect 30380 2388 30432 2440
rect 33140 2524 33192 2576
rect 33416 2524 33468 2576
rect 32220 2499 32272 2508
rect 32220 2465 32229 2499
rect 32229 2465 32263 2499
rect 32263 2465 32272 2499
rect 32220 2456 32272 2465
rect 34704 2456 34756 2508
rect 31484 2431 31536 2440
rect 31484 2397 31493 2431
rect 31493 2397 31527 2431
rect 31527 2397 31536 2431
rect 31484 2388 31536 2397
rect 25504 2320 25556 2372
rect 25596 2363 25648 2372
rect 25596 2329 25605 2363
rect 25605 2329 25639 2363
rect 25639 2329 25648 2363
rect 25596 2320 25648 2329
rect 26240 2320 26292 2372
rect 28356 2320 28408 2372
rect 33416 2431 33468 2440
rect 33416 2397 33425 2431
rect 33425 2397 33459 2431
rect 33459 2397 33468 2431
rect 33416 2388 33468 2397
rect 35256 2431 35308 2440
rect 35256 2397 35265 2431
rect 35265 2397 35299 2431
rect 35299 2397 35308 2431
rect 35256 2388 35308 2397
rect 35532 2456 35584 2508
rect 36084 2456 36136 2508
rect 39488 2456 39540 2508
rect 39948 2499 40000 2508
rect 39948 2465 39957 2499
rect 39957 2465 39991 2499
rect 39991 2465 40000 2499
rect 39948 2456 40000 2465
rect 40316 2456 40368 2508
rect 34152 2320 34204 2372
rect 36912 2388 36964 2440
rect 38384 2431 38436 2440
rect 38384 2397 38393 2431
rect 38393 2397 38427 2431
rect 38427 2397 38436 2431
rect 38384 2388 38436 2397
rect 39396 2431 39448 2440
rect 39396 2397 39405 2431
rect 39405 2397 39439 2431
rect 39439 2397 39448 2431
rect 39396 2388 39448 2397
rect 41144 2388 41196 2440
rect 41052 2320 41104 2372
rect 41972 2431 42024 2440
rect 41972 2397 41981 2431
rect 41981 2397 42015 2431
rect 42015 2397 42024 2431
rect 41972 2388 42024 2397
rect 48136 2524 48188 2576
rect 49608 2524 49660 2576
rect 46756 2499 46808 2508
rect 46756 2465 46765 2499
rect 46765 2465 46799 2499
rect 46799 2465 46808 2499
rect 46756 2456 46808 2465
rect 49792 2456 49844 2508
rect 50528 2499 50580 2508
rect 50528 2465 50537 2499
rect 50537 2465 50571 2499
rect 50571 2465 50580 2499
rect 50528 2456 50580 2465
rect 52092 2499 52144 2508
rect 52092 2465 52101 2499
rect 52101 2465 52135 2499
rect 52135 2465 52144 2499
rect 52092 2456 52144 2465
rect 54024 2499 54076 2508
rect 54024 2465 54033 2499
rect 54033 2465 54067 2499
rect 54067 2465 54076 2499
rect 54024 2456 54076 2465
rect 45836 2388 45888 2440
rect 47952 2431 48004 2440
rect 47952 2397 47961 2431
rect 47961 2397 47995 2431
rect 47995 2397 48004 2431
rect 47952 2388 48004 2397
rect 48412 2388 48464 2440
rect 49700 2431 49752 2440
rect 49700 2397 49709 2431
rect 49709 2397 49743 2431
rect 49743 2397 49752 2431
rect 49700 2388 49752 2397
rect 52828 2431 52880 2440
rect 52828 2397 52837 2431
rect 52837 2397 52871 2431
rect 52871 2397 52880 2431
rect 52828 2388 52880 2397
rect 55312 2388 55364 2440
rect 55404 2388 55456 2440
rect 58624 2431 58676 2440
rect 58624 2397 58633 2431
rect 58633 2397 58667 2431
rect 58667 2397 58676 2431
rect 58624 2388 58676 2397
rect 21088 2295 21140 2304
rect 21088 2261 21097 2295
rect 21097 2261 21131 2295
rect 21131 2261 21140 2295
rect 21088 2252 21140 2261
rect 22928 2252 22980 2304
rect 24492 2252 24544 2304
rect 33232 2295 33284 2304
rect 33232 2261 33241 2295
rect 33241 2261 33275 2295
rect 33275 2261 33284 2295
rect 33232 2252 33284 2261
rect 36360 2252 36412 2304
rect 38108 2252 38160 2304
rect 41880 2320 41932 2372
rect 57336 2320 57388 2372
rect 61752 2499 61804 2508
rect 61752 2465 61761 2499
rect 61761 2465 61795 2499
rect 61795 2465 61804 2499
rect 61752 2456 61804 2465
rect 65524 2499 65576 2508
rect 65524 2465 65533 2499
rect 65533 2465 65567 2499
rect 65567 2465 65576 2499
rect 65524 2456 65576 2465
rect 67640 2499 67692 2508
rect 67640 2465 67649 2499
rect 67649 2465 67683 2499
rect 67683 2465 67692 2499
rect 67640 2456 67692 2465
rect 69480 2499 69532 2508
rect 69480 2465 69489 2499
rect 69489 2465 69523 2499
rect 69523 2465 69532 2499
rect 69480 2456 69532 2465
rect 70308 2456 70360 2508
rect 62764 2431 62816 2440
rect 62764 2397 62773 2431
rect 62773 2397 62807 2431
rect 62807 2397 62816 2431
rect 62764 2388 62816 2397
rect 63132 2388 63184 2440
rect 66260 2431 66312 2440
rect 66260 2397 66269 2431
rect 66269 2397 66303 2431
rect 66303 2397 66312 2431
rect 66260 2388 66312 2397
rect 68284 2431 68336 2440
rect 68284 2397 68293 2431
rect 68293 2397 68327 2431
rect 68327 2397 68336 2431
rect 68284 2388 68336 2397
rect 70492 2431 70544 2440
rect 70492 2397 70501 2431
rect 70501 2397 70535 2431
rect 70535 2397 70544 2431
rect 70492 2388 70544 2397
rect 72608 2499 72660 2508
rect 72608 2465 72617 2499
rect 72617 2465 72651 2499
rect 72651 2465 72660 2499
rect 72608 2456 72660 2465
rect 72792 2456 72844 2508
rect 75460 2456 75512 2508
rect 73252 2388 73304 2440
rect 76196 2431 76248 2440
rect 76196 2397 76205 2431
rect 76205 2397 76239 2431
rect 76239 2397 76248 2431
rect 76196 2388 76248 2397
rect 41328 2252 41380 2304
rect 47584 2252 47636 2304
rect 5794 2150 5846 2202
rect 5858 2150 5910 2202
rect 5922 2150 5974 2202
rect 5986 2150 6038 2202
rect 6050 2150 6102 2202
rect 36514 2150 36566 2202
rect 36578 2150 36630 2202
rect 36642 2150 36694 2202
rect 36706 2150 36758 2202
rect 36770 2150 36822 2202
rect 67234 2150 67286 2202
rect 67298 2150 67350 2202
rect 67362 2150 67414 2202
rect 67426 2150 67478 2202
rect 67490 2150 67542 2202
rect 12256 2048 12308 2100
rect 17224 2048 17276 2100
rect 20536 2048 20588 2100
rect 30932 2048 30984 2100
rect 38108 2048 38160 2100
rect 47952 2048 48004 2100
rect 10232 1980 10284 2032
rect 12624 1980 12676 2032
rect 18972 1980 19024 2032
rect 32404 1980 32456 2032
rect 33416 1980 33468 2032
rect 40592 1980 40644 2032
rect 9864 1912 9916 1964
rect 17592 1912 17644 1964
rect 27528 1912 27580 1964
rect 38384 1912 38436 1964
rect 12072 1844 12124 1896
rect 17408 1844 17460 1896
rect 21824 1844 21876 1896
rect 5724 1776 5776 1828
rect 13912 1776 13964 1828
rect 18512 1776 18564 1828
rect 31944 1776 31996 1828
rect 33232 1844 33284 1896
rect 38292 1844 38344 1896
rect 38200 1776 38252 1828
rect 23940 1708 23992 1760
rect 40776 1708 40828 1760
rect 15660 1640 15712 1692
rect 25596 1640 25648 1692
rect 18880 1572 18932 1624
rect 31484 1572 31536 1624
rect 8024 1368 8076 1420
rect 9680 1368 9732 1420
rect 14280 1368 14332 1420
rect 21272 1368 21324 1420
rect 22192 1368 22244 1420
rect 23204 1368 23256 1420
rect 10048 1300 10100 1352
rect 16120 1300 16172 1352
rect 17040 1300 17092 1352
rect 19340 1300 19392 1352
rect 13268 1232 13320 1284
rect 18052 1232 18104 1284
rect 16948 1164 17000 1216
rect 25780 1164 25832 1216
rect 21180 280 21232 332
rect 29552 280 29604 332
rect 10692 212 10744 264
rect 21824 212 21876 264
rect 21548 144 21600 196
rect 33416 144 33468 196
rect 9588 76 9640 128
rect 23756 76 23808 128
<< metal2 >>
rect 2226 39200 2282 40000
rect 4066 39200 4122 40000
rect 5906 39200 5962 40000
rect 7746 39200 7802 40000
rect 9586 39200 9642 40000
rect 11426 39200 11482 40000
rect 13266 39200 13322 40000
rect 15106 39200 15162 40000
rect 16946 39200 17002 40000
rect 18786 39200 18842 40000
rect 20626 39200 20682 40000
rect 22466 39200 22522 40000
rect 24306 39200 24362 40000
rect 26146 39200 26202 40000
rect 27986 39200 28042 40000
rect 29826 39200 29882 40000
rect 31666 39200 31722 40000
rect 33506 39200 33562 40000
rect 35346 39200 35402 40000
rect 37186 39200 37242 40000
rect 39026 39200 39082 40000
rect 40866 39200 40922 40000
rect 42706 39200 42762 40000
rect 44546 39200 44602 40000
rect 46386 39200 46442 40000
rect 48226 39200 48282 40000
rect 50066 39200 50122 40000
rect 51906 39200 51962 40000
rect 53746 39200 53802 40000
rect 55586 39200 55642 40000
rect 57426 39200 57482 40000
rect 59266 39200 59322 40000
rect 2240 37330 2268 39200
rect 2228 37324 2280 37330
rect 2228 37266 2280 37272
rect 3516 37256 3568 37262
rect 3516 37198 3568 37204
rect 3528 24138 3556 37198
rect 4080 36854 4108 39200
rect 5134 37564 5442 37573
rect 5134 37562 5140 37564
rect 5196 37562 5220 37564
rect 5276 37562 5300 37564
rect 5356 37562 5380 37564
rect 5436 37562 5442 37564
rect 5196 37510 5198 37562
rect 5378 37510 5380 37562
rect 5134 37508 5140 37510
rect 5196 37508 5220 37510
rect 5276 37508 5300 37510
rect 5356 37508 5380 37510
rect 5436 37508 5442 37510
rect 5134 37499 5442 37508
rect 5920 37262 5948 39200
rect 7760 37618 7788 39200
rect 7760 37590 7972 37618
rect 7944 37262 7972 37590
rect 5908 37256 5960 37262
rect 5908 37198 5960 37204
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 7748 37256 7800 37262
rect 7748 37198 7800 37204
rect 7932 37256 7984 37262
rect 7932 37198 7984 37204
rect 5794 37020 6102 37029
rect 5794 37018 5800 37020
rect 5856 37018 5880 37020
rect 5936 37018 5960 37020
rect 6016 37018 6040 37020
rect 6096 37018 6102 37020
rect 5856 36966 5858 37018
rect 6038 36966 6040 37018
rect 5794 36964 5800 36966
rect 5856 36964 5880 36966
rect 5936 36964 5960 36966
rect 6016 36964 6040 36966
rect 6096 36964 6102 36966
rect 5794 36955 6102 36964
rect 4068 36848 4120 36854
rect 4068 36790 4120 36796
rect 5134 36476 5442 36485
rect 5134 36474 5140 36476
rect 5196 36474 5220 36476
rect 5276 36474 5300 36476
rect 5356 36474 5380 36476
rect 5436 36474 5442 36476
rect 5196 36422 5198 36474
rect 5378 36422 5380 36474
rect 5134 36420 5140 36422
rect 5196 36420 5220 36422
rect 5276 36420 5300 36422
rect 5356 36420 5380 36422
rect 5436 36420 5442 36422
rect 5134 36411 5442 36420
rect 5794 35932 6102 35941
rect 5794 35930 5800 35932
rect 5856 35930 5880 35932
rect 5936 35930 5960 35932
rect 6016 35930 6040 35932
rect 6096 35930 6102 35932
rect 5856 35878 5858 35930
rect 6038 35878 6040 35930
rect 5794 35876 5800 35878
rect 5856 35876 5880 35878
rect 5936 35876 5960 35878
rect 6016 35876 6040 35878
rect 6096 35876 6102 35878
rect 5794 35867 6102 35876
rect 5134 35388 5442 35397
rect 5134 35386 5140 35388
rect 5196 35386 5220 35388
rect 5276 35386 5300 35388
rect 5356 35386 5380 35388
rect 5436 35386 5442 35388
rect 5196 35334 5198 35386
rect 5378 35334 5380 35386
rect 5134 35332 5140 35334
rect 5196 35332 5220 35334
rect 5276 35332 5300 35334
rect 5356 35332 5380 35334
rect 5436 35332 5442 35334
rect 5134 35323 5442 35332
rect 5794 34844 6102 34853
rect 5794 34842 5800 34844
rect 5856 34842 5880 34844
rect 5936 34842 5960 34844
rect 6016 34842 6040 34844
rect 6096 34842 6102 34844
rect 5856 34790 5858 34842
rect 6038 34790 6040 34842
rect 5794 34788 5800 34790
rect 5856 34788 5880 34790
rect 5936 34788 5960 34790
rect 6016 34788 6040 34790
rect 6096 34788 6102 34790
rect 5794 34779 6102 34788
rect 5134 34300 5442 34309
rect 5134 34298 5140 34300
rect 5196 34298 5220 34300
rect 5276 34298 5300 34300
rect 5356 34298 5380 34300
rect 5436 34298 5442 34300
rect 5196 34246 5198 34298
rect 5378 34246 5380 34298
rect 5134 34244 5140 34246
rect 5196 34244 5220 34246
rect 5276 34244 5300 34246
rect 5356 34244 5380 34246
rect 5436 34244 5442 34246
rect 5134 34235 5442 34244
rect 5794 33756 6102 33765
rect 5794 33754 5800 33756
rect 5856 33754 5880 33756
rect 5936 33754 5960 33756
rect 6016 33754 6040 33756
rect 6096 33754 6102 33756
rect 5856 33702 5858 33754
rect 6038 33702 6040 33754
rect 5794 33700 5800 33702
rect 5856 33700 5880 33702
rect 5936 33700 5960 33702
rect 6016 33700 6040 33702
rect 6096 33700 6102 33702
rect 5794 33691 6102 33700
rect 5134 33212 5442 33221
rect 5134 33210 5140 33212
rect 5196 33210 5220 33212
rect 5276 33210 5300 33212
rect 5356 33210 5380 33212
rect 5436 33210 5442 33212
rect 5196 33158 5198 33210
rect 5378 33158 5380 33210
rect 5134 33156 5140 33158
rect 5196 33156 5220 33158
rect 5276 33156 5300 33158
rect 5356 33156 5380 33158
rect 5436 33156 5442 33158
rect 5134 33147 5442 33156
rect 5794 32668 6102 32677
rect 5794 32666 5800 32668
rect 5856 32666 5880 32668
rect 5936 32666 5960 32668
rect 6016 32666 6040 32668
rect 6096 32666 6102 32668
rect 5856 32614 5858 32666
rect 6038 32614 6040 32666
rect 5794 32612 5800 32614
rect 5856 32612 5880 32614
rect 5936 32612 5960 32614
rect 6016 32612 6040 32614
rect 6096 32612 6102 32614
rect 5794 32603 6102 32612
rect 7116 32473 7144 37198
rect 7760 36922 7788 37198
rect 7748 36916 7800 36922
rect 7748 36858 7800 36864
rect 9600 36854 9628 39200
rect 11440 37262 11468 39200
rect 13280 37330 13308 39200
rect 15120 37346 15148 39200
rect 13268 37324 13320 37330
rect 13268 37266 13320 37272
rect 15028 37318 15148 37346
rect 11428 37256 11480 37262
rect 11428 37198 11480 37204
rect 11888 37256 11940 37262
rect 11888 37198 11940 37204
rect 14556 37256 14608 37262
rect 14556 37198 14608 37204
rect 11900 36922 11928 37198
rect 11888 36916 11940 36922
rect 11888 36858 11940 36864
rect 9588 36848 9640 36854
rect 9588 36790 9640 36796
rect 10968 36780 11020 36786
rect 10968 36722 11020 36728
rect 11796 36780 11848 36786
rect 11796 36722 11848 36728
rect 7102 32464 7158 32473
rect 7102 32399 7158 32408
rect 5134 32124 5442 32133
rect 5134 32122 5140 32124
rect 5196 32122 5220 32124
rect 5276 32122 5300 32124
rect 5356 32122 5380 32124
rect 5436 32122 5442 32124
rect 5196 32070 5198 32122
rect 5378 32070 5380 32122
rect 5134 32068 5140 32070
rect 5196 32068 5220 32070
rect 5276 32068 5300 32070
rect 5356 32068 5380 32070
rect 5436 32068 5442 32070
rect 5134 32059 5442 32068
rect 5794 31580 6102 31589
rect 5794 31578 5800 31580
rect 5856 31578 5880 31580
rect 5936 31578 5960 31580
rect 6016 31578 6040 31580
rect 6096 31578 6102 31580
rect 5856 31526 5858 31578
rect 6038 31526 6040 31578
rect 5794 31524 5800 31526
rect 5856 31524 5880 31526
rect 5936 31524 5960 31526
rect 6016 31524 6040 31526
rect 6096 31524 6102 31526
rect 5794 31515 6102 31524
rect 5134 31036 5442 31045
rect 5134 31034 5140 31036
rect 5196 31034 5220 31036
rect 5276 31034 5300 31036
rect 5356 31034 5380 31036
rect 5436 31034 5442 31036
rect 5196 30982 5198 31034
rect 5378 30982 5380 31034
rect 5134 30980 5140 30982
rect 5196 30980 5220 30982
rect 5276 30980 5300 30982
rect 5356 30980 5380 30982
rect 5436 30980 5442 30982
rect 5134 30971 5442 30980
rect 5794 30492 6102 30501
rect 5794 30490 5800 30492
rect 5856 30490 5880 30492
rect 5936 30490 5960 30492
rect 6016 30490 6040 30492
rect 6096 30490 6102 30492
rect 5856 30438 5858 30490
rect 6038 30438 6040 30490
rect 5794 30436 5800 30438
rect 5856 30436 5880 30438
rect 5936 30436 5960 30438
rect 6016 30436 6040 30438
rect 6096 30436 6102 30438
rect 5794 30427 6102 30436
rect 5134 29948 5442 29957
rect 5134 29946 5140 29948
rect 5196 29946 5220 29948
rect 5276 29946 5300 29948
rect 5356 29946 5380 29948
rect 5436 29946 5442 29948
rect 5196 29894 5198 29946
rect 5378 29894 5380 29946
rect 5134 29892 5140 29894
rect 5196 29892 5220 29894
rect 5276 29892 5300 29894
rect 5356 29892 5380 29894
rect 5436 29892 5442 29894
rect 5134 29883 5442 29892
rect 10980 29617 11008 36722
rect 11808 36650 11836 36722
rect 11796 36644 11848 36650
rect 11796 36586 11848 36592
rect 10966 29608 11022 29617
rect 10966 29543 11022 29552
rect 5794 29404 6102 29413
rect 5794 29402 5800 29404
rect 5856 29402 5880 29404
rect 5936 29402 5960 29404
rect 6016 29402 6040 29404
rect 6096 29402 6102 29404
rect 5856 29350 5858 29402
rect 6038 29350 6040 29402
rect 5794 29348 5800 29350
rect 5856 29348 5880 29350
rect 5936 29348 5960 29350
rect 6016 29348 6040 29350
rect 6096 29348 6102 29350
rect 5794 29339 6102 29348
rect 5134 28860 5442 28869
rect 5134 28858 5140 28860
rect 5196 28858 5220 28860
rect 5276 28858 5300 28860
rect 5356 28858 5380 28860
rect 5436 28858 5442 28860
rect 5196 28806 5198 28858
rect 5378 28806 5380 28858
rect 5134 28804 5140 28806
rect 5196 28804 5220 28806
rect 5276 28804 5300 28806
rect 5356 28804 5380 28806
rect 5436 28804 5442 28806
rect 5134 28795 5442 28804
rect 5794 28316 6102 28325
rect 5794 28314 5800 28316
rect 5856 28314 5880 28316
rect 5936 28314 5960 28316
rect 6016 28314 6040 28316
rect 6096 28314 6102 28316
rect 5856 28262 5858 28314
rect 6038 28262 6040 28314
rect 5794 28260 5800 28262
rect 5856 28260 5880 28262
rect 5936 28260 5960 28262
rect 6016 28260 6040 28262
rect 6096 28260 6102 28262
rect 5794 28251 6102 28260
rect 5134 27772 5442 27781
rect 5134 27770 5140 27772
rect 5196 27770 5220 27772
rect 5276 27770 5300 27772
rect 5356 27770 5380 27772
rect 5436 27770 5442 27772
rect 5196 27718 5198 27770
rect 5378 27718 5380 27770
rect 5134 27716 5140 27718
rect 5196 27716 5220 27718
rect 5276 27716 5300 27718
rect 5356 27716 5380 27718
rect 5436 27716 5442 27718
rect 5134 27707 5442 27716
rect 5794 27228 6102 27237
rect 5794 27226 5800 27228
rect 5856 27226 5880 27228
rect 5936 27226 5960 27228
rect 6016 27226 6040 27228
rect 6096 27226 6102 27228
rect 5856 27174 5858 27226
rect 6038 27174 6040 27226
rect 5794 27172 5800 27174
rect 5856 27172 5880 27174
rect 5936 27172 5960 27174
rect 6016 27172 6040 27174
rect 6096 27172 6102 27174
rect 5794 27163 6102 27172
rect 5134 26684 5442 26693
rect 5134 26682 5140 26684
rect 5196 26682 5220 26684
rect 5276 26682 5300 26684
rect 5356 26682 5380 26684
rect 5436 26682 5442 26684
rect 5196 26630 5198 26682
rect 5378 26630 5380 26682
rect 5134 26628 5140 26630
rect 5196 26628 5220 26630
rect 5276 26628 5300 26630
rect 5356 26628 5380 26630
rect 5436 26628 5442 26630
rect 5134 26619 5442 26628
rect 11808 26234 11836 36586
rect 14568 36553 14596 37198
rect 15028 37194 15056 37318
rect 15108 37256 15160 37262
rect 15108 37198 15160 37204
rect 15016 37188 15068 37194
rect 15016 37130 15068 37136
rect 15120 36922 15148 37198
rect 15108 36916 15160 36922
rect 15108 36858 15160 36864
rect 16960 36854 16988 39200
rect 18800 37262 18828 39200
rect 20640 37262 20668 39200
rect 22480 37346 22508 39200
rect 22480 37318 22600 37346
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 18788 37256 18840 37262
rect 18788 37198 18840 37204
rect 20628 37256 20680 37262
rect 20628 37198 20680 37204
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 18708 36922 18736 37198
rect 18696 36916 18748 36922
rect 18696 36858 18748 36864
rect 16948 36848 17000 36854
rect 16948 36790 17000 36796
rect 18788 36780 18840 36786
rect 18788 36722 18840 36728
rect 14554 36544 14610 36553
rect 14554 36479 14610 36488
rect 18800 26994 18828 36722
rect 18788 26988 18840 26994
rect 18788 26930 18840 26936
rect 11716 26206 11836 26234
rect 5794 26140 6102 26149
rect 5794 26138 5800 26140
rect 5856 26138 5880 26140
rect 5936 26138 5960 26140
rect 6016 26138 6040 26140
rect 6096 26138 6102 26140
rect 5856 26086 5858 26138
rect 6038 26086 6040 26138
rect 5794 26084 5800 26086
rect 5856 26084 5880 26086
rect 5936 26084 5960 26086
rect 6016 26084 6040 26086
rect 6096 26084 6102 26086
rect 5794 26075 6102 26084
rect 5134 25596 5442 25605
rect 5134 25594 5140 25596
rect 5196 25594 5220 25596
rect 5276 25594 5300 25596
rect 5356 25594 5380 25596
rect 5436 25594 5442 25596
rect 5196 25542 5198 25594
rect 5378 25542 5380 25594
rect 5134 25540 5140 25542
rect 5196 25540 5220 25542
rect 5276 25540 5300 25542
rect 5356 25540 5380 25542
rect 5436 25540 5442 25542
rect 5134 25531 5442 25540
rect 5794 25052 6102 25061
rect 5794 25050 5800 25052
rect 5856 25050 5880 25052
rect 5936 25050 5960 25052
rect 6016 25050 6040 25052
rect 6096 25050 6102 25052
rect 5856 24998 5858 25050
rect 6038 24998 6040 25050
rect 5794 24996 5800 24998
rect 5856 24996 5880 24998
rect 5936 24996 5960 24998
rect 6016 24996 6040 24998
rect 6096 24996 6102 24998
rect 5794 24987 6102 24996
rect 5134 24508 5442 24517
rect 5134 24506 5140 24508
rect 5196 24506 5220 24508
rect 5276 24506 5300 24508
rect 5356 24506 5380 24508
rect 5436 24506 5442 24508
rect 5196 24454 5198 24506
rect 5378 24454 5380 24506
rect 5134 24452 5140 24454
rect 5196 24452 5220 24454
rect 5276 24452 5300 24454
rect 5356 24452 5380 24454
rect 5436 24452 5442 24454
rect 5134 24443 5442 24452
rect 3516 24132 3568 24138
rect 3516 24074 3568 24080
rect 5794 23964 6102 23973
rect 5794 23962 5800 23964
rect 5856 23962 5880 23964
rect 5936 23962 5960 23964
rect 6016 23962 6040 23964
rect 6096 23962 6102 23964
rect 5856 23910 5858 23962
rect 6038 23910 6040 23962
rect 5794 23908 5800 23910
rect 5856 23908 5880 23910
rect 5936 23908 5960 23910
rect 6016 23908 6040 23910
rect 6096 23908 6102 23910
rect 5794 23899 6102 23908
rect 5134 23420 5442 23429
rect 5134 23418 5140 23420
rect 5196 23418 5220 23420
rect 5276 23418 5300 23420
rect 5356 23418 5380 23420
rect 5436 23418 5442 23420
rect 5196 23366 5198 23418
rect 5378 23366 5380 23418
rect 5134 23364 5140 23366
rect 5196 23364 5220 23366
rect 5276 23364 5300 23366
rect 5356 23364 5380 23366
rect 5436 23364 5442 23366
rect 5134 23355 5442 23364
rect 5794 22876 6102 22885
rect 5794 22874 5800 22876
rect 5856 22874 5880 22876
rect 5936 22874 5960 22876
rect 6016 22874 6040 22876
rect 6096 22874 6102 22876
rect 5856 22822 5858 22874
rect 6038 22822 6040 22874
rect 5794 22820 5800 22822
rect 5856 22820 5880 22822
rect 5936 22820 5960 22822
rect 6016 22820 6040 22822
rect 6096 22820 6102 22822
rect 5794 22811 6102 22820
rect 5134 22332 5442 22341
rect 5134 22330 5140 22332
rect 5196 22330 5220 22332
rect 5276 22330 5300 22332
rect 5356 22330 5380 22332
rect 5436 22330 5442 22332
rect 5196 22278 5198 22330
rect 5378 22278 5380 22330
rect 5134 22276 5140 22278
rect 5196 22276 5220 22278
rect 5276 22276 5300 22278
rect 5356 22276 5380 22278
rect 5436 22276 5442 22278
rect 5134 22267 5442 22276
rect 5794 21788 6102 21797
rect 5794 21786 5800 21788
rect 5856 21786 5880 21788
rect 5936 21786 5960 21788
rect 6016 21786 6040 21788
rect 6096 21786 6102 21788
rect 5856 21734 5858 21786
rect 6038 21734 6040 21786
rect 5794 21732 5800 21734
rect 5856 21732 5880 21734
rect 5936 21732 5960 21734
rect 6016 21732 6040 21734
rect 6096 21732 6102 21734
rect 5794 21723 6102 21732
rect 5134 21244 5442 21253
rect 5134 21242 5140 21244
rect 5196 21242 5220 21244
rect 5276 21242 5300 21244
rect 5356 21242 5380 21244
rect 5436 21242 5442 21244
rect 5196 21190 5198 21242
rect 5378 21190 5380 21242
rect 5134 21188 5140 21190
rect 5196 21188 5220 21190
rect 5276 21188 5300 21190
rect 5356 21188 5380 21190
rect 5436 21188 5442 21190
rect 5134 21179 5442 21188
rect 5794 20700 6102 20709
rect 5794 20698 5800 20700
rect 5856 20698 5880 20700
rect 5936 20698 5960 20700
rect 6016 20698 6040 20700
rect 6096 20698 6102 20700
rect 5856 20646 5858 20698
rect 6038 20646 6040 20698
rect 5794 20644 5800 20646
rect 5856 20644 5880 20646
rect 5936 20644 5960 20646
rect 6016 20644 6040 20646
rect 6096 20644 6102 20646
rect 5794 20635 6102 20644
rect 5134 20156 5442 20165
rect 5134 20154 5140 20156
rect 5196 20154 5220 20156
rect 5276 20154 5300 20156
rect 5356 20154 5380 20156
rect 5436 20154 5442 20156
rect 5196 20102 5198 20154
rect 5378 20102 5380 20154
rect 5134 20100 5140 20102
rect 5196 20100 5220 20102
rect 5276 20100 5300 20102
rect 5356 20100 5380 20102
rect 5436 20100 5442 20102
rect 5134 20091 5442 20100
rect 5794 19612 6102 19621
rect 5794 19610 5800 19612
rect 5856 19610 5880 19612
rect 5936 19610 5960 19612
rect 6016 19610 6040 19612
rect 6096 19610 6102 19612
rect 5856 19558 5858 19610
rect 6038 19558 6040 19610
rect 5794 19556 5800 19558
rect 5856 19556 5880 19558
rect 5936 19556 5960 19558
rect 6016 19556 6040 19558
rect 6096 19556 6102 19558
rect 5794 19547 6102 19556
rect 5134 19068 5442 19077
rect 5134 19066 5140 19068
rect 5196 19066 5220 19068
rect 5276 19066 5300 19068
rect 5356 19066 5380 19068
rect 5436 19066 5442 19068
rect 5196 19014 5198 19066
rect 5378 19014 5380 19066
rect 5134 19012 5140 19014
rect 5196 19012 5220 19014
rect 5276 19012 5300 19014
rect 5356 19012 5380 19014
rect 5436 19012 5442 19014
rect 5134 19003 5442 19012
rect 5794 18524 6102 18533
rect 5794 18522 5800 18524
rect 5856 18522 5880 18524
rect 5936 18522 5960 18524
rect 6016 18522 6040 18524
rect 6096 18522 6102 18524
rect 5856 18470 5858 18522
rect 6038 18470 6040 18522
rect 5794 18468 5800 18470
rect 5856 18468 5880 18470
rect 5936 18468 5960 18470
rect 6016 18468 6040 18470
rect 6096 18468 6102 18470
rect 5794 18459 6102 18468
rect 5134 17980 5442 17989
rect 5134 17978 5140 17980
rect 5196 17978 5220 17980
rect 5276 17978 5300 17980
rect 5356 17978 5380 17980
rect 5436 17978 5442 17980
rect 5196 17926 5198 17978
rect 5378 17926 5380 17978
rect 5134 17924 5140 17926
rect 5196 17924 5220 17926
rect 5276 17924 5300 17926
rect 5356 17924 5380 17926
rect 5436 17924 5442 17926
rect 5134 17915 5442 17924
rect 5794 17436 6102 17445
rect 5794 17434 5800 17436
rect 5856 17434 5880 17436
rect 5936 17434 5960 17436
rect 6016 17434 6040 17436
rect 6096 17434 6102 17436
rect 5856 17382 5858 17434
rect 6038 17382 6040 17434
rect 5794 17380 5800 17382
rect 5856 17380 5880 17382
rect 5936 17380 5960 17382
rect 6016 17380 6040 17382
rect 6096 17380 6102 17382
rect 5794 17371 6102 17380
rect 5134 16892 5442 16901
rect 5134 16890 5140 16892
rect 5196 16890 5220 16892
rect 5276 16890 5300 16892
rect 5356 16890 5380 16892
rect 5436 16890 5442 16892
rect 5196 16838 5198 16890
rect 5378 16838 5380 16890
rect 5134 16836 5140 16838
rect 5196 16836 5220 16838
rect 5276 16836 5300 16838
rect 5356 16836 5380 16838
rect 5436 16836 5442 16838
rect 5134 16827 5442 16836
rect 5794 16348 6102 16357
rect 5794 16346 5800 16348
rect 5856 16346 5880 16348
rect 5936 16346 5960 16348
rect 6016 16346 6040 16348
rect 6096 16346 6102 16348
rect 5856 16294 5858 16346
rect 6038 16294 6040 16346
rect 5794 16292 5800 16294
rect 5856 16292 5880 16294
rect 5936 16292 5960 16294
rect 6016 16292 6040 16294
rect 6096 16292 6102 16294
rect 5794 16283 6102 16292
rect 5134 15804 5442 15813
rect 5134 15802 5140 15804
rect 5196 15802 5220 15804
rect 5276 15802 5300 15804
rect 5356 15802 5380 15804
rect 5436 15802 5442 15804
rect 5196 15750 5198 15802
rect 5378 15750 5380 15802
rect 5134 15748 5140 15750
rect 5196 15748 5220 15750
rect 5276 15748 5300 15750
rect 5356 15748 5380 15750
rect 5436 15748 5442 15750
rect 5134 15739 5442 15748
rect 5794 15260 6102 15269
rect 5794 15258 5800 15260
rect 5856 15258 5880 15260
rect 5936 15258 5960 15260
rect 6016 15258 6040 15260
rect 6096 15258 6102 15260
rect 5856 15206 5858 15258
rect 6038 15206 6040 15258
rect 5794 15204 5800 15206
rect 5856 15204 5880 15206
rect 5936 15204 5960 15206
rect 6016 15204 6040 15206
rect 6096 15204 6102 15206
rect 5794 15195 6102 15204
rect 5134 14716 5442 14725
rect 5134 14714 5140 14716
rect 5196 14714 5220 14716
rect 5276 14714 5300 14716
rect 5356 14714 5380 14716
rect 5436 14714 5442 14716
rect 5196 14662 5198 14714
rect 5378 14662 5380 14714
rect 5134 14660 5140 14662
rect 5196 14660 5220 14662
rect 5276 14660 5300 14662
rect 5356 14660 5380 14662
rect 5436 14660 5442 14662
rect 5134 14651 5442 14660
rect 5794 14172 6102 14181
rect 5794 14170 5800 14172
rect 5856 14170 5880 14172
rect 5936 14170 5960 14172
rect 6016 14170 6040 14172
rect 6096 14170 6102 14172
rect 5856 14118 5858 14170
rect 6038 14118 6040 14170
rect 5794 14116 5800 14118
rect 5856 14116 5880 14118
rect 5936 14116 5960 14118
rect 6016 14116 6040 14118
rect 6096 14116 6102 14118
rect 5794 14107 6102 14116
rect 5134 13628 5442 13637
rect 5134 13626 5140 13628
rect 5196 13626 5220 13628
rect 5276 13626 5300 13628
rect 5356 13626 5380 13628
rect 5436 13626 5442 13628
rect 5196 13574 5198 13626
rect 5378 13574 5380 13626
rect 5134 13572 5140 13574
rect 5196 13572 5220 13574
rect 5276 13572 5300 13574
rect 5356 13572 5380 13574
rect 5436 13572 5442 13574
rect 5134 13563 5442 13572
rect 5794 13084 6102 13093
rect 5794 13082 5800 13084
rect 5856 13082 5880 13084
rect 5936 13082 5960 13084
rect 6016 13082 6040 13084
rect 6096 13082 6102 13084
rect 5856 13030 5858 13082
rect 6038 13030 6040 13082
rect 5794 13028 5800 13030
rect 5856 13028 5880 13030
rect 5936 13028 5960 13030
rect 6016 13028 6040 13030
rect 6096 13028 6102 13030
rect 5794 13019 6102 13028
rect 5134 12540 5442 12549
rect 5134 12538 5140 12540
rect 5196 12538 5220 12540
rect 5276 12538 5300 12540
rect 5356 12538 5380 12540
rect 5436 12538 5442 12540
rect 5196 12486 5198 12538
rect 5378 12486 5380 12538
rect 5134 12484 5140 12486
rect 5196 12484 5220 12486
rect 5276 12484 5300 12486
rect 5356 12484 5380 12486
rect 5436 12484 5442 12486
rect 5134 12475 5442 12484
rect 5794 11996 6102 12005
rect 5794 11994 5800 11996
rect 5856 11994 5880 11996
rect 5936 11994 5960 11996
rect 6016 11994 6040 11996
rect 6096 11994 6102 11996
rect 5856 11942 5858 11994
rect 6038 11942 6040 11994
rect 5794 11940 5800 11942
rect 5856 11940 5880 11942
rect 5936 11940 5960 11942
rect 6016 11940 6040 11942
rect 6096 11940 6102 11942
rect 5794 11931 6102 11940
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 5134 11452 5442 11461
rect 5134 11450 5140 11452
rect 5196 11450 5220 11452
rect 5276 11450 5300 11452
rect 5356 11450 5380 11452
rect 5436 11450 5442 11452
rect 5196 11398 5198 11450
rect 5378 11398 5380 11450
rect 5134 11396 5140 11398
rect 5196 11396 5220 11398
rect 5276 11396 5300 11398
rect 5356 11396 5380 11398
rect 5436 11396 5442 11398
rect 5134 11387 5442 11396
rect 5794 10908 6102 10917
rect 5794 10906 5800 10908
rect 5856 10906 5880 10908
rect 5936 10906 5960 10908
rect 6016 10906 6040 10908
rect 6096 10906 6102 10908
rect 5856 10854 5858 10906
rect 6038 10854 6040 10906
rect 5794 10852 5800 10854
rect 5856 10852 5880 10854
rect 5936 10852 5960 10854
rect 6016 10852 6040 10854
rect 6096 10852 6102 10854
rect 5794 10843 6102 10852
rect 5134 10364 5442 10373
rect 5134 10362 5140 10364
rect 5196 10362 5220 10364
rect 5276 10362 5300 10364
rect 5356 10362 5380 10364
rect 5436 10362 5442 10364
rect 5196 10310 5198 10362
rect 5378 10310 5380 10362
rect 5134 10308 5140 10310
rect 5196 10308 5220 10310
rect 5276 10308 5300 10310
rect 5356 10308 5380 10310
rect 5436 10308 5442 10310
rect 5134 10299 5442 10308
rect 5794 9820 6102 9829
rect 5794 9818 5800 9820
rect 5856 9818 5880 9820
rect 5936 9818 5960 9820
rect 6016 9818 6040 9820
rect 6096 9818 6102 9820
rect 5856 9766 5858 9818
rect 6038 9766 6040 9818
rect 5794 9764 5800 9766
rect 5856 9764 5880 9766
rect 5936 9764 5960 9766
rect 6016 9764 6040 9766
rect 6096 9764 6102 9766
rect 5794 9755 6102 9764
rect 5134 9276 5442 9285
rect 5134 9274 5140 9276
rect 5196 9274 5220 9276
rect 5276 9274 5300 9276
rect 5356 9274 5380 9276
rect 5436 9274 5442 9276
rect 5196 9222 5198 9274
rect 5378 9222 5380 9274
rect 5134 9220 5140 9222
rect 5196 9220 5220 9222
rect 5276 9220 5300 9222
rect 5356 9220 5380 9222
rect 5436 9220 5442 9222
rect 5134 9211 5442 9220
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 2514 3280 8774
rect 5794 8732 6102 8741
rect 5794 8730 5800 8732
rect 5856 8730 5880 8732
rect 5936 8730 5960 8732
rect 6016 8730 6040 8732
rect 6096 8730 6102 8732
rect 5856 8678 5858 8730
rect 6038 8678 6040 8730
rect 5794 8676 5800 8678
rect 5856 8676 5880 8678
rect 5936 8676 5960 8678
rect 6016 8676 6040 8678
rect 6096 8676 6102 8678
rect 5794 8667 6102 8676
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3804 3194 3832 4014
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3896 2650 3924 5510
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3988 2514 4016 8298
rect 5134 8188 5442 8197
rect 5134 8186 5140 8188
rect 5196 8186 5220 8188
rect 5276 8186 5300 8188
rect 5356 8186 5380 8188
rect 5436 8186 5442 8188
rect 5196 8134 5198 8186
rect 5378 8134 5380 8186
rect 5134 8132 5140 8134
rect 5196 8132 5220 8134
rect 5276 8132 5300 8134
rect 5356 8132 5380 8134
rect 5436 8132 5442 8134
rect 5134 8123 5442 8132
rect 5794 7644 6102 7653
rect 5794 7642 5800 7644
rect 5856 7642 5880 7644
rect 5936 7642 5960 7644
rect 6016 7642 6040 7644
rect 6096 7642 6102 7644
rect 5856 7590 5858 7642
rect 6038 7590 6040 7642
rect 5794 7588 5800 7590
rect 5856 7588 5880 7590
rect 5936 7588 5960 7590
rect 6016 7588 6040 7590
rect 6096 7588 6102 7590
rect 5794 7579 6102 7588
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 5134 7100 5442 7109
rect 5134 7098 5140 7100
rect 5196 7098 5220 7100
rect 5276 7098 5300 7100
rect 5356 7098 5380 7100
rect 5436 7098 5442 7100
rect 5196 7046 5198 7098
rect 5378 7046 5380 7098
rect 5134 7044 5140 7046
rect 5196 7044 5220 7046
rect 5276 7044 5300 7046
rect 5356 7044 5380 7046
rect 5436 7044 5442 7046
rect 5134 7035 5442 7044
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 5794 6556 6102 6565
rect 5794 6554 5800 6556
rect 5856 6554 5880 6556
rect 5936 6554 5960 6556
rect 6016 6554 6040 6556
rect 6096 6554 6102 6556
rect 5856 6502 5858 6554
rect 6038 6502 6040 6554
rect 5794 6500 5800 6502
rect 5856 6500 5880 6502
rect 5936 6500 5960 6502
rect 6016 6500 6040 6502
rect 6096 6500 6102 6502
rect 5794 6491 6102 6500
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5134 6012 5442 6021
rect 5134 6010 5140 6012
rect 5196 6010 5220 6012
rect 5276 6010 5300 6012
rect 5356 6010 5380 6012
rect 5436 6010 5442 6012
rect 5196 5958 5198 6010
rect 5378 5958 5380 6010
rect 5134 5956 5140 5958
rect 5196 5956 5220 5958
rect 5276 5956 5300 5958
rect 5356 5956 5380 5958
rect 5436 5956 5442 5958
rect 5134 5947 5442 5956
rect 5134 4924 5442 4933
rect 5134 4922 5140 4924
rect 5196 4922 5220 4924
rect 5276 4922 5300 4924
rect 5356 4922 5380 4924
rect 5436 4922 5442 4924
rect 5196 4870 5198 4922
rect 5378 4870 5380 4922
rect 5134 4868 5140 4870
rect 5196 4868 5220 4870
rect 5276 4868 5300 4870
rect 5356 4868 5380 4870
rect 5436 4868 5442 4870
rect 5134 4859 5442 4868
rect 5134 3836 5442 3845
rect 5134 3834 5140 3836
rect 5196 3834 5220 3836
rect 5276 3834 5300 3836
rect 5356 3834 5380 3836
rect 5436 3834 5442 3836
rect 5196 3782 5198 3834
rect 5378 3782 5380 3834
rect 5134 3780 5140 3782
rect 5196 3780 5220 3782
rect 5276 3780 5300 3782
rect 5356 3780 5380 3782
rect 5436 3780 5442 3782
rect 5134 3771 5442 3780
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4172 2446 4200 3402
rect 5276 3194 5304 3470
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5644 2990 5672 6122
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5736 2990 5764 5782
rect 5794 5468 6102 5477
rect 5794 5466 5800 5468
rect 5856 5466 5880 5468
rect 5936 5466 5960 5468
rect 6016 5466 6040 5468
rect 6096 5466 6102 5468
rect 5856 5414 5858 5466
rect 6038 5414 6040 5466
rect 5794 5412 5800 5414
rect 5856 5412 5880 5414
rect 5936 5412 5960 5414
rect 6016 5412 6040 5414
rect 6096 5412 6102 5414
rect 5794 5403 6102 5412
rect 5794 4380 6102 4389
rect 5794 4378 5800 4380
rect 5856 4378 5880 4380
rect 5936 4378 5960 4380
rect 6016 4378 6040 4380
rect 6096 4378 6102 4380
rect 5856 4326 5858 4378
rect 6038 4326 6040 4378
rect 5794 4324 5800 4326
rect 5856 4324 5880 4326
rect 5936 4324 5960 4326
rect 6016 4324 6040 4326
rect 6096 4324 6102 4326
rect 5794 4315 6102 4324
rect 6380 4146 6408 6802
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6472 4146 6500 4422
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6656 3738 6684 6734
rect 6748 5574 6776 7346
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 5794 3292 6102 3301
rect 5794 3290 5800 3292
rect 5856 3290 5880 3292
rect 5936 3290 5960 3292
rect 6016 3290 6040 3292
rect 6096 3290 6102 3292
rect 5856 3238 5858 3290
rect 6038 3238 6040 3290
rect 5794 3236 5800 3238
rect 5856 3236 5880 3238
rect 5936 3236 5960 3238
rect 6016 3236 6040 3238
rect 6096 3236 6102 3238
rect 5794 3227 6102 3236
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5134 2748 5442 2757
rect 5134 2746 5140 2748
rect 5196 2746 5220 2748
rect 5276 2746 5300 2748
rect 5356 2746 5380 2748
rect 5436 2746 5442 2748
rect 5196 2694 5198 2746
rect 5378 2694 5380 2746
rect 5134 2692 5140 2694
rect 5196 2692 5220 2694
rect 5276 2692 5300 2694
rect 5356 2692 5380 2694
rect 5436 2692 5442 2694
rect 5134 2683 5442 2692
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4894 2408 4950 2417
rect 5552 2378 5580 2926
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 5630 2544 5686 2553
rect 5630 2479 5686 2488
rect 5644 2446 5672 2479
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 4894 2343 4950 2352
rect 5540 2372 5592 2378
rect 4908 2310 4936 2343
rect 5540 2314 5592 2320
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 5736 1834 5764 2382
rect 6472 2310 6500 2790
rect 6550 2680 6606 2689
rect 6550 2615 6606 2624
rect 6564 2514 6592 2615
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 5794 2204 6102 2213
rect 5794 2202 5800 2204
rect 5856 2202 5880 2204
rect 5936 2202 5960 2204
rect 6016 2202 6040 2204
rect 6096 2202 6102 2204
rect 5856 2150 5858 2202
rect 6038 2150 6040 2202
rect 5794 2148 5800 2150
rect 5856 2148 5880 2150
rect 5936 2148 5960 2150
rect 6016 2148 6040 2150
rect 6096 2148 6102 2150
rect 5794 2139 6102 2148
rect 5724 1828 5776 1834
rect 5724 1770 5776 1776
rect 6748 1329 6776 4558
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6840 3602 6868 4422
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6932 2990 6960 6054
rect 7104 5296 7156 5302
rect 7104 5238 7156 5244
rect 7116 2990 7144 5238
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 4282 7512 5170
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7576 3058 7604 7210
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7760 4146 7788 5714
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7838 4992 7894 5001
rect 7838 4927 7894 4936
rect 7852 4146 7880 4927
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7668 2650 7696 2926
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 8036 1426 8064 5646
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4690 8340 4966
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8206 3224 8262 3233
rect 8206 3159 8208 3168
rect 8260 3159 8262 3168
rect 8208 3130 8260 3136
rect 8404 2514 8432 5034
rect 8496 4060 8524 11766
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8588 5914 8616 6190
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8588 4214 8616 5578
rect 8680 5234 8708 6666
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8496 4032 8708 4060
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8496 3058 8524 3878
rect 8588 3738 8616 3878
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8680 2774 8708 4032
rect 8772 3534 8800 6326
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8864 3398 8892 8842
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8956 2774 8984 7414
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9048 5370 9076 5646
rect 9140 5370 9168 7278
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9140 4282 9168 4558
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 8588 2746 8708 2774
rect 8864 2746 8984 2774
rect 8588 2650 8616 2746
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8864 2582 8892 2746
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 9048 2009 9076 3334
rect 9140 2990 9168 3878
rect 9232 3194 9260 11834
rect 11610 10704 11666 10713
rect 11610 10639 11666 10648
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10414 8936 10470 8945
rect 10414 8871 10470 8880
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9600 5710 9628 6054
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9310 5400 9366 5409
rect 9310 5335 9366 5344
rect 9324 4078 9352 5335
rect 9692 5166 9720 7142
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9784 4826 9812 6258
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9508 3913 9536 4014
rect 9494 3904 9550 3913
rect 9494 3839 9550 3848
rect 9600 3398 9628 4422
rect 9784 4214 9812 4490
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9784 2774 9812 4014
rect 9876 3602 9904 5102
rect 9968 4146 9996 5510
rect 10060 5234 10088 6938
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10138 5264 10194 5273
rect 10048 5228 10100 5234
rect 10138 5199 10194 5208
rect 10048 5170 10100 5176
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10048 4072 10100 4078
rect 10046 4040 10048 4049
rect 10100 4040 10102 4049
rect 10046 3975 10102 3984
rect 10152 3618 10180 5199
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9968 3590 10180 3618
rect 9968 3194 9996 3590
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9954 3088 10010 3097
rect 9954 3023 9956 3032
rect 10008 3023 10010 3032
rect 9956 2994 10008 3000
rect 9784 2746 9904 2774
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9034 2000 9090 2009
rect 9034 1935 9090 1944
rect 8024 1420 8076 1426
rect 8024 1362 8076 1368
rect 6734 1320 6790 1329
rect 6734 1255 6790 1264
rect 9048 870 9168 898
rect 9048 800 9076 870
rect 9034 0 9090 800
rect 9140 105 9168 870
rect 9600 134 9628 2382
rect 9876 1970 9904 2746
rect 9864 1964 9916 1970
rect 9864 1906 9916 1912
rect 9680 1420 9732 1426
rect 9680 1362 9732 1368
rect 9692 800 9720 1362
rect 10060 1358 10088 3470
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10152 2854 10180 3062
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10244 2038 10272 5578
rect 10232 2032 10284 2038
rect 10232 1974 10284 1980
rect 10048 1352 10100 1358
rect 10048 1294 10100 1300
rect 10336 800 10364 6598
rect 10428 5710 10456 8871
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10520 4146 10548 8026
rect 10612 5778 10640 9046
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10980 5794 11008 6326
rect 11072 5846 11100 6394
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10796 5766 11008 5794
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10598 4720 10654 4729
rect 10598 4655 10654 4664
rect 10612 4622 10640 4655
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10428 3602 10456 4014
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10508 3460 10560 3466
rect 10508 3402 10560 3408
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10428 3194 10456 3334
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10520 3058 10548 3402
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10612 2281 10640 2382
rect 10598 2272 10654 2281
rect 10598 2207 10654 2216
rect 9588 128 9640 134
rect 9126 96 9182 105
rect 9588 70 9640 76
rect 9126 31 9182 40
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10704 270 10732 4966
rect 10796 3126 10824 5766
rect 10966 5672 11022 5681
rect 10966 5607 11022 5616
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10888 3602 10916 4966
rect 10980 4146 11008 5607
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 11072 4758 11100 5034
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10966 3496 11022 3505
rect 10966 3431 11022 3440
rect 10980 3398 11008 3431
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 11164 2774 11192 6190
rect 11256 4826 11284 8910
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11256 3369 11284 4762
rect 11334 4720 11390 4729
rect 11334 4655 11390 4664
rect 11348 4622 11376 4655
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11242 3360 11298 3369
rect 11242 3295 11298 3304
rect 11256 3126 11284 3295
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 11072 2746 11192 2774
rect 11072 2310 11100 2746
rect 11440 2378 11468 6326
rect 11532 5370 11560 6666
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11624 4162 11652 10639
rect 11716 9178 11744 26206
rect 21928 24206 21956 37198
rect 22480 36922 22508 37198
rect 22572 37194 22600 37318
rect 22560 37188 22612 37194
rect 22560 37130 22612 37136
rect 22468 36916 22520 36922
rect 22468 36858 22520 36864
rect 24320 36854 24348 39200
rect 26056 37256 26108 37262
rect 26056 37198 26108 37204
rect 26068 36922 26096 37198
rect 26160 37194 26188 39200
rect 28000 37262 28028 39200
rect 27988 37256 28040 37262
rect 27988 37198 28040 37204
rect 26148 37188 26200 37194
rect 26148 37130 26200 37136
rect 26056 36916 26108 36922
rect 26056 36858 26108 36864
rect 29840 36854 29868 39200
rect 31680 37262 31708 39200
rect 33520 37330 33548 39200
rect 33508 37324 33560 37330
rect 33508 37266 33560 37272
rect 31668 37256 31720 37262
rect 31668 37198 31720 37204
rect 32680 37256 32732 37262
rect 32680 37198 32732 37204
rect 33784 37256 33836 37262
rect 33784 37198 33836 37204
rect 24308 36848 24360 36854
rect 24308 36790 24360 36796
rect 29828 36848 29880 36854
rect 29828 36790 29880 36796
rect 25780 36780 25832 36786
rect 25780 36722 25832 36728
rect 25792 36378 25820 36722
rect 32692 36417 32720 37198
rect 33048 37188 33100 37194
rect 33048 37130 33100 37136
rect 32678 36408 32734 36417
rect 25780 36372 25832 36378
rect 32678 36343 32734 36352
rect 25780 36314 25832 36320
rect 27252 32428 27304 32434
rect 27252 32370 27304 32376
rect 24952 29640 25004 29646
rect 24952 29582 25004 29588
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 12254 8664 12310 8673
rect 11704 8628 11756 8634
rect 12254 8599 12310 8608
rect 11704 8570 11756 8576
rect 11716 5234 11744 8570
rect 12070 7304 12126 7313
rect 12070 7239 12072 7248
rect 12124 7239 12126 7248
rect 12164 7268 12216 7274
rect 12072 7210 12124 7216
rect 12164 7210 12216 7216
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 6254 11836 6598
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11886 5944 11942 5953
rect 11886 5879 11942 5888
rect 11900 5778 11928 5879
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11992 4808 12020 5646
rect 11532 4146 11652 4162
rect 11520 4140 11652 4146
rect 11572 4134 11652 4140
rect 11900 4780 12020 4808
rect 11520 4082 11572 4088
rect 11518 3768 11574 3777
rect 11518 3703 11574 3712
rect 11532 3398 11560 3703
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11900 2650 11928 4780
rect 11978 4720 12034 4729
rect 11978 4655 12034 4664
rect 11992 4622 12020 4655
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11978 4176 12034 4185
rect 11978 4111 12034 4120
rect 11992 4010 12020 4111
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 12084 2650 12112 6258
rect 12176 3194 12204 7210
rect 12268 5370 12296 8599
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12360 4758 12388 11154
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12452 5234 12480 6598
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12636 4758 12664 11630
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 12990 9344 13046 9353
rect 12990 9279 13046 9288
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12728 5098 12756 7958
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12808 5092 12860 5098
rect 12808 5034 12860 5040
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12820 4622 12848 5034
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12254 4312 12310 4321
rect 12254 4247 12310 4256
rect 12268 4146 12296 4247
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12360 3602 12388 4558
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12452 4214 12480 4422
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12360 3369 12388 3402
rect 12346 3360 12402 3369
rect 12346 3295 12402 3304
rect 12360 3194 12388 3295
rect 12622 3224 12678 3233
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12348 3188 12400 3194
rect 12728 3210 12756 4490
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12820 3777 12848 4150
rect 12806 3768 12862 3777
rect 12806 3703 12862 3712
rect 12678 3182 12756 3210
rect 12622 3159 12678 3168
rect 12348 3130 12400 3136
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 11428 2372 11480 2378
rect 11428 2314 11480 2320
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 10966 1320 11022 1329
rect 10966 1255 11022 1264
rect 10980 800 11008 1255
rect 11624 800 11652 2382
rect 12084 1902 12112 2382
rect 12176 2310 12204 3130
rect 12636 3126 12664 3159
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12256 2848 12308 2854
rect 12308 2796 12388 2802
rect 12256 2790 12388 2796
rect 12268 2774 12388 2790
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12268 2106 12296 2246
rect 12256 2100 12308 2106
rect 12256 2042 12308 2048
rect 12072 1896 12124 1902
rect 12072 1838 12124 1844
rect 12360 1442 12388 2774
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 12636 2038 12664 2314
rect 12624 2032 12676 2038
rect 12624 1974 12676 1980
rect 12268 1414 12388 1442
rect 12268 800 12296 1414
rect 12912 800 12940 4422
rect 13004 3194 13032 9279
rect 13188 4214 13216 10746
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13280 6254 13308 9658
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 13096 3194 13124 3334
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13096 3058 13124 3130
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 13280 1290 13308 5646
rect 13372 5370 13400 7278
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13556 7002 13584 7142
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13636 6928 13688 6934
rect 13636 6870 13688 6876
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13464 6458 13492 6598
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13648 6118 13676 6870
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13464 5030 13492 5578
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13542 4720 13598 4729
rect 13542 4655 13544 4664
rect 13596 4655 13598 4664
rect 13544 4626 13596 4632
rect 13740 4078 13768 10678
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13728 3732 13780 3738
rect 13832 3720 13860 7346
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13780 3692 13860 3720
rect 13728 3674 13780 3680
rect 13740 2446 13768 3674
rect 13820 3120 13872 3126
rect 13818 3088 13820 3097
rect 13872 3088 13874 3097
rect 13818 3023 13874 3032
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 13268 1284 13320 1290
rect 13268 1226 13320 1232
rect 13556 800 13584 2314
rect 13924 1834 13952 6190
rect 14016 5166 14044 8434
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14108 6390 14136 7822
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14384 7410 14412 7754
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14278 7168 14334 7177
rect 14278 7103 14334 7112
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14016 3534 14044 4218
rect 14108 4146 14136 6054
rect 14200 4146 14228 6598
rect 14292 5273 14320 7103
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14278 5264 14334 5273
rect 14278 5199 14334 5208
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14292 4690 14320 4966
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14384 4536 14412 6190
rect 14292 4508 14412 4536
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14108 2514 14136 3538
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 14108 2310 14136 2450
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 13912 1828 13964 1834
rect 13912 1770 13964 1776
rect 14292 1426 14320 4508
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14384 2446 14412 4014
rect 14476 3534 14504 7686
rect 14568 5930 14596 11290
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14660 6798 14688 8366
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 14844 6866 14872 7210
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14660 6322 14688 6598
rect 14752 6322 14780 6802
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14568 5902 14688 5930
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14568 3398 14596 5714
rect 14660 5710 14688 5902
rect 14830 5808 14886 5817
rect 14830 5743 14832 5752
rect 14884 5743 14886 5752
rect 14832 5714 14884 5720
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14936 5642 14964 10202
rect 15028 7857 15056 11562
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15212 7886 15240 8230
rect 15200 7880 15252 7886
rect 15014 7848 15070 7857
rect 15200 7822 15252 7828
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15014 7783 15070 7792
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14924 5636 14976 5642
rect 14924 5578 14976 5584
rect 15028 5273 15056 7686
rect 15304 7546 15332 7822
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15384 7472 15436 7478
rect 15304 7420 15384 7426
rect 15304 7414 15436 7420
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15304 7398 15424 7414
rect 15120 5710 15148 7346
rect 15304 7342 15332 7398
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15014 5264 15070 5273
rect 15014 5199 15070 5208
rect 14648 5160 14700 5166
rect 14646 5128 14648 5137
rect 14700 5128 14702 5137
rect 14646 5063 14702 5072
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 15028 4457 15056 4558
rect 15014 4448 15070 4457
rect 15014 4383 15070 4392
rect 14832 4208 14884 4214
rect 14738 4176 14794 4185
rect 14832 4150 14884 4156
rect 14738 4111 14740 4120
rect 14792 4111 14794 4120
rect 14740 4082 14792 4088
rect 14844 3738 14872 4150
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 15120 3641 15148 4014
rect 14646 3632 14702 3641
rect 14646 3567 14702 3576
rect 15106 3632 15162 3641
rect 15106 3567 15162 3576
rect 14660 3534 14688 3567
rect 15212 3534 15240 7278
rect 15396 7041 15424 7278
rect 15382 7032 15438 7041
rect 15382 6967 15438 6976
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15304 5710 15332 6802
rect 15488 6798 15516 10542
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15304 3738 15332 5646
rect 15396 3913 15424 6598
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15382 3904 15438 3913
rect 15382 3839 15438 3848
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14924 3460 14976 3466
rect 14924 3402 14976 3408
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14752 2854 14780 3402
rect 14936 3194 14964 3402
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 15108 3120 15160 3126
rect 15106 3088 15108 3097
rect 15160 3088 15162 3097
rect 15106 3023 15162 3032
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14280 1420 14332 1426
rect 14280 1362 14332 1368
rect 15488 800 15516 6258
rect 15580 6254 15608 9114
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15660 8016 15712 8022
rect 15660 7958 15712 7964
rect 15672 6390 15700 7958
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15856 6934 15884 7754
rect 15948 7546 15976 8978
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16132 7274 16160 7482
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15660 6384 15712 6390
rect 15660 6326 15712 6332
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15566 5536 15622 5545
rect 15566 5471 15622 5480
rect 15580 5370 15608 5471
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15764 4826 15792 6734
rect 15856 5545 15884 6870
rect 15842 5536 15898 5545
rect 15842 5471 15898 5480
rect 15842 5128 15898 5137
rect 15842 5063 15898 5072
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15856 4554 15884 5063
rect 15948 4978 15976 7142
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16040 5234 16068 6054
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 15948 4950 16068 4978
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15580 2990 15608 3470
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15672 1698 15700 4422
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15752 3936 15804 3942
rect 15750 3904 15752 3913
rect 15804 3904 15806 3913
rect 15750 3839 15806 3848
rect 15948 3738 15976 4014
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15948 3194 15976 3334
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 16040 2446 16068 4950
rect 16132 4826 16160 6734
rect 16224 6322 16252 11222
rect 16592 9722 16620 12106
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17408 10192 17460 10198
rect 17222 10160 17278 10169
rect 17408 10134 17460 10140
rect 17222 10095 17278 10104
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16304 7948 16356 7954
rect 16488 7948 16540 7954
rect 16304 7890 16356 7896
rect 16408 7908 16488 7936
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16316 5953 16344 7890
rect 16408 6458 16436 7908
rect 16488 7890 16540 7896
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 16500 7410 16528 7754
rect 16592 7410 16620 8026
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16302 5944 16358 5953
rect 16302 5879 16358 5888
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16224 5166 16252 5306
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16224 4690 16252 4966
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16316 4214 16344 5646
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16408 4321 16436 5510
rect 16500 5302 16528 7210
rect 16684 6322 16712 8842
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 16762 7304 16818 7313
rect 16762 7239 16764 7248
rect 16816 7239 16818 7248
rect 16764 7210 16816 7216
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16592 5681 16620 6054
rect 16578 5672 16634 5681
rect 16578 5607 16634 5616
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16684 5302 16712 5578
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16500 4729 16528 5102
rect 16672 5092 16724 5098
rect 16672 5034 16724 5040
rect 16486 4720 16542 4729
rect 16486 4655 16542 4664
rect 16394 4312 16450 4321
rect 16394 4247 16450 4256
rect 16304 4208 16356 4214
rect 16304 4150 16356 4156
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16132 2582 16160 3878
rect 16396 3664 16448 3670
rect 16302 3632 16358 3641
rect 16592 3652 16620 3878
rect 16448 3624 16620 3652
rect 16396 3606 16448 3612
rect 16302 3567 16358 3576
rect 16316 3534 16344 3567
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16684 2650 16712 5034
rect 16776 4758 16804 5102
rect 16764 4752 16816 4758
rect 16764 4694 16816 4700
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16776 4049 16804 4150
rect 16762 4040 16818 4049
rect 16762 3975 16818 3984
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16120 2576 16172 2582
rect 16120 2518 16172 2524
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15660 1692 15712 1698
rect 15660 1634 15712 1640
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 16132 800 16160 1294
rect 16776 800 16804 3538
rect 16868 3194 16896 8366
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16960 1222 16988 5306
rect 17052 1358 17080 8366
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17144 5953 17172 7822
rect 17130 5944 17186 5953
rect 17130 5879 17186 5888
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17236 5522 17264 10095
rect 17420 7410 17448 10134
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17144 4690 17172 5510
rect 17236 5494 17356 5522
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17144 2378 17172 4218
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 17236 2106 17264 5306
rect 17328 4185 17356 5494
rect 17314 4176 17370 4185
rect 17314 4111 17370 4120
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 17328 3913 17356 3946
rect 17314 3904 17370 3913
rect 17314 3839 17370 3848
rect 17314 3360 17370 3369
rect 17314 3295 17370 3304
rect 17328 3194 17356 3295
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17314 3088 17370 3097
rect 17314 3023 17370 3032
rect 17328 2990 17356 3023
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17316 2372 17368 2378
rect 17316 2314 17368 2320
rect 17328 2145 17356 2314
rect 17314 2136 17370 2145
rect 17224 2100 17276 2106
rect 17314 2071 17370 2080
rect 17224 2042 17276 2048
rect 17420 1902 17448 6190
rect 17512 5914 17540 6734
rect 17604 6390 17632 12038
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22008 11824 22060 11830
rect 22192 11824 22244 11830
rect 22060 11784 22192 11812
rect 22008 11766 22060 11772
rect 22192 11766 22244 11772
rect 22480 11762 22508 11834
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22744 11552 22796 11558
rect 22744 11494 22796 11500
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 21730 11384 21786 11393
rect 22296 11354 22324 11494
rect 22466 11384 22522 11393
rect 21730 11319 21786 11328
rect 22284 11348 22336 11354
rect 21744 11150 21772 11319
rect 22466 11319 22522 11328
rect 22652 11348 22704 11354
rect 22284 11290 22336 11296
rect 22480 11218 22508 11319
rect 22652 11290 22704 11296
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21824 11076 21876 11082
rect 21824 11018 21876 11024
rect 22376 11076 22428 11082
rect 22376 11018 22428 11024
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17696 7426 17724 10950
rect 21836 10849 21864 11018
rect 21822 10840 21878 10849
rect 21822 10775 21878 10784
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 17958 10568 18014 10577
rect 17868 10532 17920 10538
rect 17958 10503 18014 10512
rect 17868 10474 17920 10480
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17788 8265 17816 8434
rect 17880 8294 17908 10474
rect 17972 9217 18000 10503
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18788 9648 18840 9654
rect 18788 9590 18840 9596
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 17958 9208 18014 9217
rect 17958 9143 18014 9152
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18144 8560 18196 8566
rect 18142 8528 18144 8537
rect 18196 8528 18198 8537
rect 18052 8492 18104 8498
rect 18142 8463 18198 8472
rect 18052 8434 18104 8440
rect 17868 8288 17920 8294
rect 17774 8256 17830 8265
rect 17868 8230 17920 8236
rect 17774 8191 17830 8200
rect 17696 7398 17816 7426
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17696 6458 17724 7210
rect 17788 6882 17816 7398
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17880 7002 17908 7346
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17788 6854 17908 6882
rect 17880 6474 17908 6854
rect 18064 6662 18092 8434
rect 18142 8392 18198 8401
rect 18142 8327 18144 8336
rect 18196 8327 18198 8336
rect 18144 8298 18196 8304
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17684 6452 17736 6458
rect 17880 6446 18000 6474
rect 17684 6394 17736 6400
rect 17592 6384 17644 6390
rect 17592 6326 17644 6332
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17880 6254 17908 6326
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17972 6100 18000 6446
rect 18050 6216 18106 6225
rect 18050 6151 18106 6160
rect 17880 6072 18000 6100
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17774 5808 17830 5817
rect 17774 5743 17830 5752
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17498 5536 17554 5545
rect 17498 5471 17554 5480
rect 17512 4468 17540 5471
rect 17696 5370 17724 5646
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17788 5166 17816 5743
rect 17880 5710 17908 6072
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17776 5160 17828 5166
rect 17696 5120 17776 5148
rect 17590 4720 17646 4729
rect 17590 4655 17646 4664
rect 17604 4622 17632 4655
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17696 4536 17724 5120
rect 17776 5102 17828 5108
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 4729 17816 4966
rect 17880 4865 17908 5102
rect 17866 4856 17922 4865
rect 17866 4791 17922 4800
rect 17774 4720 17830 4729
rect 17774 4655 17830 4664
rect 17868 4548 17920 4554
rect 17696 4508 17816 4536
rect 17512 4440 17632 4468
rect 17604 4146 17632 4440
rect 17682 4448 17738 4457
rect 17682 4383 17738 4392
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17590 4040 17646 4049
rect 17512 2825 17540 4014
rect 17590 3975 17646 3984
rect 17604 3194 17632 3975
rect 17696 3369 17724 4383
rect 17788 4282 17816 4508
rect 17868 4490 17920 4496
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17774 4176 17830 4185
rect 17880 4162 17908 4490
rect 17830 4134 17908 4162
rect 17774 4111 17830 4120
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17682 3360 17738 3369
rect 17682 3295 17738 3304
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17498 2816 17554 2825
rect 17498 2751 17554 2760
rect 17880 2514 17908 3538
rect 17972 3126 18000 5306
rect 18064 5030 18092 6151
rect 18052 5024 18104 5030
rect 18156 5001 18184 6734
rect 18248 5370 18276 8774
rect 18340 5409 18368 8978
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18326 5400 18382 5409
rect 18236 5364 18288 5370
rect 18326 5335 18382 5344
rect 18236 5306 18288 5312
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 18236 5160 18288 5166
rect 18340 5148 18368 5238
rect 18288 5120 18368 5148
rect 18236 5102 18288 5108
rect 18328 5024 18380 5030
rect 18052 4966 18104 4972
rect 18142 4992 18198 5001
rect 18328 4966 18380 4972
rect 18142 4927 18198 4936
rect 18142 4720 18198 4729
rect 18142 4655 18198 4664
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 18064 3398 18092 4490
rect 18156 4010 18184 4655
rect 18340 4486 18368 4966
rect 18432 4486 18460 8910
rect 18524 7834 18552 9454
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18616 8809 18644 9318
rect 18602 8800 18658 8809
rect 18602 8735 18658 8744
rect 18708 8634 18736 9318
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18800 7954 18828 9590
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 18892 8634 18920 8910
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18524 7806 18644 7834
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18524 6633 18552 7686
rect 18616 7546 18644 7806
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18510 6624 18566 6633
rect 18510 6559 18566 6568
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18524 6089 18552 6394
rect 18510 6080 18566 6089
rect 18510 6015 18566 6024
rect 18616 5574 18644 7142
rect 18604 5568 18656 5574
rect 18510 5536 18566 5545
rect 18604 5510 18656 5516
rect 18510 5471 18566 5480
rect 18524 5302 18552 5471
rect 18512 5296 18564 5302
rect 18512 5238 18564 5244
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18432 4146 18460 4422
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18142 3904 18198 3913
rect 18142 3839 18198 3848
rect 18156 3602 18184 3839
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 18064 3058 18092 3334
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 18156 2378 18184 3538
rect 18432 2854 18460 4082
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18144 2372 18196 2378
rect 18144 2314 18196 2320
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17604 1970 17632 2246
rect 17592 1964 17644 1970
rect 17592 1906 17644 1912
rect 17408 1896 17460 1902
rect 17408 1838 17460 1844
rect 18524 1834 18552 5102
rect 18616 4010 18644 5102
rect 18708 5030 18736 7686
rect 18892 7562 18920 8298
rect 18800 7534 18920 7562
rect 18800 7342 18828 7534
rect 18984 7460 19012 10406
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19168 9178 19196 10066
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 19260 9217 19288 9386
rect 19246 9208 19302 9217
rect 19156 9172 19208 9178
rect 19246 9143 19302 9152
rect 19156 9114 19208 9120
rect 19352 9110 19380 10610
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20628 10192 20680 10198
rect 20628 10134 20680 10140
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 19708 10056 19760 10062
rect 20444 10056 20496 10062
rect 19708 9998 19760 10004
rect 20442 10024 20444 10033
rect 20496 10024 20498 10033
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19444 9586 19472 9862
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19430 9344 19486 9353
rect 19430 9279 19486 9288
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19168 7886 19196 8978
rect 19444 8809 19472 9279
rect 19430 8800 19486 8809
rect 19430 8735 19486 8744
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 18892 7432 19012 7460
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18800 6458 18828 6734
rect 18788 6452 18840 6458
rect 18892 6440 18920 7432
rect 19352 7410 19380 8230
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 18984 7002 19012 7278
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 19076 6474 19104 6870
rect 19444 6866 19472 7822
rect 19536 7478 19564 9862
rect 19628 9761 19656 9998
rect 19614 9752 19670 9761
rect 19614 9687 19670 9696
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19246 6488 19302 6497
rect 19076 6458 19196 6474
rect 19076 6452 19208 6458
rect 19076 6446 19156 6452
rect 18892 6412 19012 6440
rect 18788 6394 18840 6400
rect 18984 6236 19012 6412
rect 19246 6423 19302 6432
rect 19156 6394 19208 6400
rect 19260 6390 19288 6423
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 18892 6208 19012 6236
rect 19432 6248 19484 6254
rect 18892 5778 18920 6208
rect 19432 6190 19484 6196
rect 19156 6180 19208 6186
rect 19156 6122 19208 6128
rect 19168 6089 19196 6122
rect 19248 6112 19300 6118
rect 19154 6080 19210 6089
rect 19300 6089 19380 6100
rect 19300 6080 19394 6089
rect 19300 6072 19338 6080
rect 19248 6054 19300 6060
rect 19154 6015 19210 6024
rect 19338 6015 19394 6024
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 19246 5672 19302 5681
rect 19246 5607 19302 5616
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 18616 3398 18644 3946
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 3194 18644 3334
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18694 2000 18750 2009
rect 18694 1935 18750 1944
rect 18512 1828 18564 1834
rect 18512 1770 18564 1776
rect 17040 1352 17092 1358
rect 17040 1294 17092 1300
rect 18052 1284 18104 1290
rect 18052 1226 18104 1232
rect 16948 1216 17000 1222
rect 16948 1158 17000 1164
rect 18064 800 18092 1226
rect 18708 800 18736 1935
rect 18892 1630 18920 4966
rect 18984 2038 19012 5510
rect 19062 5400 19118 5409
rect 19062 5335 19118 5344
rect 19076 4826 19104 5335
rect 19168 5137 19196 5510
rect 19260 5302 19288 5607
rect 19248 5296 19300 5302
rect 19248 5238 19300 5244
rect 19154 5128 19210 5137
rect 19154 5063 19210 5072
rect 19444 4826 19472 6190
rect 19536 5846 19564 6734
rect 19628 6322 19656 8910
rect 19720 8022 19748 9998
rect 19800 9988 19852 9994
rect 20442 9959 20498 9968
rect 19800 9930 19852 9936
rect 19812 8974 19840 9930
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19800 8968 19852 8974
rect 19800 8910 19852 8916
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19708 8016 19760 8022
rect 19708 7958 19760 7964
rect 19708 7812 19760 7818
rect 19708 7754 19760 7760
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19524 5840 19576 5846
rect 19524 5782 19576 5788
rect 19064 4820 19116 4826
rect 19064 4762 19116 4768
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19524 4752 19576 4758
rect 19524 4694 19576 4700
rect 19536 3913 19564 4694
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19522 3904 19578 3913
rect 19522 3839 19578 3848
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19352 3126 19380 3334
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 19628 2446 19656 4422
rect 19720 2990 19748 7754
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 19812 2446 19840 8774
rect 19904 8401 19932 9454
rect 20260 9444 20312 9450
rect 20260 9386 20312 9392
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19890 8392 19946 8401
rect 19890 8327 19946 8336
rect 19996 8090 20024 8434
rect 20180 8276 20208 8910
rect 20272 8430 20300 9386
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20350 8664 20406 8673
rect 20350 8599 20406 8608
rect 20364 8430 20392 8599
rect 20260 8424 20312 8430
rect 20260 8366 20312 8372
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 20180 8248 20392 8276
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 20260 8016 20312 8022
rect 20088 7964 20260 7970
rect 20088 7958 20312 7964
rect 20088 7942 20300 7958
rect 20088 6322 20116 7942
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20180 7585 20208 7822
rect 20166 7576 20222 7585
rect 20166 7511 20222 7520
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19904 6089 19932 6190
rect 19890 6080 19946 6089
rect 19890 6015 19946 6024
rect 19892 5568 19944 5574
rect 19996 5556 20024 6190
rect 20180 5914 20208 7346
rect 20272 7177 20300 7822
rect 20258 7168 20314 7177
rect 20258 7103 20314 7112
rect 20364 7018 20392 8248
rect 20272 6990 20392 7018
rect 20272 5914 20300 6990
rect 20456 6866 20484 8910
rect 20534 8392 20590 8401
rect 20534 8327 20590 8336
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20352 6180 20404 6186
rect 20352 6122 20404 6128
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 19944 5528 20024 5556
rect 20076 5568 20128 5574
rect 19892 5510 19944 5516
rect 20076 5510 20128 5516
rect 19892 4752 19944 4758
rect 19892 4694 19944 4700
rect 19904 4486 19932 4694
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19982 4312 20038 4321
rect 19982 4247 19984 4256
rect 20036 4247 20038 4256
rect 19984 4218 20036 4224
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 19904 4049 19932 4082
rect 19890 4040 19946 4049
rect 19890 3975 19946 3984
rect 20088 3738 20116 5510
rect 20180 4554 20208 5646
rect 20272 5370 20300 5850
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20168 4548 20220 4554
rect 20168 4490 20220 4496
rect 20364 4162 20392 6122
rect 20442 5944 20498 5953
rect 20442 5879 20498 5888
rect 20180 4134 20392 4162
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19904 3618 19932 3674
rect 19904 3590 20024 3618
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19904 2514 19932 3470
rect 19996 2514 20024 3590
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19800 2440 19852 2446
rect 19800 2382 19852 2388
rect 18972 2032 19024 2038
rect 18972 1974 19024 1980
rect 18880 1624 18932 1630
rect 18880 1566 18932 1572
rect 19340 1352 19392 1358
rect 19340 1294 19392 1300
rect 19352 800 19380 1294
rect 20088 1170 20116 3538
rect 20180 3233 20208 4134
rect 20260 4072 20312 4078
rect 20312 4032 20392 4060
rect 20260 4014 20312 4020
rect 20258 3768 20314 3777
rect 20258 3703 20314 3712
rect 20272 3466 20300 3703
rect 20260 3460 20312 3466
rect 20260 3402 20312 3408
rect 20166 3224 20222 3233
rect 20166 3159 20222 3168
rect 20364 2774 20392 4032
rect 20456 3942 20484 5879
rect 20548 5846 20576 8327
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20536 5296 20588 5302
rect 20536 5238 20588 5244
rect 20548 4282 20576 5238
rect 20640 4690 20668 10134
rect 20812 9920 20864 9926
rect 20810 9888 20812 9897
rect 20864 9888 20866 9897
rect 20810 9823 20866 9832
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20732 5370 20760 9454
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20824 7410 20852 9318
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20824 6066 20852 7142
rect 20916 7002 20944 10406
rect 21008 9178 21036 10610
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 21640 10532 21692 10538
rect 21640 10474 21692 10480
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21192 10305 21220 10406
rect 21178 10296 21234 10305
rect 21178 10231 21234 10240
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 21100 8090 21128 9590
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 21178 8256 21234 8265
rect 21178 8191 21234 8200
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 21192 7970 21220 8191
rect 21284 8090 21312 8978
rect 21468 8974 21496 10406
rect 21652 10062 21680 10474
rect 21824 10464 21876 10470
rect 22204 10441 22232 10542
rect 21824 10406 21876 10412
rect 22190 10432 22246 10441
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 21376 8634 21404 8774
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21560 8566 21588 9862
rect 21836 9761 21864 10406
rect 22190 10367 22246 10376
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 21822 9752 21878 9761
rect 21732 9716 21784 9722
rect 21822 9687 21878 9696
rect 21732 9658 21784 9664
rect 21744 9518 21772 9658
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21640 9104 21692 9110
rect 21640 9046 21692 9052
rect 21744 9058 21772 9454
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 21548 8560 21600 8566
rect 21548 8502 21600 8508
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21100 7942 21220 7970
rect 20994 7712 21050 7721
rect 20994 7647 21050 7656
rect 21008 7546 21036 7647
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 20996 7268 21048 7274
rect 20996 7210 21048 7216
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20824 6038 20944 6066
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20824 5817 20852 5850
rect 20810 5808 20866 5817
rect 20810 5743 20866 5752
rect 20810 5672 20866 5681
rect 20810 5607 20866 5616
rect 20824 5574 20852 5607
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20916 5409 20944 6038
rect 20902 5400 20958 5409
rect 20720 5364 20772 5370
rect 20902 5335 20958 5344
rect 20720 5306 20772 5312
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20824 3398 20852 5170
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20916 4457 20944 4558
rect 20902 4448 20958 4457
rect 20902 4383 20958 4392
rect 21008 3602 21036 7210
rect 21100 6390 21128 7942
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21192 7546 21220 7822
rect 21364 7812 21416 7818
rect 21364 7754 21416 7760
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21180 7336 21232 7342
rect 21178 7304 21180 7313
rect 21232 7304 21234 7313
rect 21178 7239 21234 7248
rect 21376 6730 21404 7754
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21454 7576 21510 7585
rect 21454 7511 21510 7520
rect 21468 7478 21496 7511
rect 21456 7472 21508 7478
rect 21456 7414 21508 7420
rect 21560 7274 21588 7686
rect 21548 7268 21600 7274
rect 21548 7210 21600 7216
rect 21364 6724 21416 6730
rect 21192 6684 21364 6712
rect 21088 6384 21140 6390
rect 21088 6326 21140 6332
rect 21192 5794 21220 6684
rect 21364 6666 21416 6672
rect 21548 6656 21600 6662
rect 21454 6624 21510 6633
rect 21548 6598 21600 6604
rect 21454 6559 21510 6568
rect 21362 6488 21418 6497
rect 21362 6423 21364 6432
rect 21416 6423 21418 6432
rect 21364 6394 21416 6400
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21100 5766 21220 5794
rect 21100 5234 21128 5766
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 21100 3194 21128 4082
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 20364 2746 20576 2774
rect 20548 2106 20576 2746
rect 20718 2680 20774 2689
rect 20718 2615 20720 2624
rect 20772 2615 20774 2624
rect 20720 2586 20772 2592
rect 21088 2304 21140 2310
rect 21086 2272 21088 2281
rect 21140 2272 21142 2281
rect 21086 2207 21142 2216
rect 20536 2100 20588 2106
rect 20536 2042 20588 2048
rect 19996 1142 20116 1170
rect 19996 800 20024 1142
rect 10692 264 10744 270
rect 10692 206 10744 212
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21192 338 21220 5646
rect 21376 5370 21404 6258
rect 21468 5914 21496 6559
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21362 5264 21418 5273
rect 21560 5234 21588 6598
rect 21652 6254 21680 9046
rect 21744 9030 21956 9058
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 21744 6186 21772 8502
rect 21732 6180 21784 6186
rect 21732 6122 21784 6128
rect 21836 6118 21864 8910
rect 21928 7562 21956 9030
rect 22020 8838 22048 9386
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 22008 8288 22060 8294
rect 22008 8230 22060 8236
rect 22020 7954 22048 8230
rect 22008 7948 22060 7954
rect 22008 7890 22060 7896
rect 21928 7534 22048 7562
rect 21914 7168 21970 7177
rect 21914 7103 21970 7112
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21652 5234 21680 5510
rect 21928 5370 21956 7103
rect 22020 6662 22048 7534
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 22020 6458 22048 6598
rect 22008 6452 22060 6458
rect 22008 6394 22060 6400
rect 22008 5908 22060 5914
rect 22008 5850 22060 5856
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21362 5199 21418 5208
rect 21548 5228 21600 5234
rect 21376 5166 21404 5199
rect 21548 5170 21600 5176
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21822 5128 21878 5137
rect 21822 5063 21878 5072
rect 21270 4856 21326 4865
rect 21270 4791 21326 4800
rect 21456 4820 21508 4826
rect 21284 3466 21312 4791
rect 21456 4762 21508 4768
rect 21364 4072 21416 4078
rect 21362 4040 21364 4049
rect 21416 4040 21418 4049
rect 21362 3975 21418 3984
rect 21272 3460 21324 3466
rect 21272 3402 21324 3408
rect 21468 3398 21496 4762
rect 21836 4758 21864 5063
rect 21732 4752 21784 4758
rect 21732 4694 21784 4700
rect 21824 4752 21876 4758
rect 21824 4694 21876 4700
rect 21548 4616 21600 4622
rect 21744 4593 21772 4694
rect 21916 4616 21968 4622
rect 21548 4558 21600 4564
rect 21730 4584 21786 4593
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21272 1420 21324 1426
rect 21272 1362 21324 1368
rect 21284 800 21312 1362
rect 21180 332 21232 338
rect 21180 274 21232 280
rect 21270 0 21326 800
rect 21560 202 21588 4558
rect 21916 4558 21968 4564
rect 21730 4519 21786 4528
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21652 3913 21680 4082
rect 21744 4078 21772 4519
rect 21928 4282 21956 4558
rect 21916 4276 21968 4282
rect 21916 4218 21968 4224
rect 21732 4072 21784 4078
rect 21732 4014 21784 4020
rect 21824 3936 21876 3942
rect 21638 3904 21694 3913
rect 21824 3878 21876 3884
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 21638 3839 21694 3848
rect 21836 3058 21864 3878
rect 21928 3466 21956 3878
rect 21916 3460 21968 3466
rect 21916 3402 21968 3408
rect 22020 3176 22048 5850
rect 21928 3148 22048 3176
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 21836 2446 21864 2790
rect 21928 2650 21956 3148
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 22020 2553 22048 2994
rect 22112 2774 22140 9862
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22204 7018 22232 8774
rect 22296 8498 22324 8774
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22388 8362 22416 11018
rect 22560 10736 22612 10742
rect 22560 10678 22612 10684
rect 22572 9586 22600 10678
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22664 8974 22692 11290
rect 22756 11257 22784 11494
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 22742 11248 22798 11257
rect 22742 11183 22744 11192
rect 22796 11183 22798 11192
rect 23202 11248 23258 11257
rect 23202 11183 23258 11192
rect 22744 11154 22796 11160
rect 23216 11082 23244 11183
rect 23204 11076 23256 11082
rect 23204 11018 23256 11024
rect 22744 11008 22796 11014
rect 22744 10950 22796 10956
rect 22756 10130 22784 10950
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 22836 10532 22888 10538
rect 22836 10474 22888 10480
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22744 9512 22796 9518
rect 22744 9454 22796 9460
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22572 8634 22600 8910
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22664 8566 22692 8910
rect 22652 8560 22704 8566
rect 22652 8502 22704 8508
rect 22560 8492 22612 8498
rect 22464 8452 22560 8480
rect 22376 8356 22428 8362
rect 22464 8344 22492 8452
rect 22560 8434 22612 8440
rect 22464 8316 22508 8344
rect 22376 8298 22428 8304
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22296 7546 22324 8230
rect 22388 7954 22416 8298
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22388 7410 22416 7890
rect 22480 7818 22508 8316
rect 22756 8294 22784 9454
rect 22848 8974 22876 10474
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22848 8634 22876 8774
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 22664 8266 22784 8294
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22468 7472 22520 7478
rect 22466 7440 22468 7449
rect 22520 7440 22522 7449
rect 22376 7404 22428 7410
rect 22466 7375 22522 7384
rect 22376 7346 22428 7352
rect 22282 7032 22338 7041
rect 22204 6990 22282 7018
rect 22282 6967 22338 6976
rect 22190 6760 22246 6769
rect 22296 6746 22324 6967
rect 22388 6866 22416 7346
rect 22664 6984 22692 8266
rect 22742 7984 22798 7993
rect 22742 7919 22798 7928
rect 22480 6956 22692 6984
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22296 6718 22416 6746
rect 22190 6695 22246 6704
rect 22204 6118 22232 6695
rect 22284 6656 22336 6662
rect 22284 6598 22336 6604
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22296 5846 22324 6598
rect 22388 6390 22416 6718
rect 22376 6384 22428 6390
rect 22376 6326 22428 6332
rect 22284 5840 22336 5846
rect 22284 5782 22336 5788
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22204 5574 22232 5646
rect 22192 5568 22244 5574
rect 22480 5545 22508 6956
rect 22558 6896 22614 6905
rect 22558 6831 22614 6840
rect 22572 6798 22600 6831
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22652 6724 22704 6730
rect 22652 6666 22704 6672
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22572 5778 22600 6598
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 22192 5510 22244 5516
rect 22466 5536 22522 5545
rect 22466 5471 22522 5480
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22190 4312 22246 4321
rect 22190 4247 22246 4256
rect 22204 3466 22232 4247
rect 22296 4078 22324 4422
rect 22480 4282 22508 5471
rect 22664 5386 22692 6666
rect 22756 6254 22784 7919
rect 22744 6248 22796 6254
rect 22744 6190 22796 6196
rect 22572 5358 22692 5386
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22376 4004 22428 4010
rect 22376 3946 22428 3952
rect 22388 3670 22416 3946
rect 22376 3664 22428 3670
rect 22376 3606 22428 3612
rect 22192 3460 22244 3466
rect 22192 3402 22244 3408
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 22112 2746 22232 2774
rect 22006 2544 22062 2553
rect 22006 2479 22062 2488
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 21836 1902 21864 2382
rect 21824 1896 21876 1902
rect 21824 1838 21876 1844
rect 22204 1426 22232 2746
rect 22480 2446 22508 3402
rect 22572 2582 22600 5358
rect 22744 5296 22796 5302
rect 22744 5238 22796 5244
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 22664 3194 22692 4558
rect 22756 4214 22784 5238
rect 22744 4208 22796 4214
rect 22744 4150 22796 4156
rect 22744 4004 22796 4010
rect 22848 3992 22876 8434
rect 22940 7154 22968 10610
rect 23032 9926 23060 10610
rect 23308 10606 23336 11290
rect 23492 11286 23520 11494
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23952 11218 23980 11766
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 24216 11552 24268 11558
rect 24216 11494 24268 11500
rect 24228 11218 24256 11494
rect 23940 11212 23992 11218
rect 23940 11154 23992 11160
rect 24216 11212 24268 11218
rect 24216 11154 24268 11160
rect 23386 11112 23442 11121
rect 23386 11047 23388 11056
rect 23440 11047 23442 11056
rect 23480 11076 23532 11082
rect 23388 11018 23440 11024
rect 23480 11018 23532 11024
rect 23296 10600 23348 10606
rect 23296 10542 23348 10548
rect 23112 10464 23164 10470
rect 23112 10406 23164 10412
rect 23124 10266 23152 10406
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 23020 9920 23072 9926
rect 23020 9862 23072 9868
rect 23018 8936 23074 8945
rect 23018 8871 23020 8880
rect 23072 8871 23074 8880
rect 23112 8900 23164 8906
rect 23020 8842 23072 8848
rect 23112 8842 23164 8848
rect 23124 8294 23152 8842
rect 23112 8288 23164 8294
rect 23112 8230 23164 8236
rect 22940 7126 23152 7154
rect 22928 6996 22980 7002
rect 22928 6938 22980 6944
rect 22796 3964 22876 3992
rect 22744 3946 22796 3952
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22836 2848 22888 2854
rect 22836 2790 22888 2796
rect 22560 2576 22612 2582
rect 22560 2518 22612 2524
rect 22468 2440 22520 2446
rect 22468 2382 22520 2388
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 22192 1420 22244 1426
rect 22192 1362 22244 1368
rect 21836 870 21956 898
rect 21836 270 21864 870
rect 21928 800 21956 870
rect 22572 800 22600 2382
rect 22848 2009 22876 2790
rect 22940 2774 22968 6938
rect 23018 5672 23074 5681
rect 23018 5607 23074 5616
rect 23032 5370 23060 5607
rect 23020 5364 23072 5370
rect 23020 5306 23072 5312
rect 23124 5030 23152 7126
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 23032 3194 23060 4558
rect 23124 3942 23152 4966
rect 23216 4826 23244 10066
rect 23308 10062 23336 10542
rect 23296 10056 23348 10062
rect 23492 10033 23520 11018
rect 24032 11008 24084 11014
rect 24032 10950 24084 10956
rect 24124 11008 24176 11014
rect 24124 10950 24176 10956
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 23296 9998 23348 10004
rect 23478 10024 23534 10033
rect 23478 9959 23534 9968
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23480 9920 23532 9926
rect 23584 9908 23612 10542
rect 24044 10266 24072 10950
rect 24136 10606 24164 10950
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24124 10464 24176 10470
rect 24124 10406 24176 10412
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 23756 9988 23808 9994
rect 23756 9930 23808 9936
rect 23532 9880 23612 9908
rect 23480 9862 23532 9868
rect 23308 8974 23336 9862
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23400 8820 23428 9522
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23308 8792 23428 8820
rect 23308 6497 23336 8792
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23400 7206 23428 8570
rect 23492 8022 23520 9318
rect 23480 8016 23532 8022
rect 23480 7958 23532 7964
rect 23584 7954 23612 9880
rect 23768 9450 23796 9930
rect 23756 9444 23808 9450
rect 23756 9386 23808 9392
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23388 6928 23440 6934
rect 23388 6870 23440 6876
rect 23294 6488 23350 6497
rect 23294 6423 23296 6432
rect 23348 6423 23350 6432
rect 23296 6394 23348 6400
rect 23400 6322 23428 6870
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 23202 4312 23258 4321
rect 23202 4247 23204 4256
rect 23256 4247 23258 4256
rect 23204 4218 23256 4224
rect 23308 4162 23336 6258
rect 23388 5772 23440 5778
rect 23388 5714 23440 5720
rect 23400 5545 23428 5714
rect 23386 5536 23442 5545
rect 23386 5471 23442 5480
rect 23492 5370 23520 7346
rect 23584 7342 23612 7890
rect 23572 7336 23624 7342
rect 23572 7278 23624 7284
rect 23572 7200 23624 7206
rect 23572 7142 23624 7148
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23584 5098 23612 7142
rect 23388 5092 23440 5098
rect 23388 5034 23440 5040
rect 23572 5092 23624 5098
rect 23572 5034 23624 5040
rect 23400 4622 23428 5034
rect 23570 4856 23626 4865
rect 23570 4791 23626 4800
rect 23584 4690 23612 4791
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 23676 4162 23704 9318
rect 23756 8968 23808 8974
rect 23756 8910 23808 8916
rect 23768 7721 23796 8910
rect 23860 8566 23888 9318
rect 23940 8900 23992 8906
rect 23940 8842 23992 8848
rect 23848 8560 23900 8566
rect 23848 8502 23900 8508
rect 23848 8288 23900 8294
rect 23848 8230 23900 8236
rect 23860 7818 23888 8230
rect 23848 7812 23900 7818
rect 23848 7754 23900 7760
rect 23754 7712 23810 7721
rect 23754 7647 23810 7656
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 23768 7002 23796 7278
rect 23846 7032 23902 7041
rect 23756 6996 23808 7002
rect 23846 6967 23902 6976
rect 23756 6938 23808 6944
rect 23754 6488 23810 6497
rect 23754 6423 23810 6432
rect 23768 6322 23796 6423
rect 23860 6322 23888 6967
rect 23952 6866 23980 8842
rect 24032 7744 24084 7750
rect 24032 7686 24084 7692
rect 24044 7313 24072 7686
rect 24030 7304 24086 7313
rect 24030 7239 24086 7248
rect 24032 6996 24084 7002
rect 24032 6938 24084 6944
rect 23940 6860 23992 6866
rect 23940 6802 23992 6808
rect 24044 6458 24072 6938
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 24030 6352 24086 6361
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23848 6316 23900 6322
rect 24030 6287 24086 6296
rect 23848 6258 23900 6264
rect 23940 6248 23992 6254
rect 23940 6190 23992 6196
rect 23952 5914 23980 6190
rect 24044 5953 24072 6287
rect 24030 5944 24086 5953
rect 23940 5908 23992 5914
rect 24030 5879 24086 5888
rect 23940 5850 23992 5856
rect 23756 5840 23808 5846
rect 24136 5794 24164 10406
rect 24228 9625 24256 11154
rect 24214 9616 24270 9625
rect 24214 9551 24270 9560
rect 24216 9444 24268 9450
rect 24216 9386 24268 9392
rect 24228 8974 24256 9386
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 24216 8832 24268 8838
rect 24320 8809 24348 11698
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 24688 11150 24716 11494
rect 24872 11354 24900 14418
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24872 11150 24900 11290
rect 24964 11150 24992 29582
rect 26240 26920 26292 26926
rect 26240 26862 26292 26868
rect 26252 16574 26280 26862
rect 27264 16574 27292 32370
rect 28724 21412 28776 21418
rect 28724 21354 28776 21360
rect 26252 16546 26372 16574
rect 25320 12096 25372 12102
rect 25320 12038 25372 12044
rect 25228 11552 25280 11558
rect 25226 11520 25228 11529
rect 25280 11520 25282 11529
rect 25226 11455 25282 11464
rect 25240 11218 25268 11455
rect 25332 11354 25360 12038
rect 25964 11552 26016 11558
rect 25964 11494 26016 11500
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25228 11212 25280 11218
rect 25228 11154 25280 11160
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 24964 11014 24992 11086
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 24400 10668 24452 10674
rect 24400 10610 24452 10616
rect 24412 9110 24440 10610
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24492 10056 24544 10062
rect 24492 9998 24544 10004
rect 24400 9104 24452 9110
rect 24400 9046 24452 9052
rect 24216 8774 24268 8780
rect 24306 8800 24362 8809
rect 24228 8566 24256 8774
rect 24306 8735 24362 8744
rect 24398 8664 24454 8673
rect 24308 8628 24360 8634
rect 24398 8599 24454 8608
rect 24308 8570 24360 8576
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 24320 7834 24348 8570
rect 23756 5782 23808 5788
rect 23216 4134 23336 4162
rect 23388 4140 23440 4146
rect 23112 3936 23164 3942
rect 23112 3878 23164 3884
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 22940 2746 23060 2774
rect 22926 2680 22982 2689
rect 22926 2615 22982 2624
rect 22940 2310 22968 2615
rect 23032 2446 23060 2746
rect 23216 2650 23244 4134
rect 23388 4082 23440 4088
rect 23584 4134 23704 4162
rect 23400 4026 23428 4082
rect 23584 4026 23612 4134
rect 23400 3998 23612 4026
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 23400 3058 23428 3470
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23204 2644 23256 2650
rect 23204 2586 23256 2592
rect 23676 2582 23704 4014
rect 23768 2990 23796 5782
rect 24044 5766 24164 5794
rect 24228 7806 24348 7834
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23860 4214 23888 5170
rect 24044 4622 24072 5766
rect 24228 5710 24256 7806
rect 24306 7712 24362 7721
rect 24306 7647 24362 7656
rect 24320 7546 24348 7647
rect 24308 7540 24360 7546
rect 24308 7482 24360 7488
rect 24412 7426 24440 8599
rect 24320 7398 24440 7426
rect 24320 5914 24348 7398
rect 24398 6488 24454 6497
rect 24398 6423 24400 6432
rect 24452 6423 24454 6432
rect 24400 6394 24452 6400
rect 24308 5908 24360 5914
rect 24308 5850 24360 5856
rect 24308 5772 24360 5778
rect 24308 5714 24360 5720
rect 24216 5704 24268 5710
rect 24122 5672 24178 5681
rect 24216 5646 24268 5652
rect 24122 5607 24178 5616
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 23848 4208 23900 4214
rect 23848 4150 23900 4156
rect 24032 4208 24084 4214
rect 24032 4150 24084 4156
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 23664 2576 23716 2582
rect 23664 2518 23716 2524
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 22928 2304 22980 2310
rect 22928 2246 22980 2252
rect 22834 2000 22890 2009
rect 22834 1935 22890 1944
rect 23952 1766 23980 4082
rect 24044 3534 24072 4150
rect 24136 4078 24164 5607
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24228 4146 24256 5306
rect 24320 5001 24348 5714
rect 24400 5092 24452 5098
rect 24400 5034 24452 5040
rect 24306 4992 24362 5001
rect 24306 4927 24362 4936
rect 24308 4684 24360 4690
rect 24308 4626 24360 4632
rect 24320 4593 24348 4626
rect 24306 4584 24362 4593
rect 24306 4519 24362 4528
rect 24320 4282 24348 4519
rect 24308 4276 24360 4282
rect 24308 4218 24360 4224
rect 24216 4140 24268 4146
rect 24216 4082 24268 4088
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 24228 3398 24256 4082
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24412 2854 24440 5034
rect 24504 4826 24532 9998
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24492 4820 24544 4826
rect 24492 4762 24544 4768
rect 24596 4706 24624 9862
rect 24688 9761 24716 9862
rect 24674 9752 24730 9761
rect 24674 9687 24730 9696
rect 24780 9450 24808 10474
rect 24858 10024 24914 10033
rect 24858 9959 24914 9968
rect 24768 9444 24820 9450
rect 24768 9386 24820 9392
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24688 6610 24716 9114
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24780 8265 24808 8910
rect 24766 8256 24822 8265
rect 24766 8191 24822 8200
rect 24768 7948 24820 7954
rect 24768 7890 24820 7896
rect 24780 7857 24808 7890
rect 24766 7848 24822 7857
rect 24766 7783 24822 7792
rect 24768 7472 24820 7478
rect 24768 7414 24820 7420
rect 24780 6730 24808 7414
rect 24872 6866 24900 9959
rect 25056 7721 25084 11086
rect 25318 10840 25374 10849
rect 25318 10775 25374 10784
rect 25228 10464 25280 10470
rect 25228 10406 25280 10412
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25148 9586 25176 9862
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 25148 8090 25176 8774
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 25042 7712 25098 7721
rect 25042 7647 25098 7656
rect 24950 7576 25006 7585
rect 24950 7511 25006 7520
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 24688 6582 24808 6610
rect 24674 6488 24730 6497
rect 24674 6423 24730 6432
rect 24688 5846 24716 6423
rect 24676 5840 24728 5846
rect 24676 5782 24728 5788
rect 24674 5400 24730 5409
rect 24674 5335 24730 5344
rect 24504 4678 24624 4706
rect 24504 3126 24532 4678
rect 24688 4622 24716 5335
rect 24780 4690 24808 6582
rect 24964 5574 24992 7511
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 25056 6118 25084 6258
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 25136 6112 25188 6118
rect 25136 6054 25188 6060
rect 25056 5642 25084 6054
rect 25148 5846 25176 6054
rect 25136 5840 25188 5846
rect 25136 5782 25188 5788
rect 25134 5672 25190 5681
rect 25044 5636 25096 5642
rect 25134 5607 25190 5616
rect 25044 5578 25096 5584
rect 24952 5568 25004 5574
rect 24952 5510 25004 5516
rect 24858 5264 24914 5273
rect 24858 5199 24860 5208
rect 24912 5199 24914 5208
rect 24860 5170 24912 5176
rect 25056 4690 25084 5578
rect 24768 4684 24820 4690
rect 24768 4626 24820 4632
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 24676 4616 24728 4622
rect 24676 4558 24728 4564
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24582 4176 24638 4185
rect 24582 4111 24638 4120
rect 24596 4078 24624 4111
rect 24584 4072 24636 4078
rect 24584 4014 24636 4020
rect 24780 3641 24808 4422
rect 24964 4214 24992 4490
rect 24952 4208 25004 4214
rect 24952 4150 25004 4156
rect 24950 3904 25006 3913
rect 24950 3839 25006 3848
rect 24964 3670 24992 3839
rect 24952 3664 25004 3670
rect 24766 3632 24822 3641
rect 24952 3606 25004 3612
rect 24766 3567 24822 3576
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24492 3120 24544 3126
rect 24492 3062 24544 3068
rect 24780 3058 24808 3334
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 24860 3052 24912 3058
rect 25148 3040 25176 5607
rect 25240 3534 25268 10406
rect 25332 9586 25360 10775
rect 25976 9674 26004 11494
rect 26054 11384 26110 11393
rect 26054 11319 26056 11328
rect 26108 11319 26110 11328
rect 26056 11290 26108 11296
rect 26238 11248 26294 11257
rect 26238 11183 26240 11192
rect 26292 11183 26294 11192
rect 26240 11154 26292 11160
rect 26054 10704 26110 10713
rect 26054 10639 26056 10648
rect 26108 10639 26110 10648
rect 26056 10610 26108 10616
rect 26344 10130 26372 16546
rect 26988 16546 27292 16574
rect 26988 12434 27016 16546
rect 27436 14544 27488 14550
rect 27436 14486 27488 14492
rect 27448 12434 27476 14486
rect 28736 12434 28764 21354
rect 26712 12406 27016 12434
rect 27356 12406 27476 12434
rect 28552 12406 28764 12434
rect 26424 11824 26476 11830
rect 26424 11766 26476 11772
rect 26436 10606 26464 11766
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26528 10674 26556 11494
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 26424 10600 26476 10606
rect 26424 10542 26476 10548
rect 26332 10124 26384 10130
rect 26332 10066 26384 10072
rect 26344 9761 26372 10066
rect 26330 9752 26386 9761
rect 26436 9722 26464 10542
rect 26516 10532 26568 10538
rect 26516 10474 26568 10480
rect 26330 9687 26386 9696
rect 26424 9716 26476 9722
rect 25596 9648 25648 9654
rect 25976 9646 26096 9674
rect 26424 9658 26476 9664
rect 25596 9590 25648 9596
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 25320 8968 25372 8974
rect 25320 8910 25372 8916
rect 25332 8401 25360 8910
rect 25318 8392 25374 8401
rect 25318 8327 25374 8336
rect 25412 8084 25464 8090
rect 25412 8026 25464 8032
rect 25320 7880 25372 7886
rect 25320 7822 25372 7828
rect 25332 7750 25360 7822
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25424 6934 25452 8026
rect 25412 6928 25464 6934
rect 25412 6870 25464 6876
rect 25320 6248 25372 6254
rect 25320 6190 25372 6196
rect 25332 5778 25360 6190
rect 25320 5772 25372 5778
rect 25320 5714 25372 5720
rect 25320 3664 25372 3670
rect 25320 3606 25372 3612
rect 25332 3534 25360 3606
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 25424 3398 25452 6870
rect 25504 6792 25556 6798
rect 25502 6760 25504 6769
rect 25556 6760 25558 6769
rect 25502 6695 25558 6704
rect 25504 5772 25556 5778
rect 25504 5714 25556 5720
rect 25516 5681 25544 5714
rect 25502 5672 25558 5681
rect 25502 5607 25558 5616
rect 25608 5574 25636 9590
rect 25964 9512 26016 9518
rect 25962 9480 25964 9489
rect 26016 9480 26018 9489
rect 25962 9415 26018 9424
rect 25872 9376 25924 9382
rect 25872 9318 25924 9324
rect 25884 8945 25912 9318
rect 25870 8936 25926 8945
rect 25870 8871 25926 8880
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 25884 8566 25912 8774
rect 25872 8560 25924 8566
rect 25872 8502 25924 8508
rect 25780 8356 25832 8362
rect 25780 8298 25832 8304
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25700 7886 25728 8026
rect 25792 7886 25820 8298
rect 25884 8129 25912 8502
rect 25964 8424 26016 8430
rect 26068 8412 26096 9646
rect 26240 8832 26292 8838
rect 26240 8774 26292 8780
rect 26252 8566 26280 8774
rect 26528 8616 26556 10474
rect 26620 9586 26648 11494
rect 26608 9580 26660 9586
rect 26608 9522 26660 9528
rect 26712 9466 26740 12406
rect 27252 11892 27304 11898
rect 27252 11834 27304 11840
rect 26884 11620 26936 11626
rect 26884 11562 26936 11568
rect 26896 11286 26924 11562
rect 26884 11280 26936 11286
rect 26884 11222 26936 11228
rect 26976 11144 27028 11150
rect 26976 11086 27028 11092
rect 26884 11076 26936 11082
rect 26884 11018 26936 11024
rect 26792 10736 26844 10742
rect 26792 10678 26844 10684
rect 26620 9438 26740 9466
rect 26620 8838 26648 9438
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26344 8588 26556 8616
rect 26240 8560 26292 8566
rect 26240 8502 26292 8508
rect 26016 8384 26096 8412
rect 26344 8378 26372 8588
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 25964 8366 26016 8372
rect 25870 8120 25926 8129
rect 25870 8055 25926 8064
rect 25872 8016 25924 8022
rect 25872 7958 25924 7964
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 25780 7880 25832 7886
rect 25780 7822 25832 7828
rect 25780 7744 25832 7750
rect 25686 7712 25742 7721
rect 25780 7686 25832 7692
rect 25686 7647 25742 7656
rect 25700 6798 25728 7647
rect 25792 6905 25820 7686
rect 25778 6896 25834 6905
rect 25778 6831 25834 6840
rect 25688 6792 25740 6798
rect 25688 6734 25740 6740
rect 25686 6080 25742 6089
rect 25686 6015 25742 6024
rect 25700 5710 25728 6015
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25596 5568 25648 5574
rect 25792 5556 25820 6831
rect 25884 5778 25912 7958
rect 25976 7750 26004 8366
rect 26252 8350 26372 8378
rect 26056 8288 26108 8294
rect 26056 8230 26108 8236
rect 26068 7954 26096 8230
rect 26056 7948 26108 7954
rect 26056 7890 26108 7896
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 25964 7336 26016 7342
rect 25964 7278 26016 7284
rect 25976 6934 26004 7278
rect 26056 7200 26108 7206
rect 26056 7142 26108 7148
rect 26146 7168 26202 7177
rect 26068 7002 26096 7142
rect 26146 7103 26202 7112
rect 26056 6996 26108 7002
rect 26056 6938 26108 6944
rect 25964 6928 26016 6934
rect 25964 6870 26016 6876
rect 26160 6322 26188 7103
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 25872 5772 25924 5778
rect 25872 5714 25924 5720
rect 26148 5704 26200 5710
rect 26148 5646 26200 5652
rect 25872 5636 25924 5642
rect 25872 5578 25924 5584
rect 25596 5510 25648 5516
rect 25700 5528 25820 5556
rect 25502 5400 25558 5409
rect 25502 5335 25504 5344
rect 25556 5335 25558 5344
rect 25504 5306 25556 5312
rect 25594 4312 25650 4321
rect 25594 4247 25650 4256
rect 25608 3942 25636 4247
rect 25596 3936 25648 3942
rect 25596 3878 25648 3884
rect 25594 3768 25650 3777
rect 25594 3703 25650 3712
rect 25608 3466 25636 3703
rect 25700 3670 25728 5528
rect 25884 5234 25912 5578
rect 26160 5522 26188 5646
rect 25976 5494 26188 5522
rect 25872 5228 25924 5234
rect 25872 5170 25924 5176
rect 25870 4448 25926 4457
rect 25870 4383 25926 4392
rect 25688 3664 25740 3670
rect 25688 3606 25740 3612
rect 25884 3466 25912 4383
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 25872 3460 25924 3466
rect 25872 3402 25924 3408
rect 25412 3392 25464 3398
rect 25688 3392 25740 3398
rect 25412 3334 25464 3340
rect 25686 3360 25688 3369
rect 25740 3360 25742 3369
rect 25686 3295 25742 3304
rect 25504 3120 25556 3126
rect 25504 3062 25556 3068
rect 25228 3052 25280 3058
rect 25148 3012 25228 3040
rect 24860 2994 24912 3000
rect 25228 2994 25280 3000
rect 24400 2848 24452 2854
rect 24400 2790 24452 2796
rect 24780 2514 24808 2994
rect 24872 2922 24900 2994
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 24768 2508 24820 2514
rect 24768 2450 24820 2456
rect 25516 2378 25544 3062
rect 25884 2632 25912 3402
rect 25976 3194 26004 5494
rect 26148 5364 26200 5370
rect 26148 5306 26200 5312
rect 26160 5148 26188 5306
rect 26252 5250 26280 8350
rect 26332 8288 26384 8294
rect 26332 8230 26384 8236
rect 26344 5914 26372 8230
rect 26436 7410 26464 8434
rect 26620 8430 26648 8774
rect 26608 8424 26660 8430
rect 26608 8366 26660 8372
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26608 7744 26660 7750
rect 26608 7686 26660 7692
rect 26424 7404 26476 7410
rect 26424 7346 26476 7352
rect 26332 5908 26384 5914
rect 26332 5850 26384 5856
rect 26436 5370 26464 7346
rect 26516 7336 26568 7342
rect 26516 7278 26568 7284
rect 26528 6866 26556 7278
rect 26620 7002 26648 7686
rect 26608 6996 26660 7002
rect 26608 6938 26660 6944
rect 26606 6896 26662 6905
rect 26516 6860 26568 6866
rect 26606 6831 26662 6840
rect 26516 6802 26568 6808
rect 26620 6662 26648 6831
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 26424 5364 26476 5370
rect 26424 5306 26476 5312
rect 26252 5222 26556 5250
rect 26160 5120 26280 5148
rect 26252 4554 26280 5120
rect 26422 4720 26478 4729
rect 26332 4684 26384 4690
rect 26422 4655 26424 4664
rect 26332 4626 26384 4632
rect 26476 4655 26478 4664
rect 26424 4626 26476 4632
rect 26240 4548 26292 4554
rect 26240 4490 26292 4496
rect 26148 4072 26200 4078
rect 26148 4014 26200 4020
rect 26160 3913 26188 4014
rect 26146 3904 26202 3913
rect 26068 3862 26146 3890
rect 25964 3188 26016 3194
rect 25964 3130 26016 3136
rect 26068 3126 26096 3862
rect 26146 3839 26202 3848
rect 26146 3496 26202 3505
rect 26146 3431 26148 3440
rect 26200 3431 26202 3440
rect 26148 3402 26200 3408
rect 26252 3398 26280 4490
rect 26344 3913 26372 4626
rect 26424 4140 26476 4146
rect 26424 4082 26476 4088
rect 26330 3904 26386 3913
rect 26330 3839 26386 3848
rect 26436 3602 26464 4082
rect 26528 3670 26556 5222
rect 26516 3664 26568 3670
rect 26516 3606 26568 3612
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26056 3120 26108 3126
rect 26056 3062 26108 3068
rect 25964 2644 26016 2650
rect 25884 2604 25964 2632
rect 25964 2586 26016 2592
rect 26252 2378 26280 3334
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 25504 2372 25556 2378
rect 25504 2314 25556 2320
rect 25596 2372 25648 2378
rect 25596 2314 25648 2320
rect 26240 2372 26292 2378
rect 26240 2314 26292 2320
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 23940 1760 23992 1766
rect 23940 1702 23992 1708
rect 23204 1420 23256 1426
rect 23204 1362 23256 1368
rect 23216 800 23244 1362
rect 23768 870 23888 898
rect 21824 264 21876 270
rect 21824 206 21876 212
rect 21548 196 21600 202
rect 21548 138 21600 144
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23768 134 23796 870
rect 23860 800 23888 870
rect 24504 800 24532 2246
rect 25608 1698 25636 2314
rect 25596 1692 25648 1698
rect 25596 1634 25648 1640
rect 25780 1216 25832 1222
rect 25780 1158 25832 1164
rect 25056 870 25176 898
rect 23756 128 23808 134
rect 23756 70 23808 76
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25056 241 25084 870
rect 25148 800 25176 870
rect 25792 800 25820 1158
rect 26436 800 26464 2926
rect 26528 2922 26556 3606
rect 26516 2916 26568 2922
rect 26516 2858 26568 2864
rect 26620 2774 26648 6598
rect 26712 6458 26740 7822
rect 26700 6452 26752 6458
rect 26700 6394 26752 6400
rect 26804 6390 26832 10678
rect 26896 9586 26924 11018
rect 26884 9580 26936 9586
rect 26884 9522 26936 9528
rect 26884 8356 26936 8362
rect 26884 8298 26936 8304
rect 26896 7954 26924 8298
rect 26884 7948 26936 7954
rect 26884 7890 26936 7896
rect 26884 7744 26936 7750
rect 26884 7686 26936 7692
rect 26896 7478 26924 7686
rect 26884 7472 26936 7478
rect 26884 7414 26936 7420
rect 26792 6384 26844 6390
rect 26792 6326 26844 6332
rect 26792 6248 26844 6254
rect 26792 6190 26844 6196
rect 26700 5568 26752 5574
rect 26700 5510 26752 5516
rect 26712 3058 26740 5510
rect 26700 3052 26752 3058
rect 26700 2994 26752 3000
rect 26804 2990 26832 6190
rect 26988 5794 27016 11086
rect 27068 10600 27120 10606
rect 27068 10542 27120 10548
rect 27080 10266 27108 10542
rect 27068 10260 27120 10266
rect 27068 10202 27120 10208
rect 27264 10146 27292 11834
rect 27080 10118 27292 10146
rect 27080 7993 27108 10118
rect 27356 10010 27384 12406
rect 27436 11892 27488 11898
rect 27436 11834 27488 11840
rect 27448 11694 27476 11834
rect 27896 11756 27948 11762
rect 27896 11698 27948 11704
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27436 11008 27488 11014
rect 27436 10950 27488 10956
rect 27448 10062 27476 10950
rect 27528 10464 27580 10470
rect 27528 10406 27580 10412
rect 27620 10464 27672 10470
rect 27620 10406 27672 10412
rect 27172 9982 27384 10010
rect 27436 10056 27488 10062
rect 27436 9998 27488 10004
rect 27172 8430 27200 9982
rect 27540 9926 27568 10406
rect 27632 10169 27660 10406
rect 27618 10160 27674 10169
rect 27618 10095 27674 10104
rect 27712 10124 27764 10130
rect 27712 10066 27764 10072
rect 27724 10033 27752 10066
rect 27710 10024 27766 10033
rect 27620 9988 27672 9994
rect 27710 9959 27766 9968
rect 27620 9930 27672 9936
rect 27252 9920 27304 9926
rect 27252 9862 27304 9868
rect 27528 9920 27580 9926
rect 27528 9862 27580 9868
rect 27160 8424 27212 8430
rect 27160 8366 27212 8372
rect 27172 8090 27200 8366
rect 27160 8084 27212 8090
rect 27160 8026 27212 8032
rect 27066 7984 27122 7993
rect 27066 7919 27122 7928
rect 27068 7880 27120 7886
rect 27068 7822 27120 7828
rect 27080 5914 27108 7822
rect 27172 7750 27200 8026
rect 27160 7744 27212 7750
rect 27160 7686 27212 7692
rect 27160 7404 27212 7410
rect 27160 7346 27212 7352
rect 27068 5908 27120 5914
rect 27068 5850 27120 5856
rect 26988 5766 27108 5794
rect 26884 5024 26936 5030
rect 26884 4966 26936 4972
rect 26976 5024 27028 5030
rect 26976 4966 27028 4972
rect 26896 4690 26924 4966
rect 26884 4684 26936 4690
rect 26884 4626 26936 4632
rect 26988 4214 27016 4966
rect 26976 4208 27028 4214
rect 26976 4150 27028 4156
rect 26884 4072 26936 4078
rect 26884 4014 26936 4020
rect 26896 3058 26924 4014
rect 26974 3360 27030 3369
rect 26974 3295 27030 3304
rect 26988 3194 27016 3295
rect 26976 3188 27028 3194
rect 26976 3130 27028 3136
rect 26884 3052 26936 3058
rect 26884 2994 26936 3000
rect 26792 2984 26844 2990
rect 26792 2926 26844 2932
rect 26988 2854 27016 3130
rect 26976 2848 27028 2854
rect 26976 2790 27028 2796
rect 26620 2746 26832 2774
rect 26804 2514 26832 2746
rect 26792 2508 26844 2514
rect 26792 2450 26844 2456
rect 27080 800 27108 5766
rect 27172 2650 27200 7346
rect 27264 3466 27292 9862
rect 27344 9376 27396 9382
rect 27344 9318 27396 9324
rect 27356 8090 27384 9318
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 27448 8673 27476 9114
rect 27434 8664 27490 8673
rect 27434 8599 27490 8608
rect 27528 8560 27580 8566
rect 27528 8502 27580 8508
rect 27434 8256 27490 8265
rect 27434 8191 27490 8200
rect 27344 8084 27396 8090
rect 27344 8026 27396 8032
rect 27448 6100 27476 8191
rect 27540 6390 27568 8502
rect 27632 7546 27660 9930
rect 27908 9586 27936 11698
rect 28448 11688 28500 11694
rect 28446 11656 28448 11665
rect 28500 11656 28502 11665
rect 28446 11591 28502 11600
rect 28356 11552 28408 11558
rect 28356 11494 28408 11500
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 27896 9580 27948 9586
rect 27896 9522 27948 9528
rect 27896 9444 27948 9450
rect 27896 9386 27948 9392
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27816 9042 27844 9318
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 27712 8424 27764 8430
rect 27712 8366 27764 8372
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27724 6458 27752 8366
rect 27712 6452 27764 6458
rect 27712 6394 27764 6400
rect 27528 6384 27580 6390
rect 27528 6326 27580 6332
rect 27620 6384 27672 6390
rect 27620 6326 27672 6332
rect 27448 6072 27568 6100
rect 27436 5908 27488 5914
rect 27436 5850 27488 5856
rect 27342 5808 27398 5817
rect 27342 5743 27344 5752
rect 27396 5743 27398 5752
rect 27344 5714 27396 5720
rect 27448 5681 27476 5850
rect 27434 5672 27490 5681
rect 27434 5607 27490 5616
rect 27436 5568 27488 5574
rect 27436 5510 27488 5516
rect 27344 5160 27396 5166
rect 27344 5102 27396 5108
rect 27356 4321 27384 5102
rect 27448 4622 27476 5510
rect 27540 5137 27568 6072
rect 27632 5545 27660 6326
rect 27618 5536 27674 5545
rect 27618 5471 27674 5480
rect 27526 5128 27582 5137
rect 27526 5063 27582 5072
rect 27712 5024 27764 5030
rect 27618 4992 27674 5001
rect 27712 4966 27764 4972
rect 27618 4927 27674 4936
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 27528 4548 27580 4554
rect 27528 4490 27580 4496
rect 27342 4312 27398 4321
rect 27342 4247 27398 4256
rect 27436 3596 27488 3602
rect 27436 3538 27488 3544
rect 27252 3460 27304 3466
rect 27252 3402 27304 3408
rect 27448 3194 27476 3538
rect 27436 3188 27488 3194
rect 27436 3130 27488 3136
rect 27344 3052 27396 3058
rect 27344 2994 27396 3000
rect 27356 2961 27384 2994
rect 27342 2952 27398 2961
rect 27342 2887 27398 2896
rect 27160 2644 27212 2650
rect 27160 2586 27212 2592
rect 27540 1970 27568 4490
rect 27632 4486 27660 4927
rect 27620 4480 27672 4486
rect 27620 4422 27672 4428
rect 27724 4282 27752 4966
rect 27712 4276 27764 4282
rect 27712 4218 27764 4224
rect 27816 4162 27844 8434
rect 27908 7410 27936 9386
rect 27896 7404 27948 7410
rect 27896 7346 27948 7352
rect 27894 5536 27950 5545
rect 27894 5471 27950 5480
rect 27908 5234 27936 5471
rect 27896 5228 27948 5234
rect 27896 5170 27948 5176
rect 27896 5092 27948 5098
rect 27896 5034 27948 5040
rect 27724 4134 27844 4162
rect 27724 3738 27752 4134
rect 27908 3942 27936 5034
rect 28000 4826 28028 9998
rect 28092 9654 28120 10610
rect 28264 10464 28316 10470
rect 28264 10406 28316 10412
rect 28080 9648 28132 9654
rect 28080 9590 28132 9596
rect 28080 8968 28132 8974
rect 28080 8910 28132 8916
rect 28092 8294 28120 8910
rect 28276 8906 28304 10406
rect 28264 8900 28316 8906
rect 28264 8842 28316 8848
rect 28172 8832 28224 8838
rect 28172 8774 28224 8780
rect 28080 8288 28132 8294
rect 28080 8230 28132 8236
rect 28080 5568 28132 5574
rect 28080 5510 28132 5516
rect 27988 4820 28040 4826
rect 27988 4762 28040 4768
rect 27988 4616 28040 4622
rect 27986 4584 27988 4593
rect 28040 4584 28042 4593
rect 27986 4519 28042 4528
rect 28092 4146 28120 5510
rect 28184 4690 28212 8774
rect 28264 8288 28316 8294
rect 28264 8230 28316 8236
rect 28276 7478 28304 8230
rect 28264 7472 28316 7478
rect 28264 7414 28316 7420
rect 28368 7342 28396 11494
rect 28448 11144 28500 11150
rect 28448 11086 28500 11092
rect 28460 10810 28488 11086
rect 28448 10804 28500 10810
rect 28448 10746 28500 10752
rect 28448 9580 28500 9586
rect 28448 9522 28500 9528
rect 28460 8537 28488 9522
rect 28446 8528 28502 8537
rect 28552 8498 28580 12406
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 31024 12232 31076 12238
rect 31024 12174 31076 12180
rect 28644 11762 28672 12174
rect 30012 12164 30064 12170
rect 30012 12106 30064 12112
rect 28908 12096 28960 12102
rect 28908 12038 28960 12044
rect 28814 11928 28870 11937
rect 28920 11898 28948 12038
rect 28814 11863 28870 11872
rect 28908 11892 28960 11898
rect 28632 11756 28684 11762
rect 28632 11698 28684 11704
rect 28724 11688 28776 11694
rect 28724 11630 28776 11636
rect 28736 10010 28764 11630
rect 28828 11354 28856 11863
rect 28908 11834 28960 11840
rect 30024 11830 30052 12106
rect 30564 12096 30616 12102
rect 30564 12038 30616 12044
rect 30576 11830 30604 12038
rect 30012 11824 30064 11830
rect 30012 11766 30064 11772
rect 30564 11824 30616 11830
rect 30564 11766 30616 11772
rect 29092 11756 29144 11762
rect 29092 11698 29144 11704
rect 29184 11756 29236 11762
rect 29184 11698 29236 11704
rect 30472 11756 30524 11762
rect 30472 11698 30524 11704
rect 28908 11620 28960 11626
rect 28908 11562 28960 11568
rect 28816 11348 28868 11354
rect 28816 11290 28868 11296
rect 28816 10600 28868 10606
rect 28814 10568 28816 10577
rect 28868 10568 28870 10577
rect 28814 10503 28870 10512
rect 28736 9982 28856 10010
rect 28724 9920 28776 9926
rect 28724 9862 28776 9868
rect 28632 9512 28684 9518
rect 28632 9454 28684 9460
rect 28644 9178 28672 9454
rect 28632 9172 28684 9178
rect 28632 9114 28684 9120
rect 28446 8463 28502 8472
rect 28540 8492 28592 8498
rect 28540 8434 28592 8440
rect 28448 8424 28500 8430
rect 28448 8366 28500 8372
rect 28460 8129 28488 8366
rect 28446 8120 28502 8129
rect 28446 8055 28502 8064
rect 28356 7336 28408 7342
rect 28262 7304 28318 7313
rect 28356 7278 28408 7284
rect 28262 7239 28318 7248
rect 28276 5030 28304 7239
rect 28460 6361 28488 8055
rect 28552 6866 28580 8434
rect 28540 6860 28592 6866
rect 28540 6802 28592 6808
rect 28552 6769 28580 6802
rect 28538 6760 28594 6769
rect 28538 6695 28594 6704
rect 28446 6352 28502 6361
rect 28446 6287 28502 6296
rect 28630 6352 28686 6361
rect 28630 6287 28686 6296
rect 28354 5264 28410 5273
rect 28354 5199 28410 5208
rect 28368 5166 28396 5199
rect 28356 5160 28408 5166
rect 28356 5102 28408 5108
rect 28264 5024 28316 5030
rect 28460 5012 28488 6287
rect 28540 6112 28592 6118
rect 28540 6054 28592 6060
rect 28552 5234 28580 6054
rect 28540 5228 28592 5234
rect 28540 5170 28592 5176
rect 28264 4966 28316 4972
rect 28368 4984 28488 5012
rect 28172 4684 28224 4690
rect 28172 4626 28224 4632
rect 28264 4616 28316 4622
rect 28264 4558 28316 4564
rect 28276 4214 28304 4558
rect 28264 4208 28316 4214
rect 28264 4150 28316 4156
rect 28080 4140 28132 4146
rect 28080 4082 28132 4088
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 27712 3732 27764 3738
rect 27712 3674 27764 3680
rect 28080 3732 28132 3738
rect 28080 3674 28132 3680
rect 27988 3664 28040 3670
rect 27988 3606 28040 3612
rect 28000 3058 28028 3606
rect 28092 3534 28120 3674
rect 28080 3528 28132 3534
rect 28080 3470 28132 3476
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 28264 2440 28316 2446
rect 28262 2408 28264 2417
rect 28316 2408 28318 2417
rect 28368 2378 28396 4984
rect 28448 4480 28500 4486
rect 28448 4422 28500 4428
rect 28460 3670 28488 4422
rect 28540 4208 28592 4214
rect 28540 4150 28592 4156
rect 28448 3664 28500 3670
rect 28448 3606 28500 3612
rect 28552 3194 28580 4150
rect 28448 3188 28500 3194
rect 28448 3130 28500 3136
rect 28540 3188 28592 3194
rect 28540 3130 28592 3136
rect 28460 2836 28488 3130
rect 28552 2961 28580 3130
rect 28644 2990 28672 6287
rect 28736 4146 28764 9862
rect 28828 9178 28856 9982
rect 28816 9172 28868 9178
rect 28816 9114 28868 9120
rect 28920 7970 28948 11562
rect 29000 10464 29052 10470
rect 29000 10406 29052 10412
rect 29012 9625 29040 10406
rect 28998 9616 29054 9625
rect 28998 9551 29054 9560
rect 29104 8412 29132 11698
rect 29196 11218 29224 11698
rect 29368 11552 29420 11558
rect 29368 11494 29420 11500
rect 30288 11552 30340 11558
rect 30288 11494 30340 11500
rect 29184 11212 29236 11218
rect 29184 11154 29236 11160
rect 28828 7942 28948 7970
rect 29012 8384 29132 8412
rect 28828 7342 28856 7942
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 28920 7546 28948 7822
rect 28908 7540 28960 7546
rect 28908 7482 28960 7488
rect 28816 7336 28868 7342
rect 28816 7278 28868 7284
rect 29012 7274 29040 8384
rect 29092 7744 29144 7750
rect 29092 7686 29144 7692
rect 29000 7268 29052 7274
rect 29000 7210 29052 7216
rect 29012 7002 29040 7210
rect 29000 6996 29052 7002
rect 29000 6938 29052 6944
rect 29104 6866 29132 7686
rect 29092 6860 29144 6866
rect 29092 6802 29144 6808
rect 29000 6316 29052 6322
rect 29000 6258 29052 6264
rect 28908 6248 28960 6254
rect 28908 6190 28960 6196
rect 28920 5710 28948 6190
rect 28908 5704 28960 5710
rect 28908 5646 28960 5652
rect 28816 5160 28868 5166
rect 28816 5102 28868 5108
rect 28724 4140 28776 4146
rect 28724 4082 28776 4088
rect 28724 3528 28776 3534
rect 28722 3496 28724 3505
rect 28776 3496 28778 3505
rect 28722 3431 28778 3440
rect 28736 3233 28764 3431
rect 28722 3224 28778 3233
rect 28722 3159 28778 3168
rect 28724 3120 28776 3126
rect 28724 3062 28776 3068
rect 28632 2984 28684 2990
rect 28538 2952 28594 2961
rect 28632 2926 28684 2932
rect 28538 2887 28594 2896
rect 28736 2836 28764 3062
rect 28460 2808 28764 2836
rect 28828 2650 28856 5102
rect 28906 4992 28962 5001
rect 28906 4927 28962 4936
rect 28920 4690 28948 4927
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 29012 4593 29040 6258
rect 29090 5808 29146 5817
rect 29090 5743 29146 5752
rect 29104 5642 29132 5743
rect 29092 5636 29144 5642
rect 29092 5578 29144 5584
rect 28998 4584 29054 4593
rect 28998 4519 29054 4528
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 28908 4072 28960 4078
rect 28908 4014 28960 4020
rect 28920 3233 28948 4014
rect 28906 3224 28962 3233
rect 28906 3159 28962 3168
rect 29012 2922 29040 4082
rect 29092 4072 29144 4078
rect 29092 4014 29144 4020
rect 29104 3534 29132 4014
rect 29092 3528 29144 3534
rect 29092 3470 29144 3476
rect 29000 2916 29052 2922
rect 29000 2858 29052 2864
rect 29196 2774 29224 11154
rect 29276 10464 29328 10470
rect 29276 10406 29328 10412
rect 29288 7585 29316 10406
rect 29274 7576 29330 7585
rect 29274 7511 29330 7520
rect 29380 6746 29408 11494
rect 30196 11212 30248 11218
rect 30196 11154 30248 11160
rect 29552 11076 29604 11082
rect 29552 11018 29604 11024
rect 29564 10849 29592 11018
rect 29550 10840 29606 10849
rect 29550 10775 29606 10784
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 29564 10130 29592 10406
rect 29552 10124 29604 10130
rect 29552 10066 29604 10072
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 29460 9376 29512 9382
rect 29460 9318 29512 9324
rect 29472 8498 29500 9318
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 29460 8492 29512 8498
rect 29460 8434 29512 8440
rect 29460 8356 29512 8362
rect 29460 8298 29512 8304
rect 29288 6718 29408 6746
rect 29288 5137 29316 6718
rect 29368 6656 29420 6662
rect 29368 6598 29420 6604
rect 29274 5128 29330 5137
rect 29274 5063 29330 5072
rect 29380 4740 29408 6598
rect 29472 6390 29500 8298
rect 29564 6866 29592 8910
rect 29644 8288 29696 8294
rect 29644 8230 29696 8236
rect 29656 7410 29684 8230
rect 29736 7744 29788 7750
rect 29736 7686 29788 7692
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29748 7041 29776 7686
rect 29734 7032 29790 7041
rect 29734 6967 29790 6976
rect 29552 6860 29604 6866
rect 29552 6802 29604 6808
rect 29734 6760 29790 6769
rect 29734 6695 29790 6704
rect 29552 6656 29604 6662
rect 29552 6598 29604 6604
rect 29460 6384 29512 6390
rect 29460 6326 29512 6332
rect 29564 6186 29592 6598
rect 29748 6390 29776 6695
rect 29736 6384 29788 6390
rect 29736 6326 29788 6332
rect 29644 6248 29696 6254
rect 29644 6190 29696 6196
rect 29552 6180 29604 6186
rect 29552 6122 29604 6128
rect 29550 5944 29606 5953
rect 29550 5879 29606 5888
rect 29458 5808 29514 5817
rect 29564 5778 29592 5879
rect 29458 5743 29460 5752
rect 29512 5743 29514 5752
rect 29552 5772 29604 5778
rect 29460 5714 29512 5720
rect 29552 5714 29604 5720
rect 29656 5681 29684 6190
rect 29736 6112 29788 6118
rect 29736 6054 29788 6060
rect 29642 5672 29698 5681
rect 29642 5607 29698 5616
rect 29656 5302 29684 5607
rect 29748 5370 29776 6054
rect 29736 5364 29788 5370
rect 29736 5306 29788 5312
rect 29644 5296 29696 5302
rect 29644 5238 29696 5244
rect 29644 5092 29696 5098
rect 29644 5034 29696 5040
rect 29656 4826 29684 5034
rect 29644 4820 29696 4826
rect 29644 4762 29696 4768
rect 29380 4712 29592 4740
rect 29564 4672 29592 4712
rect 29564 4644 29776 4672
rect 29368 4616 29420 4622
rect 29368 4558 29420 4564
rect 29642 4584 29698 4593
rect 29276 4548 29328 4554
rect 29276 4490 29328 4496
rect 29288 2854 29316 4490
rect 29380 4146 29408 4558
rect 29642 4519 29698 4528
rect 29552 4480 29604 4486
rect 29552 4422 29604 4428
rect 29564 4214 29592 4422
rect 29552 4208 29604 4214
rect 29656 4185 29684 4519
rect 29552 4150 29604 4156
rect 29642 4176 29698 4185
rect 29368 4140 29420 4146
rect 29642 4111 29698 4120
rect 29368 4082 29420 4088
rect 29748 4078 29776 4644
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 29840 3924 29868 9998
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 29920 9172 29972 9178
rect 29920 9114 29972 9120
rect 29932 8634 29960 9114
rect 29920 8628 29972 8634
rect 29920 8570 29972 8576
rect 29920 8424 29972 8430
rect 29920 8366 29972 8372
rect 29932 8090 29960 8366
rect 29920 8084 29972 8090
rect 29920 8026 29972 8032
rect 29918 7168 29974 7177
rect 29918 7103 29974 7112
rect 29932 6254 29960 7103
rect 29920 6248 29972 6254
rect 29920 6190 29972 6196
rect 29932 6089 29960 6190
rect 29918 6080 29974 6089
rect 29918 6015 29974 6024
rect 29920 5772 29972 5778
rect 29920 5714 29972 5720
rect 29932 4622 29960 5714
rect 29920 4616 29972 4622
rect 29920 4558 29972 4564
rect 29920 3936 29972 3942
rect 29840 3896 29920 3924
rect 29920 3878 29972 3884
rect 29552 3732 29604 3738
rect 29552 3674 29604 3680
rect 29458 3632 29514 3641
rect 29368 3596 29420 3602
rect 29458 3567 29514 3576
rect 29368 3538 29420 3544
rect 29276 2848 29328 2854
rect 29276 2790 29328 2796
rect 29012 2746 29224 2774
rect 28816 2644 28868 2650
rect 28816 2586 28868 2592
rect 28262 2343 28318 2352
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 27528 1964 27580 1970
rect 27528 1906 27580 1912
rect 27710 1592 27766 1601
rect 27710 1527 27766 1536
rect 27724 800 27752 1527
rect 28354 1456 28410 1465
rect 28354 1391 28410 1400
rect 28368 800 28396 1391
rect 29012 800 29040 2746
rect 29380 1465 29408 3538
rect 29472 3398 29500 3567
rect 29460 3392 29512 3398
rect 29460 3334 29512 3340
rect 29564 3126 29592 3674
rect 29918 3360 29974 3369
rect 29918 3295 29974 3304
rect 29552 3120 29604 3126
rect 29552 3062 29604 3068
rect 29932 2990 29960 3295
rect 30024 3126 30052 9862
rect 30208 9602 30236 11154
rect 30116 9574 30236 9602
rect 30116 9518 30144 9574
rect 30104 9512 30156 9518
rect 30104 9454 30156 9460
rect 30196 9512 30248 9518
rect 30196 9454 30248 9460
rect 30208 9382 30236 9454
rect 30196 9376 30248 9382
rect 30196 9318 30248 9324
rect 30104 8628 30156 8634
rect 30104 8570 30156 8576
rect 30116 7546 30144 8570
rect 30208 8566 30236 9318
rect 30300 9042 30328 11494
rect 30484 11121 30512 11698
rect 30470 11112 30526 11121
rect 30470 11047 30526 11056
rect 30472 10600 30524 10606
rect 30472 10542 30524 10548
rect 30484 10441 30512 10542
rect 30470 10432 30526 10441
rect 30470 10367 30526 10376
rect 30380 10260 30432 10266
rect 30380 10202 30432 10208
rect 30392 10169 30420 10202
rect 30378 10160 30434 10169
rect 30576 10146 30604 11766
rect 31036 11762 31064 12174
rect 32128 11892 32180 11898
rect 32128 11834 32180 11840
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 30656 11688 30708 11694
rect 30656 11630 30708 11636
rect 30378 10095 30434 10104
rect 30484 10118 30604 10146
rect 30288 9036 30340 9042
rect 30288 8978 30340 8984
rect 30196 8560 30248 8566
rect 30196 8502 30248 8508
rect 30484 8344 30512 10118
rect 30564 9920 30616 9926
rect 30562 9888 30564 9897
rect 30616 9888 30618 9897
rect 30562 9823 30618 9832
rect 30564 8968 30616 8974
rect 30564 8910 30616 8916
rect 30208 8316 30512 8344
rect 30104 7540 30156 7546
rect 30104 7482 30156 7488
rect 30102 7440 30158 7449
rect 30102 7375 30158 7384
rect 30116 6458 30144 7375
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 30102 5128 30158 5137
rect 30102 5063 30158 5072
rect 30116 3942 30144 5063
rect 30208 4826 30236 8316
rect 30576 8276 30604 8910
rect 30668 8634 30696 11630
rect 30748 11076 30800 11082
rect 30748 11018 30800 11024
rect 30760 9586 30788 11018
rect 30748 9580 30800 9586
rect 30748 9522 30800 9528
rect 30840 9376 30892 9382
rect 30840 9318 30892 9324
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 30392 8248 30604 8276
rect 30288 7812 30340 7818
rect 30288 7754 30340 7760
rect 30300 6934 30328 7754
rect 30392 7177 30420 8248
rect 30562 7984 30618 7993
rect 30562 7919 30618 7928
rect 30472 7880 30524 7886
rect 30470 7848 30472 7857
rect 30524 7848 30526 7857
rect 30470 7783 30526 7792
rect 30472 7336 30524 7342
rect 30472 7278 30524 7284
rect 30378 7168 30434 7177
rect 30378 7103 30434 7112
rect 30288 6928 30340 6934
rect 30288 6870 30340 6876
rect 30380 6928 30432 6934
rect 30380 6870 30432 6876
rect 30392 6662 30420 6870
rect 30380 6656 30432 6662
rect 30380 6598 30432 6604
rect 30392 6458 30420 6598
rect 30380 6452 30432 6458
rect 30380 6394 30432 6400
rect 30288 6384 30340 6390
rect 30288 6326 30340 6332
rect 30300 5370 30328 6326
rect 30380 6112 30432 6118
rect 30380 6054 30432 6060
rect 30288 5364 30340 5370
rect 30288 5306 30340 5312
rect 30196 4820 30248 4826
rect 30196 4762 30248 4768
rect 30208 4010 30236 4762
rect 30288 4616 30340 4622
rect 30288 4558 30340 4564
rect 30196 4004 30248 4010
rect 30196 3946 30248 3952
rect 30104 3936 30156 3942
rect 30104 3878 30156 3884
rect 30104 3596 30156 3602
rect 30104 3538 30156 3544
rect 30116 3126 30144 3538
rect 30012 3120 30064 3126
rect 30012 3062 30064 3068
rect 30104 3120 30156 3126
rect 30104 3062 30156 3068
rect 29920 2984 29972 2990
rect 29920 2926 29972 2932
rect 30300 2854 30328 4558
rect 30392 3670 30420 6054
rect 30484 5914 30512 7278
rect 30472 5908 30524 5914
rect 30472 5850 30524 5856
rect 30576 5250 30604 7919
rect 30656 7880 30708 7886
rect 30656 7822 30708 7828
rect 30668 7206 30696 7822
rect 30656 7200 30708 7206
rect 30656 7142 30708 7148
rect 30746 6896 30802 6905
rect 30746 6831 30802 6840
rect 30656 6656 30708 6662
rect 30656 6598 30708 6604
rect 30484 5222 30604 5250
rect 30484 5030 30512 5222
rect 30472 5024 30524 5030
rect 30472 4966 30524 4972
rect 30564 4820 30616 4826
rect 30564 4762 30616 4768
rect 30472 4684 30524 4690
rect 30472 4626 30524 4632
rect 30484 4486 30512 4626
rect 30472 4480 30524 4486
rect 30472 4422 30524 4428
rect 30380 3664 30432 3670
rect 30380 3606 30432 3612
rect 30380 3460 30432 3466
rect 30380 3402 30432 3408
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 30196 2508 30248 2514
rect 30196 2450 30248 2456
rect 29366 1456 29422 1465
rect 29366 1391 29422 1400
rect 30208 1170 30236 2450
rect 30392 2446 30420 3402
rect 30484 2854 30512 4422
rect 30576 3126 30604 4762
rect 30668 3602 30696 6598
rect 30760 4690 30788 6831
rect 30852 5352 30880 9318
rect 30932 8900 30984 8906
rect 30932 8842 30984 8848
rect 30944 8362 30972 8842
rect 30932 8356 30984 8362
rect 30932 8298 30984 8304
rect 31036 8294 31064 11698
rect 31392 11144 31444 11150
rect 31392 11086 31444 11092
rect 31404 10538 31432 11086
rect 31392 10532 31444 10538
rect 31392 10474 31444 10480
rect 31116 10056 31168 10062
rect 31116 9998 31168 10004
rect 31128 9489 31156 9998
rect 31208 9512 31260 9518
rect 31114 9480 31170 9489
rect 31208 9454 31260 9460
rect 31114 9415 31170 9424
rect 31116 8832 31168 8838
rect 31116 8774 31168 8780
rect 31024 8288 31076 8294
rect 31024 8230 31076 8236
rect 31128 8090 31156 8774
rect 31116 8084 31168 8090
rect 31116 8026 31168 8032
rect 31116 7880 31168 7886
rect 31116 7822 31168 7828
rect 31024 7744 31076 7750
rect 30944 7704 31024 7732
rect 30944 7546 30972 7704
rect 31024 7686 31076 7692
rect 31128 7562 31156 7822
rect 31036 7546 31156 7562
rect 30932 7540 30984 7546
rect 30932 7482 30984 7488
rect 31024 7540 31156 7546
rect 31076 7534 31156 7540
rect 31024 7482 31076 7488
rect 30944 6730 30972 7482
rect 31024 7336 31076 7342
rect 31024 7278 31076 7284
rect 30932 6724 30984 6730
rect 30932 6666 30984 6672
rect 30930 6624 30986 6633
rect 30930 6559 30986 6568
rect 30944 6322 30972 6559
rect 30932 6316 30984 6322
rect 30932 6258 30984 6264
rect 30932 5772 30984 5778
rect 31036 5760 31064 7278
rect 30984 5732 31064 5760
rect 30932 5714 30984 5720
rect 30852 5324 31064 5352
rect 30838 5264 30894 5273
rect 30838 5199 30894 5208
rect 30748 4684 30800 4690
rect 30748 4626 30800 4632
rect 30748 4548 30800 4554
rect 30748 4490 30800 4496
rect 30760 4078 30788 4490
rect 30852 4146 30880 5199
rect 30840 4140 30892 4146
rect 30840 4082 30892 4088
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 30748 4072 30800 4078
rect 30748 4014 30800 4020
rect 30944 3913 30972 4082
rect 30930 3904 30986 3913
rect 30930 3839 30986 3848
rect 30930 3768 30986 3777
rect 30930 3703 30986 3712
rect 30656 3596 30708 3602
rect 30656 3538 30708 3544
rect 30840 3392 30892 3398
rect 30840 3334 30892 3340
rect 30852 3194 30880 3334
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 30564 3120 30616 3126
rect 30564 3062 30616 3068
rect 30760 2961 30788 3130
rect 30944 3126 30972 3703
rect 30932 3120 30984 3126
rect 30932 3062 30984 3068
rect 31036 3058 31064 5324
rect 31128 3534 31156 7534
rect 31220 4826 31248 9454
rect 31298 9208 31354 9217
rect 31298 9143 31354 9152
rect 31312 8566 31340 9143
rect 31300 8560 31352 8566
rect 31300 8502 31352 8508
rect 31300 8288 31352 8294
rect 31300 8230 31352 8236
rect 31312 7041 31340 8230
rect 31298 7032 31354 7041
rect 31298 6967 31354 6976
rect 31300 6656 31352 6662
rect 31300 6598 31352 6604
rect 31312 6458 31340 6598
rect 31300 6452 31352 6458
rect 31300 6394 31352 6400
rect 31312 5302 31340 6394
rect 31300 5296 31352 5302
rect 31300 5238 31352 5244
rect 31208 4820 31260 4826
rect 31208 4762 31260 4768
rect 31208 4684 31260 4690
rect 31208 4626 31260 4632
rect 31220 3777 31248 4626
rect 31206 3768 31262 3777
rect 31312 3738 31340 5238
rect 31404 4026 31432 10474
rect 31484 10464 31536 10470
rect 31484 10406 31536 10412
rect 31576 10464 31628 10470
rect 31576 10406 31628 10412
rect 31496 10198 31524 10406
rect 31484 10192 31536 10198
rect 31484 10134 31536 10140
rect 31588 9625 31616 10406
rect 31944 10056 31996 10062
rect 31944 9998 31996 10004
rect 31852 9920 31904 9926
rect 31852 9862 31904 9868
rect 31668 9648 31720 9654
rect 31574 9616 31630 9625
rect 31668 9590 31720 9596
rect 31574 9551 31630 9560
rect 31576 9512 31628 9518
rect 31576 9454 31628 9460
rect 31484 9376 31536 9382
rect 31484 9318 31536 9324
rect 31496 4298 31524 9318
rect 31588 9110 31616 9454
rect 31680 9110 31708 9590
rect 31576 9104 31628 9110
rect 31576 9046 31628 9052
rect 31668 9104 31720 9110
rect 31668 9046 31720 9052
rect 31576 8968 31628 8974
rect 31576 8910 31628 8916
rect 31588 7342 31616 8910
rect 31668 8900 31720 8906
rect 31668 8842 31720 8848
rect 31680 7954 31708 8842
rect 31760 8288 31812 8294
rect 31760 8230 31812 8236
rect 31772 8022 31800 8230
rect 31760 8016 31812 8022
rect 31760 7958 31812 7964
rect 31668 7948 31720 7954
rect 31668 7890 31720 7896
rect 31758 7576 31814 7585
rect 31758 7511 31814 7520
rect 31772 7478 31800 7511
rect 31760 7472 31812 7478
rect 31760 7414 31812 7420
rect 31668 7404 31720 7410
rect 31668 7346 31720 7352
rect 31576 7336 31628 7342
rect 31576 7278 31628 7284
rect 31574 7032 31630 7041
rect 31574 6967 31630 6976
rect 31588 5710 31616 6967
rect 31680 6934 31708 7346
rect 31668 6928 31720 6934
rect 31668 6870 31720 6876
rect 31772 6866 31800 7414
rect 31760 6860 31812 6866
rect 31760 6802 31812 6808
rect 31666 6488 31722 6497
rect 31666 6423 31722 6432
rect 31680 5817 31708 6423
rect 31772 6390 31800 6802
rect 31760 6384 31812 6390
rect 31760 6326 31812 6332
rect 31760 6248 31812 6254
rect 31760 6190 31812 6196
rect 31772 6089 31800 6190
rect 31758 6080 31814 6089
rect 31758 6015 31814 6024
rect 31666 5808 31722 5817
rect 31666 5743 31722 5752
rect 31576 5704 31628 5710
rect 31576 5646 31628 5652
rect 31588 4690 31616 5646
rect 31668 5636 31720 5642
rect 31668 5578 31720 5584
rect 31680 5545 31708 5578
rect 31666 5536 31722 5545
rect 31666 5471 31722 5480
rect 31864 4690 31892 9862
rect 31956 9722 31984 9998
rect 31944 9716 31996 9722
rect 31944 9658 31996 9664
rect 32036 8560 32088 8566
rect 32036 8502 32088 8508
rect 31942 8120 31998 8129
rect 31942 8055 31998 8064
rect 31956 7857 31984 8055
rect 31942 7848 31998 7857
rect 31942 7783 31998 7792
rect 31944 7404 31996 7410
rect 31944 7346 31996 7352
rect 31956 7177 31984 7346
rect 31942 7168 31998 7177
rect 31942 7103 31998 7112
rect 32048 6866 32076 8502
rect 32036 6860 32088 6866
rect 32036 6802 32088 6808
rect 32036 6724 32088 6730
rect 32036 6666 32088 6672
rect 31942 6216 31998 6225
rect 31942 6151 31998 6160
rect 31956 5914 31984 6151
rect 31944 5908 31996 5914
rect 31944 5850 31996 5856
rect 32048 5778 32076 6666
rect 32140 6254 32168 11834
rect 33060 11626 33088 37130
rect 33796 36922 33824 37198
rect 33784 36916 33836 36922
rect 33784 36858 33836 36864
rect 35360 36718 35388 39200
rect 35854 37564 36162 37573
rect 35854 37562 35860 37564
rect 35916 37562 35940 37564
rect 35996 37562 36020 37564
rect 36076 37562 36100 37564
rect 36156 37562 36162 37564
rect 35916 37510 35918 37562
rect 36098 37510 36100 37562
rect 35854 37508 35860 37510
rect 35916 37508 35940 37510
rect 35996 37508 36020 37510
rect 36076 37508 36100 37510
rect 36156 37508 36162 37510
rect 35854 37499 36162 37508
rect 37200 37262 37228 39200
rect 39040 37330 39068 39200
rect 40880 37618 40908 39200
rect 40880 37590 41092 37618
rect 39028 37324 39080 37330
rect 39028 37266 39080 37272
rect 41064 37262 41092 37590
rect 37004 37256 37056 37262
rect 37004 37198 37056 37204
rect 37188 37256 37240 37262
rect 37188 37198 37240 37204
rect 39120 37256 39172 37262
rect 39120 37198 39172 37204
rect 40868 37256 40920 37262
rect 40868 37198 40920 37204
rect 41052 37256 41104 37262
rect 41052 37198 41104 37204
rect 36514 37020 36822 37029
rect 36514 37018 36520 37020
rect 36576 37018 36600 37020
rect 36656 37018 36680 37020
rect 36736 37018 36760 37020
rect 36816 37018 36822 37020
rect 36576 36966 36578 37018
rect 36758 36966 36760 37018
rect 36514 36964 36520 36966
rect 36576 36964 36600 36966
rect 36656 36964 36680 36966
rect 36736 36964 36760 36966
rect 36816 36964 36822 36966
rect 36514 36955 36822 36964
rect 37016 36922 37044 37198
rect 37004 36916 37056 36922
rect 37004 36858 37056 36864
rect 35440 36780 35492 36786
rect 35440 36722 35492 36728
rect 35348 36712 35400 36718
rect 35348 36654 35400 36660
rect 33232 36372 33284 36378
rect 33232 36314 33284 36320
rect 33244 11830 33272 36314
rect 34796 26988 34848 26994
rect 34796 26930 34848 26936
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 33232 11824 33284 11830
rect 33232 11766 33284 11772
rect 33336 11762 33364 24142
rect 33876 11824 33928 11830
rect 33876 11766 33928 11772
rect 33324 11756 33376 11762
rect 33324 11698 33376 11704
rect 33232 11688 33284 11694
rect 33232 11630 33284 11636
rect 33048 11620 33100 11626
rect 33048 11562 33100 11568
rect 32588 11212 32640 11218
rect 32588 11154 32640 11160
rect 32404 9580 32456 9586
rect 32404 9522 32456 9528
rect 32312 9376 32364 9382
rect 32312 9318 32364 9324
rect 32218 8664 32274 8673
rect 32218 8599 32220 8608
rect 32272 8599 32274 8608
rect 32220 8570 32272 8576
rect 32220 8492 32272 8498
rect 32220 8434 32272 8440
rect 32232 7546 32260 8434
rect 32220 7540 32272 7546
rect 32220 7482 32272 7488
rect 32218 7440 32274 7449
rect 32218 7375 32220 7384
rect 32272 7375 32274 7384
rect 32220 7346 32272 7352
rect 32218 7168 32274 7177
rect 32218 7103 32274 7112
rect 32128 6248 32180 6254
rect 32128 6190 32180 6196
rect 32232 5896 32260 7103
rect 32140 5868 32260 5896
rect 32036 5772 32088 5778
rect 32036 5714 32088 5720
rect 32034 5536 32090 5545
rect 32034 5471 32090 5480
rect 32048 5166 32076 5471
rect 32140 5234 32168 5868
rect 32220 5704 32272 5710
rect 32220 5646 32272 5652
rect 32128 5228 32180 5234
rect 32128 5170 32180 5176
rect 32036 5160 32088 5166
rect 32088 5108 32168 5114
rect 32036 5102 32168 5108
rect 32048 5086 32168 5102
rect 32232 5098 32260 5646
rect 32036 5024 32088 5030
rect 32036 4966 32088 4972
rect 31576 4684 31628 4690
rect 31576 4626 31628 4632
rect 31852 4684 31904 4690
rect 31852 4626 31904 4632
rect 31944 4684 31996 4690
rect 31944 4626 31996 4632
rect 31956 4570 31984 4626
rect 31680 4554 31800 4570
rect 31680 4548 31812 4554
rect 31680 4542 31760 4548
rect 31680 4486 31708 4542
rect 31760 4490 31812 4496
rect 31864 4542 31984 4570
rect 31668 4480 31720 4486
rect 31668 4422 31720 4428
rect 31496 4270 31708 4298
rect 31404 3998 31616 4026
rect 31392 3936 31444 3942
rect 31392 3878 31444 3884
rect 31206 3703 31262 3712
rect 31300 3732 31352 3738
rect 31300 3674 31352 3680
rect 31208 3596 31260 3602
rect 31208 3538 31260 3544
rect 31116 3528 31168 3534
rect 31116 3470 31168 3476
rect 31024 3052 31076 3058
rect 31024 2994 31076 3000
rect 31220 2990 31248 3538
rect 31312 3058 31340 3674
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 31208 2984 31260 2990
rect 30746 2952 30802 2961
rect 31208 2926 31260 2932
rect 30746 2887 30802 2896
rect 30472 2848 30524 2854
rect 31404 2825 31432 3878
rect 30472 2790 30524 2796
rect 31390 2816 31446 2825
rect 31390 2751 31446 2760
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 31484 2440 31536 2446
rect 31484 2382 31536 2388
rect 30932 2100 30984 2106
rect 30932 2042 30984 2048
rect 30208 1142 30328 1170
rect 29564 870 29684 898
rect 25042 232 25098 241
rect 25042 167 25098 176
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29564 338 29592 870
rect 29656 800 29684 870
rect 30300 800 30328 1142
rect 30944 800 30972 2042
rect 31496 1630 31524 2382
rect 31484 1624 31536 1630
rect 31484 1566 31536 1572
rect 31588 800 31616 3998
rect 31680 3534 31708 4270
rect 31864 4010 31892 4542
rect 31944 4072 31996 4078
rect 31944 4014 31996 4020
rect 31852 4004 31904 4010
rect 31852 3946 31904 3952
rect 31668 3528 31720 3534
rect 31668 3470 31720 3476
rect 31864 2990 31892 3946
rect 31852 2984 31904 2990
rect 31852 2926 31904 2932
rect 31956 1834 31984 4014
rect 32048 3670 32076 4966
rect 32036 3664 32088 3670
rect 32036 3606 32088 3612
rect 32140 3602 32168 5086
rect 32220 5092 32272 5098
rect 32220 5034 32272 5040
rect 32128 3596 32180 3602
rect 32128 3538 32180 3544
rect 32324 3126 32352 9318
rect 32416 9178 32444 9522
rect 32404 9172 32456 9178
rect 32404 9114 32456 9120
rect 32416 8906 32444 9114
rect 32404 8900 32456 8906
rect 32404 8842 32456 8848
rect 32404 8424 32456 8430
rect 32404 8366 32456 8372
rect 32494 8392 32550 8401
rect 32416 7818 32444 8366
rect 32494 8327 32550 8336
rect 32508 8294 32536 8327
rect 32496 8288 32548 8294
rect 32496 8230 32548 8236
rect 32404 7812 32456 7818
rect 32404 7754 32456 7760
rect 32404 7472 32456 7478
rect 32404 7414 32456 7420
rect 32416 7206 32444 7414
rect 32600 7410 32628 11154
rect 33060 11082 33088 11562
rect 33244 11286 33272 11630
rect 33232 11280 33284 11286
rect 33232 11222 33284 11228
rect 33048 11076 33100 11082
rect 33048 11018 33100 11024
rect 32772 10600 32824 10606
rect 32772 10542 32824 10548
rect 32784 9761 32812 10542
rect 32956 10192 33008 10198
rect 32956 10134 33008 10140
rect 32864 9920 32916 9926
rect 32864 9862 32916 9868
rect 32770 9752 32826 9761
rect 32770 9687 32826 9696
rect 32680 9376 32732 9382
rect 32680 9318 32732 9324
rect 32692 8294 32720 9318
rect 32772 9172 32824 9178
rect 32772 9114 32824 9120
rect 32680 8288 32732 8294
rect 32680 8230 32732 8236
rect 32680 7472 32732 7478
rect 32680 7414 32732 7420
rect 32588 7404 32640 7410
rect 32588 7346 32640 7352
rect 32404 7200 32456 7206
rect 32404 7142 32456 7148
rect 32402 7032 32458 7041
rect 32402 6967 32458 6976
rect 32416 5302 32444 6967
rect 32496 6860 32548 6866
rect 32496 6802 32548 6808
rect 32508 5642 32536 6802
rect 32588 6792 32640 6798
rect 32588 6734 32640 6740
rect 32600 6186 32628 6734
rect 32588 6180 32640 6186
rect 32588 6122 32640 6128
rect 32588 5704 32640 5710
rect 32586 5672 32588 5681
rect 32640 5672 32642 5681
rect 32496 5636 32548 5642
rect 32586 5607 32642 5616
rect 32496 5578 32548 5584
rect 32404 5296 32456 5302
rect 32404 5238 32456 5244
rect 32508 4842 32536 5578
rect 32508 4814 32628 4842
rect 32496 4752 32548 4758
rect 32496 4694 32548 4700
rect 32404 4072 32456 4078
rect 32404 4014 32456 4020
rect 32312 3120 32364 3126
rect 32312 3062 32364 3068
rect 32220 2508 32272 2514
rect 32220 2450 32272 2456
rect 31944 1828 31996 1834
rect 31944 1770 31996 1776
rect 32232 800 32260 2450
rect 32416 2038 32444 4014
rect 32508 3942 32536 4694
rect 32600 4554 32628 4814
rect 32588 4548 32640 4554
rect 32588 4490 32640 4496
rect 32496 3936 32548 3942
rect 32496 3878 32548 3884
rect 32588 3596 32640 3602
rect 32588 3538 32640 3544
rect 32600 3040 32628 3538
rect 32692 3466 32720 7414
rect 32784 7342 32812 9114
rect 32876 7478 32904 9862
rect 32968 8378 32996 10134
rect 33060 9042 33088 11018
rect 33140 10464 33192 10470
rect 33140 10406 33192 10412
rect 33048 9036 33100 9042
rect 33048 8978 33100 8984
rect 33152 8945 33180 10406
rect 33244 9625 33272 11222
rect 33416 11144 33468 11150
rect 33416 11086 33468 11092
rect 33322 10976 33378 10985
rect 33322 10911 33378 10920
rect 33336 10810 33364 10911
rect 33324 10804 33376 10810
rect 33324 10746 33376 10752
rect 33428 10690 33456 11086
rect 33888 11082 33916 11766
rect 33968 11756 34020 11762
rect 33968 11698 34020 11704
rect 33980 11150 34008 11698
rect 34808 11150 34836 26930
rect 35348 24132 35400 24138
rect 35348 24074 35400 24080
rect 33968 11144 34020 11150
rect 33968 11086 34020 11092
rect 34520 11144 34572 11150
rect 34520 11086 34572 11092
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 33876 11076 33928 11082
rect 33876 11018 33928 11024
rect 33336 10662 33456 10690
rect 33336 10606 33364 10662
rect 33324 10600 33376 10606
rect 33324 10542 33376 10548
rect 33230 9616 33286 9625
rect 33230 9551 33286 9560
rect 33138 8936 33194 8945
rect 33048 8900 33100 8906
rect 33138 8871 33194 8880
rect 33048 8842 33100 8848
rect 33060 8537 33088 8842
rect 33232 8832 33284 8838
rect 33232 8774 33284 8780
rect 33244 8537 33272 8774
rect 33046 8528 33102 8537
rect 33046 8463 33102 8472
rect 33230 8528 33286 8537
rect 33230 8463 33286 8472
rect 33232 8424 33284 8430
rect 32968 8350 33088 8378
rect 33232 8366 33284 8372
rect 32956 8288 33008 8294
rect 32956 8230 33008 8236
rect 33060 8242 33088 8350
rect 33140 8288 33192 8294
rect 33060 8236 33140 8242
rect 33060 8230 33192 8236
rect 32968 7954 32996 8230
rect 33060 8214 33180 8230
rect 32956 7948 33008 7954
rect 32956 7890 33008 7896
rect 32864 7472 32916 7478
rect 32864 7414 32916 7420
rect 32772 7336 32824 7342
rect 32824 7296 32904 7324
rect 32772 7278 32824 7284
rect 32876 6202 32904 7296
rect 32968 6254 32996 7890
rect 33152 7410 33180 8214
rect 33140 7404 33192 7410
rect 33140 7346 33192 7352
rect 33048 7268 33100 7274
rect 33100 7228 33180 7256
rect 33048 7210 33100 7216
rect 33046 7168 33102 7177
rect 33046 7103 33102 7112
rect 32784 6174 32904 6202
rect 32956 6248 33008 6254
rect 32956 6190 33008 6196
rect 32784 5030 32812 6174
rect 32968 5914 32996 6190
rect 32956 5908 33008 5914
rect 32956 5850 33008 5856
rect 32864 5636 32916 5642
rect 32864 5578 32916 5584
rect 32772 5024 32824 5030
rect 32772 4966 32824 4972
rect 32784 4826 32812 4966
rect 32876 4826 32904 5578
rect 32968 5545 32996 5850
rect 32954 5536 33010 5545
rect 32954 5471 33010 5480
rect 32772 4820 32824 4826
rect 32772 4762 32824 4768
rect 32864 4820 32916 4826
rect 32864 4762 32916 4768
rect 33060 4690 33088 7103
rect 33152 6866 33180 7228
rect 33140 6860 33192 6866
rect 33140 6802 33192 6808
rect 33244 6662 33272 8366
rect 33336 7177 33364 10542
rect 33600 10192 33652 10198
rect 33598 10160 33600 10169
rect 33652 10160 33654 10169
rect 33598 10095 33654 10104
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33428 8401 33456 9998
rect 33690 9208 33746 9217
rect 33690 9143 33746 9152
rect 33508 8832 33560 8838
rect 33508 8774 33560 8780
rect 33414 8392 33470 8401
rect 33414 8327 33470 8336
rect 33416 8016 33468 8022
rect 33416 7958 33468 7964
rect 33428 7449 33456 7958
rect 33414 7440 33470 7449
rect 33414 7375 33470 7384
rect 33322 7168 33378 7177
rect 33322 7103 33378 7112
rect 33324 6792 33376 6798
rect 33324 6734 33376 6740
rect 33232 6656 33284 6662
rect 33232 6598 33284 6604
rect 33140 6112 33192 6118
rect 33140 6054 33192 6060
rect 33152 5302 33180 6054
rect 33336 5370 33364 6734
rect 33416 6248 33468 6254
rect 33416 6190 33468 6196
rect 33428 5710 33456 6190
rect 33416 5704 33468 5710
rect 33416 5646 33468 5652
rect 33324 5364 33376 5370
rect 33324 5306 33376 5312
rect 33140 5296 33192 5302
rect 33140 5238 33192 5244
rect 32864 4684 32916 4690
rect 32864 4626 32916 4632
rect 33048 4684 33100 4690
rect 33048 4626 33100 4632
rect 33232 4684 33284 4690
rect 33232 4626 33284 4632
rect 32680 3460 32732 3466
rect 32680 3402 32732 3408
rect 32772 3120 32824 3126
rect 32772 3062 32824 3068
rect 32680 3052 32732 3058
rect 32600 3012 32680 3040
rect 32680 2994 32732 3000
rect 32784 2961 32812 3062
rect 32770 2952 32826 2961
rect 32770 2887 32826 2896
rect 32404 2032 32456 2038
rect 32404 1974 32456 1980
rect 32876 800 32904 4626
rect 33138 4584 33194 4593
rect 33138 4519 33140 4528
rect 33192 4519 33194 4528
rect 33140 4490 33192 4496
rect 33244 4010 33272 4626
rect 33336 4622 33364 5306
rect 33416 5228 33468 5234
rect 33416 5170 33468 5176
rect 33428 5030 33456 5170
rect 33416 5024 33468 5030
rect 33416 4966 33468 4972
rect 33324 4616 33376 4622
rect 33324 4558 33376 4564
rect 33416 4072 33468 4078
rect 33416 4014 33468 4020
rect 33232 4004 33284 4010
rect 33232 3946 33284 3952
rect 33324 4004 33376 4010
rect 33324 3946 33376 3952
rect 33048 3732 33100 3738
rect 33048 3674 33100 3680
rect 33060 3466 33088 3674
rect 33048 3460 33100 3466
rect 33048 3402 33100 3408
rect 33046 2952 33102 2961
rect 33046 2887 33102 2896
rect 33060 2854 33088 2887
rect 33048 2848 33100 2854
rect 33048 2790 33100 2796
rect 33336 2774 33364 3946
rect 33152 2746 33364 2774
rect 33152 2582 33180 2746
rect 33428 2582 33456 4014
rect 33520 3398 33548 8774
rect 33704 8566 33732 9143
rect 33692 8560 33744 8566
rect 33692 8502 33744 8508
rect 33784 8492 33836 8498
rect 33784 8434 33836 8440
rect 33692 8084 33744 8090
rect 33692 8026 33744 8032
rect 33600 7948 33652 7954
rect 33600 7890 33652 7896
rect 33612 5370 33640 7890
rect 33600 5364 33652 5370
rect 33600 5306 33652 5312
rect 33704 5250 33732 8026
rect 33796 5914 33824 8434
rect 33888 7818 33916 11018
rect 33980 9217 34008 11086
rect 34244 10056 34296 10062
rect 34244 9998 34296 10004
rect 34256 9761 34284 9998
rect 34336 9920 34388 9926
rect 34336 9862 34388 9868
rect 34242 9752 34298 9761
rect 34242 9687 34298 9696
rect 34348 9586 34376 9862
rect 34336 9580 34388 9586
rect 34336 9522 34388 9528
rect 34336 9444 34388 9450
rect 34336 9386 34388 9392
rect 34060 9376 34112 9382
rect 34060 9318 34112 9324
rect 33966 9208 34022 9217
rect 33966 9143 34022 9152
rect 33968 8968 34020 8974
rect 33968 8910 34020 8916
rect 33876 7812 33928 7818
rect 33876 7754 33928 7760
rect 33888 7585 33916 7754
rect 33874 7576 33930 7585
rect 33874 7511 33930 7520
rect 33888 7410 33916 7511
rect 33876 7404 33928 7410
rect 33876 7346 33928 7352
rect 33874 7168 33930 7177
rect 33874 7103 33930 7112
rect 33888 6934 33916 7103
rect 33876 6928 33928 6934
rect 33876 6870 33928 6876
rect 33784 5908 33836 5914
rect 33784 5850 33836 5856
rect 33704 5222 33824 5250
rect 33692 5160 33744 5166
rect 33692 5102 33744 5108
rect 33704 4826 33732 5102
rect 33692 4820 33744 4826
rect 33692 4762 33744 4768
rect 33796 4146 33824 5222
rect 33784 4140 33836 4146
rect 33784 4082 33836 4088
rect 33888 4026 33916 6870
rect 33796 3998 33916 4026
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 33508 3392 33560 3398
rect 33508 3334 33560 3340
rect 33612 2990 33640 3538
rect 33796 2990 33824 3998
rect 33876 3936 33928 3942
rect 33876 3878 33928 3884
rect 33888 3466 33916 3878
rect 33980 3738 34008 8910
rect 34072 4146 34100 9318
rect 34152 8832 34204 8838
rect 34152 8774 34204 8780
rect 34164 6633 34192 8774
rect 34242 8120 34298 8129
rect 34242 8055 34298 8064
rect 34256 7886 34284 8055
rect 34348 7993 34376 9386
rect 34532 9178 34560 11086
rect 35256 11076 35308 11082
rect 35256 11018 35308 11024
rect 34796 10600 34848 10606
rect 34796 10542 34848 10548
rect 34978 10568 35034 10577
rect 34704 9580 34756 9586
rect 34704 9522 34756 9528
rect 34520 9172 34572 9178
rect 34520 9114 34572 9120
rect 34428 9104 34480 9110
rect 34428 9046 34480 9052
rect 34610 9072 34666 9081
rect 34334 7984 34390 7993
rect 34334 7919 34390 7928
rect 34244 7880 34296 7886
rect 34244 7822 34296 7828
rect 34256 6798 34284 7822
rect 34336 7812 34388 7818
rect 34336 7754 34388 7760
rect 34348 7041 34376 7754
rect 34440 7478 34468 9046
rect 34610 9007 34612 9016
rect 34664 9007 34666 9016
rect 34612 8978 34664 8984
rect 34612 8424 34664 8430
rect 34612 8366 34664 8372
rect 34520 7744 34572 7750
rect 34520 7686 34572 7692
rect 34428 7472 34480 7478
rect 34428 7414 34480 7420
rect 34334 7032 34390 7041
rect 34334 6967 34390 6976
rect 34244 6792 34296 6798
rect 34244 6734 34296 6740
rect 34150 6624 34206 6633
rect 34150 6559 34206 6568
rect 34256 5710 34284 6734
rect 34532 6361 34560 7686
rect 34624 7546 34652 8366
rect 34612 7540 34664 7546
rect 34612 7482 34664 7488
rect 34612 6928 34664 6934
rect 34612 6870 34664 6876
rect 34518 6352 34574 6361
rect 34518 6287 34574 6296
rect 34336 6180 34388 6186
rect 34336 6122 34388 6128
rect 34244 5704 34296 5710
rect 34244 5646 34296 5652
rect 34348 5302 34376 6122
rect 34428 5840 34480 5846
rect 34426 5808 34428 5817
rect 34480 5808 34482 5817
rect 34426 5743 34482 5752
rect 34532 5710 34560 6287
rect 34520 5704 34572 5710
rect 34520 5646 34572 5652
rect 34624 5642 34652 6870
rect 34612 5636 34664 5642
rect 34612 5578 34664 5584
rect 34624 5522 34652 5578
rect 34532 5494 34652 5522
rect 34336 5296 34388 5302
rect 34336 5238 34388 5244
rect 34152 5160 34204 5166
rect 34152 5102 34204 5108
rect 34060 4140 34112 4146
rect 34060 4082 34112 4088
rect 33968 3732 34020 3738
rect 33968 3674 34020 3680
rect 33876 3460 33928 3466
rect 33876 3402 33928 3408
rect 33874 3360 33930 3369
rect 33874 3295 33930 3304
rect 33888 3058 33916 3295
rect 33980 3126 34008 3674
rect 34164 3534 34192 5102
rect 34532 4486 34560 5494
rect 34716 5001 34744 9522
rect 34808 8265 34836 10542
rect 34978 10503 34980 10512
rect 35032 10503 35034 10512
rect 34980 10474 35032 10480
rect 34888 10056 34940 10062
rect 34888 9998 34940 10004
rect 34900 9722 34928 9998
rect 34888 9716 34940 9722
rect 34888 9658 34940 9664
rect 34888 9512 34940 9518
rect 34888 9454 34940 9460
rect 34900 9382 34928 9454
rect 34888 9376 34940 9382
rect 34888 9318 34940 9324
rect 34978 9344 35034 9353
rect 34794 8256 34850 8265
rect 34794 8191 34850 8200
rect 34794 7848 34850 7857
rect 34794 7783 34850 7792
rect 34808 7410 34836 7783
rect 34796 7404 34848 7410
rect 34796 7346 34848 7352
rect 34900 7313 34928 9318
rect 34978 9279 35034 9288
rect 34992 9110 35020 9279
rect 35162 9208 35218 9217
rect 35162 9143 35218 9152
rect 34980 9104 35032 9110
rect 34980 9046 35032 9052
rect 34992 7993 35020 9046
rect 35176 8974 35204 9143
rect 35268 8974 35296 11018
rect 35164 8968 35216 8974
rect 35256 8968 35308 8974
rect 35164 8910 35216 8916
rect 35254 8936 35256 8945
rect 35308 8936 35310 8945
rect 35072 8900 35124 8906
rect 35254 8871 35310 8880
rect 35072 8842 35124 8848
rect 35084 8673 35112 8842
rect 35070 8664 35126 8673
rect 35070 8599 35126 8608
rect 35256 8628 35308 8634
rect 35256 8570 35308 8576
rect 35072 8560 35124 8566
rect 35072 8502 35124 8508
rect 34978 7984 35034 7993
rect 34978 7919 35034 7928
rect 34980 7540 35032 7546
rect 35084 7528 35112 8502
rect 35164 8424 35216 8430
rect 35164 8366 35216 8372
rect 35176 8090 35204 8366
rect 35164 8084 35216 8090
rect 35164 8026 35216 8032
rect 35268 7954 35296 8570
rect 35256 7948 35308 7954
rect 35256 7890 35308 7896
rect 35164 7880 35216 7886
rect 35164 7822 35216 7828
rect 35032 7500 35112 7528
rect 34980 7482 35032 7488
rect 34980 7336 35032 7342
rect 34886 7304 34942 7313
rect 34980 7278 35032 7284
rect 34886 7239 34942 7248
rect 34888 6792 34940 6798
rect 34888 6734 34940 6740
rect 34796 6656 34848 6662
rect 34796 6598 34848 6604
rect 34808 5234 34836 6598
rect 34900 6390 34928 6734
rect 34888 6384 34940 6390
rect 34888 6326 34940 6332
rect 34888 6248 34940 6254
rect 34888 6190 34940 6196
rect 34796 5228 34848 5234
rect 34796 5170 34848 5176
rect 34794 5128 34850 5137
rect 34794 5063 34850 5072
rect 34702 4992 34758 5001
rect 34702 4927 34758 4936
rect 34612 4616 34664 4622
rect 34612 4558 34664 4564
rect 34520 4480 34572 4486
rect 34520 4422 34572 4428
rect 34152 3528 34204 3534
rect 34532 3516 34560 4422
rect 34624 3641 34652 4558
rect 34702 4312 34758 4321
rect 34702 4247 34758 4256
rect 34716 3738 34744 4247
rect 34704 3732 34756 3738
rect 34704 3674 34756 3680
rect 34610 3632 34666 3641
rect 34610 3567 34666 3576
rect 34532 3488 34652 3516
rect 34152 3470 34204 3476
rect 34152 3392 34204 3398
rect 34152 3334 34204 3340
rect 33968 3120 34020 3126
rect 33968 3062 34020 3068
rect 33876 3052 33928 3058
rect 33876 2994 33928 3000
rect 33600 2984 33652 2990
rect 33600 2926 33652 2932
rect 33784 2984 33836 2990
rect 33784 2926 33836 2932
rect 34164 2922 34192 3334
rect 34152 2916 34204 2922
rect 34152 2858 34204 2864
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 34532 2650 34560 2790
rect 34624 2774 34652 3488
rect 34624 2746 34744 2774
rect 34520 2644 34572 2650
rect 34520 2586 34572 2592
rect 33140 2576 33192 2582
rect 33140 2518 33192 2524
rect 33416 2576 33468 2582
rect 33416 2518 33468 2524
rect 34716 2514 34744 2746
rect 34704 2508 34756 2514
rect 34704 2450 34756 2456
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 33232 2304 33284 2310
rect 33232 2246 33284 2252
rect 33244 1902 33272 2246
rect 33428 2038 33456 2382
rect 34152 2372 34204 2378
rect 34152 2314 34204 2320
rect 33416 2032 33468 2038
rect 33416 1974 33468 1980
rect 33232 1896 33284 1902
rect 33232 1838 33284 1844
rect 33428 870 33548 898
rect 29552 332 29604 338
rect 29552 274 29604 280
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33428 202 33456 870
rect 33520 800 33548 870
rect 34164 800 34192 2314
rect 34808 800 34836 5063
rect 34900 3534 34928 6190
rect 34992 5846 35020 7278
rect 35072 7200 35124 7206
rect 35072 7142 35124 7148
rect 35084 7002 35112 7142
rect 35072 6996 35124 7002
rect 35072 6938 35124 6944
rect 35176 6934 35204 7822
rect 35256 7540 35308 7546
rect 35256 7482 35308 7488
rect 35164 6928 35216 6934
rect 35164 6870 35216 6876
rect 35268 6798 35296 7482
rect 35360 7410 35388 24074
rect 35452 8566 35480 36722
rect 35854 36476 36162 36485
rect 35854 36474 35860 36476
rect 35916 36474 35940 36476
rect 35996 36474 36020 36476
rect 36076 36474 36100 36476
rect 36156 36474 36162 36476
rect 35916 36422 35918 36474
rect 36098 36422 36100 36474
rect 35854 36420 35860 36422
rect 35916 36420 35940 36422
rect 35996 36420 36020 36422
rect 36076 36420 36100 36422
rect 36156 36420 36162 36422
rect 35854 36411 36162 36420
rect 36514 35932 36822 35941
rect 36514 35930 36520 35932
rect 36576 35930 36600 35932
rect 36656 35930 36680 35932
rect 36736 35930 36760 35932
rect 36816 35930 36822 35932
rect 36576 35878 36578 35930
rect 36758 35878 36760 35930
rect 36514 35876 36520 35878
rect 36576 35876 36600 35878
rect 36656 35876 36680 35878
rect 36736 35876 36760 35878
rect 36816 35876 36822 35878
rect 36514 35867 36822 35876
rect 35854 35388 36162 35397
rect 35854 35386 35860 35388
rect 35916 35386 35940 35388
rect 35996 35386 36020 35388
rect 36076 35386 36100 35388
rect 36156 35386 36162 35388
rect 35916 35334 35918 35386
rect 36098 35334 36100 35386
rect 35854 35332 35860 35334
rect 35916 35332 35940 35334
rect 35996 35332 36020 35334
rect 36076 35332 36100 35334
rect 36156 35332 36162 35334
rect 35854 35323 36162 35332
rect 36514 34844 36822 34853
rect 36514 34842 36520 34844
rect 36576 34842 36600 34844
rect 36656 34842 36680 34844
rect 36736 34842 36760 34844
rect 36816 34842 36822 34844
rect 36576 34790 36578 34842
rect 36758 34790 36760 34842
rect 36514 34788 36520 34790
rect 36576 34788 36600 34790
rect 36656 34788 36680 34790
rect 36736 34788 36760 34790
rect 36816 34788 36822 34790
rect 36514 34779 36822 34788
rect 35854 34300 36162 34309
rect 35854 34298 35860 34300
rect 35916 34298 35940 34300
rect 35996 34298 36020 34300
rect 36076 34298 36100 34300
rect 36156 34298 36162 34300
rect 35916 34246 35918 34298
rect 36098 34246 36100 34298
rect 35854 34244 35860 34246
rect 35916 34244 35940 34246
rect 35996 34244 36020 34246
rect 36076 34244 36100 34246
rect 36156 34244 36162 34246
rect 35854 34235 36162 34244
rect 36514 33756 36822 33765
rect 36514 33754 36520 33756
rect 36576 33754 36600 33756
rect 36656 33754 36680 33756
rect 36736 33754 36760 33756
rect 36816 33754 36822 33756
rect 36576 33702 36578 33754
rect 36758 33702 36760 33754
rect 36514 33700 36520 33702
rect 36576 33700 36600 33702
rect 36656 33700 36680 33702
rect 36736 33700 36760 33702
rect 36816 33700 36822 33702
rect 36514 33691 36822 33700
rect 35854 33212 36162 33221
rect 35854 33210 35860 33212
rect 35916 33210 35940 33212
rect 35996 33210 36020 33212
rect 36076 33210 36100 33212
rect 36156 33210 36162 33212
rect 35916 33158 35918 33210
rect 36098 33158 36100 33210
rect 35854 33156 35860 33158
rect 35916 33156 35940 33158
rect 35996 33156 36020 33158
rect 36076 33156 36100 33158
rect 36156 33156 36162 33158
rect 35854 33147 36162 33156
rect 36514 32668 36822 32677
rect 36514 32666 36520 32668
rect 36576 32666 36600 32668
rect 36656 32666 36680 32668
rect 36736 32666 36760 32668
rect 36816 32666 36822 32668
rect 36576 32614 36578 32666
rect 36758 32614 36760 32666
rect 36514 32612 36520 32614
rect 36576 32612 36600 32614
rect 36656 32612 36680 32614
rect 36736 32612 36760 32614
rect 36816 32612 36822 32614
rect 36514 32603 36822 32612
rect 35854 32124 36162 32133
rect 35854 32122 35860 32124
rect 35916 32122 35940 32124
rect 35996 32122 36020 32124
rect 36076 32122 36100 32124
rect 36156 32122 36162 32124
rect 35916 32070 35918 32122
rect 36098 32070 36100 32122
rect 35854 32068 35860 32070
rect 35916 32068 35940 32070
rect 35996 32068 36020 32070
rect 36076 32068 36100 32070
rect 36156 32068 36162 32070
rect 35854 32059 36162 32068
rect 36514 31580 36822 31589
rect 36514 31578 36520 31580
rect 36576 31578 36600 31580
rect 36656 31578 36680 31580
rect 36736 31578 36760 31580
rect 36816 31578 36822 31580
rect 36576 31526 36578 31578
rect 36758 31526 36760 31578
rect 36514 31524 36520 31526
rect 36576 31524 36600 31526
rect 36656 31524 36680 31526
rect 36736 31524 36760 31526
rect 36816 31524 36822 31526
rect 36514 31515 36822 31524
rect 35854 31036 36162 31045
rect 35854 31034 35860 31036
rect 35916 31034 35940 31036
rect 35996 31034 36020 31036
rect 36076 31034 36100 31036
rect 36156 31034 36162 31036
rect 35916 30982 35918 31034
rect 36098 30982 36100 31034
rect 35854 30980 35860 30982
rect 35916 30980 35940 30982
rect 35996 30980 36020 30982
rect 36076 30980 36100 30982
rect 36156 30980 36162 30982
rect 35854 30971 36162 30980
rect 36514 30492 36822 30501
rect 36514 30490 36520 30492
rect 36576 30490 36600 30492
rect 36656 30490 36680 30492
rect 36736 30490 36760 30492
rect 36816 30490 36822 30492
rect 36576 30438 36578 30490
rect 36758 30438 36760 30490
rect 36514 30436 36520 30438
rect 36576 30436 36600 30438
rect 36656 30436 36680 30438
rect 36736 30436 36760 30438
rect 36816 30436 36822 30438
rect 36514 30427 36822 30436
rect 35854 29948 36162 29957
rect 35854 29946 35860 29948
rect 35916 29946 35940 29948
rect 35996 29946 36020 29948
rect 36076 29946 36100 29948
rect 36156 29946 36162 29948
rect 35916 29894 35918 29946
rect 36098 29894 36100 29946
rect 35854 29892 35860 29894
rect 35916 29892 35940 29894
rect 35996 29892 36020 29894
rect 36076 29892 36100 29894
rect 36156 29892 36162 29894
rect 35854 29883 36162 29892
rect 36514 29404 36822 29413
rect 36514 29402 36520 29404
rect 36576 29402 36600 29404
rect 36656 29402 36680 29404
rect 36736 29402 36760 29404
rect 36816 29402 36822 29404
rect 36576 29350 36578 29402
rect 36758 29350 36760 29402
rect 36514 29348 36520 29350
rect 36576 29348 36600 29350
rect 36656 29348 36680 29350
rect 36736 29348 36760 29350
rect 36816 29348 36822 29350
rect 36514 29339 36822 29348
rect 35854 28860 36162 28869
rect 35854 28858 35860 28860
rect 35916 28858 35940 28860
rect 35996 28858 36020 28860
rect 36076 28858 36100 28860
rect 36156 28858 36162 28860
rect 35916 28806 35918 28858
rect 36098 28806 36100 28858
rect 35854 28804 35860 28806
rect 35916 28804 35940 28806
rect 35996 28804 36020 28806
rect 36076 28804 36100 28806
rect 36156 28804 36162 28806
rect 35854 28795 36162 28804
rect 36514 28316 36822 28325
rect 36514 28314 36520 28316
rect 36576 28314 36600 28316
rect 36656 28314 36680 28316
rect 36736 28314 36760 28316
rect 36816 28314 36822 28316
rect 36576 28262 36578 28314
rect 36758 28262 36760 28314
rect 36514 28260 36520 28262
rect 36576 28260 36600 28262
rect 36656 28260 36680 28262
rect 36736 28260 36760 28262
rect 36816 28260 36822 28262
rect 36514 28251 36822 28260
rect 35854 27772 36162 27781
rect 35854 27770 35860 27772
rect 35916 27770 35940 27772
rect 35996 27770 36020 27772
rect 36076 27770 36100 27772
rect 36156 27770 36162 27772
rect 35916 27718 35918 27770
rect 36098 27718 36100 27770
rect 35854 27716 35860 27718
rect 35916 27716 35940 27718
rect 35996 27716 36020 27718
rect 36076 27716 36100 27718
rect 36156 27716 36162 27718
rect 35854 27707 36162 27716
rect 36514 27228 36822 27237
rect 36514 27226 36520 27228
rect 36576 27226 36600 27228
rect 36656 27226 36680 27228
rect 36736 27226 36760 27228
rect 36816 27226 36822 27228
rect 36576 27174 36578 27226
rect 36758 27174 36760 27226
rect 36514 27172 36520 27174
rect 36576 27172 36600 27174
rect 36656 27172 36680 27174
rect 36736 27172 36760 27174
rect 36816 27172 36822 27174
rect 36514 27163 36822 27172
rect 35854 26684 36162 26693
rect 35854 26682 35860 26684
rect 35916 26682 35940 26684
rect 35996 26682 36020 26684
rect 36076 26682 36100 26684
rect 36156 26682 36162 26684
rect 35916 26630 35918 26682
rect 36098 26630 36100 26682
rect 35854 26628 35860 26630
rect 35916 26628 35940 26630
rect 35996 26628 36020 26630
rect 36076 26628 36100 26630
rect 36156 26628 36162 26630
rect 35854 26619 36162 26628
rect 36514 26140 36822 26149
rect 36514 26138 36520 26140
rect 36576 26138 36600 26140
rect 36656 26138 36680 26140
rect 36736 26138 36760 26140
rect 36816 26138 36822 26140
rect 36576 26086 36578 26138
rect 36758 26086 36760 26138
rect 36514 26084 36520 26086
rect 36576 26084 36600 26086
rect 36656 26084 36680 26086
rect 36736 26084 36760 26086
rect 36816 26084 36822 26086
rect 36514 26075 36822 26084
rect 35854 25596 36162 25605
rect 35854 25594 35860 25596
rect 35916 25594 35940 25596
rect 35996 25594 36020 25596
rect 36076 25594 36100 25596
rect 36156 25594 36162 25596
rect 35916 25542 35918 25594
rect 36098 25542 36100 25594
rect 35854 25540 35860 25542
rect 35916 25540 35940 25542
rect 35996 25540 36020 25542
rect 36076 25540 36100 25542
rect 36156 25540 36162 25542
rect 35854 25531 36162 25540
rect 36514 25052 36822 25061
rect 36514 25050 36520 25052
rect 36576 25050 36600 25052
rect 36656 25050 36680 25052
rect 36736 25050 36760 25052
rect 36816 25050 36822 25052
rect 36576 24998 36578 25050
rect 36758 24998 36760 25050
rect 36514 24996 36520 24998
rect 36576 24996 36600 24998
rect 36656 24996 36680 24998
rect 36736 24996 36760 24998
rect 36816 24996 36822 24998
rect 36514 24987 36822 24996
rect 35854 24508 36162 24517
rect 35854 24506 35860 24508
rect 35916 24506 35940 24508
rect 35996 24506 36020 24508
rect 36076 24506 36100 24508
rect 36156 24506 36162 24508
rect 35916 24454 35918 24506
rect 36098 24454 36100 24506
rect 35854 24452 35860 24454
rect 35916 24452 35940 24454
rect 35996 24452 36020 24454
rect 36076 24452 36100 24454
rect 36156 24452 36162 24454
rect 35854 24443 36162 24452
rect 36514 23964 36822 23973
rect 36514 23962 36520 23964
rect 36576 23962 36600 23964
rect 36656 23962 36680 23964
rect 36736 23962 36760 23964
rect 36816 23962 36822 23964
rect 36576 23910 36578 23962
rect 36758 23910 36760 23962
rect 36514 23908 36520 23910
rect 36576 23908 36600 23910
rect 36656 23908 36680 23910
rect 36736 23908 36760 23910
rect 36816 23908 36822 23910
rect 36514 23899 36822 23908
rect 35854 23420 36162 23429
rect 35854 23418 35860 23420
rect 35916 23418 35940 23420
rect 35996 23418 36020 23420
rect 36076 23418 36100 23420
rect 36156 23418 36162 23420
rect 35916 23366 35918 23418
rect 36098 23366 36100 23418
rect 35854 23364 35860 23366
rect 35916 23364 35940 23366
rect 35996 23364 36020 23366
rect 36076 23364 36100 23366
rect 36156 23364 36162 23366
rect 35854 23355 36162 23364
rect 36514 22876 36822 22885
rect 36514 22874 36520 22876
rect 36576 22874 36600 22876
rect 36656 22874 36680 22876
rect 36736 22874 36760 22876
rect 36816 22874 36822 22876
rect 36576 22822 36578 22874
rect 36758 22822 36760 22874
rect 36514 22820 36520 22822
rect 36576 22820 36600 22822
rect 36656 22820 36680 22822
rect 36736 22820 36760 22822
rect 36816 22820 36822 22822
rect 36514 22811 36822 22820
rect 35854 22332 36162 22341
rect 35854 22330 35860 22332
rect 35916 22330 35940 22332
rect 35996 22330 36020 22332
rect 36076 22330 36100 22332
rect 36156 22330 36162 22332
rect 35916 22278 35918 22330
rect 36098 22278 36100 22330
rect 35854 22276 35860 22278
rect 35916 22276 35940 22278
rect 35996 22276 36020 22278
rect 36076 22276 36100 22278
rect 36156 22276 36162 22278
rect 35854 22267 36162 22276
rect 36514 21788 36822 21797
rect 36514 21786 36520 21788
rect 36576 21786 36600 21788
rect 36656 21786 36680 21788
rect 36736 21786 36760 21788
rect 36816 21786 36822 21788
rect 36576 21734 36578 21786
rect 36758 21734 36760 21786
rect 36514 21732 36520 21734
rect 36576 21732 36600 21734
rect 36656 21732 36680 21734
rect 36736 21732 36760 21734
rect 36816 21732 36822 21734
rect 36514 21723 36822 21732
rect 39132 21418 39160 37198
rect 40880 36922 40908 37198
rect 42720 37194 42748 39200
rect 43352 37256 43404 37262
rect 43352 37198 43404 37204
rect 42708 37188 42760 37194
rect 42708 37130 42760 37136
rect 40868 36916 40920 36922
rect 40868 36858 40920 36864
rect 39120 21412 39172 21418
rect 39120 21354 39172 21360
rect 35854 21244 36162 21253
rect 35854 21242 35860 21244
rect 35916 21242 35940 21244
rect 35996 21242 36020 21244
rect 36076 21242 36100 21244
rect 36156 21242 36162 21244
rect 35916 21190 35918 21242
rect 36098 21190 36100 21242
rect 35854 21188 35860 21190
rect 35916 21188 35940 21190
rect 35996 21188 36020 21190
rect 36076 21188 36100 21190
rect 36156 21188 36162 21190
rect 35854 21179 36162 21188
rect 36514 20700 36822 20709
rect 36514 20698 36520 20700
rect 36576 20698 36600 20700
rect 36656 20698 36680 20700
rect 36736 20698 36760 20700
rect 36816 20698 36822 20700
rect 36576 20646 36578 20698
rect 36758 20646 36760 20698
rect 36514 20644 36520 20646
rect 36576 20644 36600 20646
rect 36656 20644 36680 20646
rect 36736 20644 36760 20646
rect 36816 20644 36822 20646
rect 36514 20635 36822 20644
rect 35854 20156 36162 20165
rect 35854 20154 35860 20156
rect 35916 20154 35940 20156
rect 35996 20154 36020 20156
rect 36076 20154 36100 20156
rect 36156 20154 36162 20156
rect 35916 20102 35918 20154
rect 36098 20102 36100 20154
rect 35854 20100 35860 20102
rect 35916 20100 35940 20102
rect 35996 20100 36020 20102
rect 36076 20100 36100 20102
rect 36156 20100 36162 20102
rect 35854 20091 36162 20100
rect 36514 19612 36822 19621
rect 36514 19610 36520 19612
rect 36576 19610 36600 19612
rect 36656 19610 36680 19612
rect 36736 19610 36760 19612
rect 36816 19610 36822 19612
rect 36576 19558 36578 19610
rect 36758 19558 36760 19610
rect 36514 19556 36520 19558
rect 36576 19556 36600 19558
rect 36656 19556 36680 19558
rect 36736 19556 36760 19558
rect 36816 19556 36822 19558
rect 36514 19547 36822 19556
rect 35854 19068 36162 19077
rect 35854 19066 35860 19068
rect 35916 19066 35940 19068
rect 35996 19066 36020 19068
rect 36076 19066 36100 19068
rect 36156 19066 36162 19068
rect 35916 19014 35918 19066
rect 36098 19014 36100 19066
rect 35854 19012 35860 19014
rect 35916 19012 35940 19014
rect 35996 19012 36020 19014
rect 36076 19012 36100 19014
rect 36156 19012 36162 19014
rect 35854 19003 36162 19012
rect 36514 18524 36822 18533
rect 36514 18522 36520 18524
rect 36576 18522 36600 18524
rect 36656 18522 36680 18524
rect 36736 18522 36760 18524
rect 36816 18522 36822 18524
rect 36576 18470 36578 18522
rect 36758 18470 36760 18522
rect 36514 18468 36520 18470
rect 36576 18468 36600 18470
rect 36656 18468 36680 18470
rect 36736 18468 36760 18470
rect 36816 18468 36822 18470
rect 36514 18459 36822 18468
rect 35854 17980 36162 17989
rect 35854 17978 35860 17980
rect 35916 17978 35940 17980
rect 35996 17978 36020 17980
rect 36076 17978 36100 17980
rect 36156 17978 36162 17980
rect 35916 17926 35918 17978
rect 36098 17926 36100 17978
rect 35854 17924 35860 17926
rect 35916 17924 35940 17926
rect 35996 17924 36020 17926
rect 36076 17924 36100 17926
rect 36156 17924 36162 17926
rect 35854 17915 36162 17924
rect 36514 17436 36822 17445
rect 36514 17434 36520 17436
rect 36576 17434 36600 17436
rect 36656 17434 36680 17436
rect 36736 17434 36760 17436
rect 36816 17434 36822 17436
rect 36576 17382 36578 17434
rect 36758 17382 36760 17434
rect 36514 17380 36520 17382
rect 36576 17380 36600 17382
rect 36656 17380 36680 17382
rect 36736 17380 36760 17382
rect 36816 17380 36822 17382
rect 36514 17371 36822 17380
rect 35854 16892 36162 16901
rect 35854 16890 35860 16892
rect 35916 16890 35940 16892
rect 35996 16890 36020 16892
rect 36076 16890 36100 16892
rect 36156 16890 36162 16892
rect 35916 16838 35918 16890
rect 36098 16838 36100 16890
rect 35854 16836 35860 16838
rect 35916 16836 35940 16838
rect 35996 16836 36020 16838
rect 36076 16836 36100 16838
rect 36156 16836 36162 16838
rect 35854 16827 36162 16836
rect 36514 16348 36822 16357
rect 36514 16346 36520 16348
rect 36576 16346 36600 16348
rect 36656 16346 36680 16348
rect 36736 16346 36760 16348
rect 36816 16346 36822 16348
rect 36576 16294 36578 16346
rect 36758 16294 36760 16346
rect 36514 16292 36520 16294
rect 36576 16292 36600 16294
rect 36656 16292 36680 16294
rect 36736 16292 36760 16294
rect 36816 16292 36822 16294
rect 36514 16283 36822 16292
rect 35854 15804 36162 15813
rect 35854 15802 35860 15804
rect 35916 15802 35940 15804
rect 35996 15802 36020 15804
rect 36076 15802 36100 15804
rect 36156 15802 36162 15804
rect 35916 15750 35918 15802
rect 36098 15750 36100 15802
rect 35854 15748 35860 15750
rect 35916 15748 35940 15750
rect 35996 15748 36020 15750
rect 36076 15748 36100 15750
rect 36156 15748 36162 15750
rect 35854 15739 36162 15748
rect 36514 15260 36822 15269
rect 36514 15258 36520 15260
rect 36576 15258 36600 15260
rect 36656 15258 36680 15260
rect 36736 15258 36760 15260
rect 36816 15258 36822 15260
rect 36576 15206 36578 15258
rect 36758 15206 36760 15258
rect 36514 15204 36520 15206
rect 36576 15204 36600 15206
rect 36656 15204 36680 15206
rect 36736 15204 36760 15206
rect 36816 15204 36822 15206
rect 36514 15195 36822 15204
rect 35854 14716 36162 14725
rect 35854 14714 35860 14716
rect 35916 14714 35940 14716
rect 35996 14714 36020 14716
rect 36076 14714 36100 14716
rect 36156 14714 36162 14716
rect 35916 14662 35918 14714
rect 36098 14662 36100 14714
rect 35854 14660 35860 14662
rect 35916 14660 35940 14662
rect 35996 14660 36020 14662
rect 36076 14660 36100 14662
rect 36156 14660 36162 14662
rect 35854 14651 36162 14660
rect 43364 14550 43392 37198
rect 44560 36666 44588 39200
rect 46400 37194 46428 39200
rect 48240 37346 48268 39200
rect 48148 37318 48268 37346
rect 46480 37256 46532 37262
rect 46480 37198 46532 37204
rect 46388 37188 46440 37194
rect 46388 37130 46440 37136
rect 44732 36712 44784 36718
rect 44560 36660 44732 36666
rect 44560 36654 44784 36660
rect 44560 36638 44772 36654
rect 46492 26926 46520 37198
rect 48148 37194 48176 37318
rect 48228 37256 48280 37262
rect 48228 37198 48280 37204
rect 48136 37188 48188 37194
rect 48136 37130 48188 37136
rect 48240 36922 48268 37198
rect 48228 36916 48280 36922
rect 48228 36858 48280 36864
rect 50080 36718 50108 39200
rect 51920 37618 51948 39200
rect 51920 37590 52132 37618
rect 52104 37262 52132 37590
rect 51908 37256 51960 37262
rect 51908 37198 51960 37204
rect 52092 37256 52144 37262
rect 52092 37198 52144 37204
rect 51920 36922 51948 37198
rect 53760 37194 53788 39200
rect 55600 37346 55628 39200
rect 55600 37318 55720 37346
rect 53840 37256 53892 37262
rect 53840 37198 53892 37204
rect 55588 37256 55640 37262
rect 55588 37198 55640 37204
rect 53748 37188 53800 37194
rect 53748 37130 53800 37136
rect 51908 36916 51960 36922
rect 51908 36858 51960 36864
rect 50160 36780 50212 36786
rect 50160 36722 50212 36728
rect 50068 36712 50120 36718
rect 50068 36654 50120 36660
rect 50172 32434 50200 36722
rect 50160 32428 50212 32434
rect 50160 32370 50212 32376
rect 53852 29646 53880 37198
rect 55600 36922 55628 37198
rect 55692 37194 55720 37318
rect 57440 37194 57468 39200
rect 58808 37256 58860 37262
rect 58808 37198 58860 37204
rect 55680 37188 55732 37194
rect 55680 37130 55732 37136
rect 57428 37188 57480 37194
rect 57428 37130 57480 37136
rect 55588 36916 55640 36922
rect 55588 36858 55640 36864
rect 53840 29640 53892 29646
rect 53840 29582 53892 29588
rect 46480 26920 46532 26926
rect 46480 26862 46532 26868
rect 43352 14544 43404 14550
rect 43352 14486 43404 14492
rect 58820 14482 58848 37198
rect 59280 36854 59308 39200
rect 66574 37564 66882 37573
rect 66574 37562 66580 37564
rect 66636 37562 66660 37564
rect 66716 37562 66740 37564
rect 66796 37562 66820 37564
rect 66876 37562 66882 37564
rect 66636 37510 66638 37562
rect 66818 37510 66820 37562
rect 66574 37508 66580 37510
rect 66636 37508 66660 37510
rect 66716 37508 66740 37510
rect 66796 37508 66820 37510
rect 66876 37508 66882 37510
rect 66574 37499 66882 37508
rect 67234 37020 67542 37029
rect 67234 37018 67240 37020
rect 67296 37018 67320 37020
rect 67376 37018 67400 37020
rect 67456 37018 67480 37020
rect 67536 37018 67542 37020
rect 67296 36966 67298 37018
rect 67478 36966 67480 37018
rect 67234 36964 67240 36966
rect 67296 36964 67320 36966
rect 67376 36964 67400 36966
rect 67456 36964 67480 36966
rect 67536 36964 67542 36966
rect 67234 36955 67542 36964
rect 59268 36848 59320 36854
rect 59268 36790 59320 36796
rect 66574 36476 66882 36485
rect 66574 36474 66580 36476
rect 66636 36474 66660 36476
rect 66716 36474 66740 36476
rect 66796 36474 66820 36476
rect 66876 36474 66882 36476
rect 66636 36422 66638 36474
rect 66818 36422 66820 36474
rect 66574 36420 66580 36422
rect 66636 36420 66660 36422
rect 66716 36420 66740 36422
rect 66796 36420 66820 36422
rect 66876 36420 66882 36422
rect 66574 36411 66882 36420
rect 67234 35932 67542 35941
rect 67234 35930 67240 35932
rect 67296 35930 67320 35932
rect 67376 35930 67400 35932
rect 67456 35930 67480 35932
rect 67536 35930 67542 35932
rect 67296 35878 67298 35930
rect 67478 35878 67480 35930
rect 67234 35876 67240 35878
rect 67296 35876 67320 35878
rect 67376 35876 67400 35878
rect 67456 35876 67480 35878
rect 67536 35876 67542 35878
rect 67234 35867 67542 35876
rect 66574 35388 66882 35397
rect 66574 35386 66580 35388
rect 66636 35386 66660 35388
rect 66716 35386 66740 35388
rect 66796 35386 66820 35388
rect 66876 35386 66882 35388
rect 66636 35334 66638 35386
rect 66818 35334 66820 35386
rect 66574 35332 66580 35334
rect 66636 35332 66660 35334
rect 66716 35332 66740 35334
rect 66796 35332 66820 35334
rect 66876 35332 66882 35334
rect 66574 35323 66882 35332
rect 67234 34844 67542 34853
rect 67234 34842 67240 34844
rect 67296 34842 67320 34844
rect 67376 34842 67400 34844
rect 67456 34842 67480 34844
rect 67536 34842 67542 34844
rect 67296 34790 67298 34842
rect 67478 34790 67480 34842
rect 67234 34788 67240 34790
rect 67296 34788 67320 34790
rect 67376 34788 67400 34790
rect 67456 34788 67480 34790
rect 67536 34788 67542 34790
rect 67234 34779 67542 34788
rect 66574 34300 66882 34309
rect 66574 34298 66580 34300
rect 66636 34298 66660 34300
rect 66716 34298 66740 34300
rect 66796 34298 66820 34300
rect 66876 34298 66882 34300
rect 66636 34246 66638 34298
rect 66818 34246 66820 34298
rect 66574 34244 66580 34246
rect 66636 34244 66660 34246
rect 66716 34244 66740 34246
rect 66796 34244 66820 34246
rect 66876 34244 66882 34246
rect 66574 34235 66882 34244
rect 67234 33756 67542 33765
rect 67234 33754 67240 33756
rect 67296 33754 67320 33756
rect 67376 33754 67400 33756
rect 67456 33754 67480 33756
rect 67536 33754 67542 33756
rect 67296 33702 67298 33754
rect 67478 33702 67480 33754
rect 67234 33700 67240 33702
rect 67296 33700 67320 33702
rect 67376 33700 67400 33702
rect 67456 33700 67480 33702
rect 67536 33700 67542 33702
rect 67234 33691 67542 33700
rect 66574 33212 66882 33221
rect 66574 33210 66580 33212
rect 66636 33210 66660 33212
rect 66716 33210 66740 33212
rect 66796 33210 66820 33212
rect 66876 33210 66882 33212
rect 66636 33158 66638 33210
rect 66818 33158 66820 33210
rect 66574 33156 66580 33158
rect 66636 33156 66660 33158
rect 66716 33156 66740 33158
rect 66796 33156 66820 33158
rect 66876 33156 66882 33158
rect 66574 33147 66882 33156
rect 67234 32668 67542 32677
rect 67234 32666 67240 32668
rect 67296 32666 67320 32668
rect 67376 32666 67400 32668
rect 67456 32666 67480 32668
rect 67536 32666 67542 32668
rect 67296 32614 67298 32666
rect 67478 32614 67480 32666
rect 67234 32612 67240 32614
rect 67296 32612 67320 32614
rect 67376 32612 67400 32614
rect 67456 32612 67480 32614
rect 67536 32612 67542 32614
rect 67234 32603 67542 32612
rect 66574 32124 66882 32133
rect 66574 32122 66580 32124
rect 66636 32122 66660 32124
rect 66716 32122 66740 32124
rect 66796 32122 66820 32124
rect 66876 32122 66882 32124
rect 66636 32070 66638 32122
rect 66818 32070 66820 32122
rect 66574 32068 66580 32070
rect 66636 32068 66660 32070
rect 66716 32068 66740 32070
rect 66796 32068 66820 32070
rect 66876 32068 66882 32070
rect 66574 32059 66882 32068
rect 67234 31580 67542 31589
rect 67234 31578 67240 31580
rect 67296 31578 67320 31580
rect 67376 31578 67400 31580
rect 67456 31578 67480 31580
rect 67536 31578 67542 31580
rect 67296 31526 67298 31578
rect 67478 31526 67480 31578
rect 67234 31524 67240 31526
rect 67296 31524 67320 31526
rect 67376 31524 67400 31526
rect 67456 31524 67480 31526
rect 67536 31524 67542 31526
rect 67234 31515 67542 31524
rect 66574 31036 66882 31045
rect 66574 31034 66580 31036
rect 66636 31034 66660 31036
rect 66716 31034 66740 31036
rect 66796 31034 66820 31036
rect 66876 31034 66882 31036
rect 66636 30982 66638 31034
rect 66818 30982 66820 31034
rect 66574 30980 66580 30982
rect 66636 30980 66660 30982
rect 66716 30980 66740 30982
rect 66796 30980 66820 30982
rect 66876 30980 66882 30982
rect 66574 30971 66882 30980
rect 67234 30492 67542 30501
rect 67234 30490 67240 30492
rect 67296 30490 67320 30492
rect 67376 30490 67400 30492
rect 67456 30490 67480 30492
rect 67536 30490 67542 30492
rect 67296 30438 67298 30490
rect 67478 30438 67480 30490
rect 67234 30436 67240 30438
rect 67296 30436 67320 30438
rect 67376 30436 67400 30438
rect 67456 30436 67480 30438
rect 67536 30436 67542 30438
rect 67234 30427 67542 30436
rect 66574 29948 66882 29957
rect 66574 29946 66580 29948
rect 66636 29946 66660 29948
rect 66716 29946 66740 29948
rect 66796 29946 66820 29948
rect 66876 29946 66882 29948
rect 66636 29894 66638 29946
rect 66818 29894 66820 29946
rect 66574 29892 66580 29894
rect 66636 29892 66660 29894
rect 66716 29892 66740 29894
rect 66796 29892 66820 29894
rect 66876 29892 66882 29894
rect 66574 29883 66882 29892
rect 67234 29404 67542 29413
rect 67234 29402 67240 29404
rect 67296 29402 67320 29404
rect 67376 29402 67400 29404
rect 67456 29402 67480 29404
rect 67536 29402 67542 29404
rect 67296 29350 67298 29402
rect 67478 29350 67480 29402
rect 67234 29348 67240 29350
rect 67296 29348 67320 29350
rect 67376 29348 67400 29350
rect 67456 29348 67480 29350
rect 67536 29348 67542 29350
rect 67234 29339 67542 29348
rect 66574 28860 66882 28869
rect 66574 28858 66580 28860
rect 66636 28858 66660 28860
rect 66716 28858 66740 28860
rect 66796 28858 66820 28860
rect 66876 28858 66882 28860
rect 66636 28806 66638 28858
rect 66818 28806 66820 28858
rect 66574 28804 66580 28806
rect 66636 28804 66660 28806
rect 66716 28804 66740 28806
rect 66796 28804 66820 28806
rect 66876 28804 66882 28806
rect 66574 28795 66882 28804
rect 67234 28316 67542 28325
rect 67234 28314 67240 28316
rect 67296 28314 67320 28316
rect 67376 28314 67400 28316
rect 67456 28314 67480 28316
rect 67536 28314 67542 28316
rect 67296 28262 67298 28314
rect 67478 28262 67480 28314
rect 67234 28260 67240 28262
rect 67296 28260 67320 28262
rect 67376 28260 67400 28262
rect 67456 28260 67480 28262
rect 67536 28260 67542 28262
rect 67234 28251 67542 28260
rect 66574 27772 66882 27781
rect 66574 27770 66580 27772
rect 66636 27770 66660 27772
rect 66716 27770 66740 27772
rect 66796 27770 66820 27772
rect 66876 27770 66882 27772
rect 66636 27718 66638 27770
rect 66818 27718 66820 27770
rect 66574 27716 66580 27718
rect 66636 27716 66660 27718
rect 66716 27716 66740 27718
rect 66796 27716 66820 27718
rect 66876 27716 66882 27718
rect 66574 27707 66882 27716
rect 67234 27228 67542 27237
rect 67234 27226 67240 27228
rect 67296 27226 67320 27228
rect 67376 27226 67400 27228
rect 67456 27226 67480 27228
rect 67536 27226 67542 27228
rect 67296 27174 67298 27226
rect 67478 27174 67480 27226
rect 67234 27172 67240 27174
rect 67296 27172 67320 27174
rect 67376 27172 67400 27174
rect 67456 27172 67480 27174
rect 67536 27172 67542 27174
rect 67234 27163 67542 27172
rect 66574 26684 66882 26693
rect 66574 26682 66580 26684
rect 66636 26682 66660 26684
rect 66716 26682 66740 26684
rect 66796 26682 66820 26684
rect 66876 26682 66882 26684
rect 66636 26630 66638 26682
rect 66818 26630 66820 26682
rect 66574 26628 66580 26630
rect 66636 26628 66660 26630
rect 66716 26628 66740 26630
rect 66796 26628 66820 26630
rect 66876 26628 66882 26630
rect 66574 26619 66882 26628
rect 67234 26140 67542 26149
rect 67234 26138 67240 26140
rect 67296 26138 67320 26140
rect 67376 26138 67400 26140
rect 67456 26138 67480 26140
rect 67536 26138 67542 26140
rect 67296 26086 67298 26138
rect 67478 26086 67480 26138
rect 67234 26084 67240 26086
rect 67296 26084 67320 26086
rect 67376 26084 67400 26086
rect 67456 26084 67480 26086
rect 67536 26084 67542 26086
rect 67234 26075 67542 26084
rect 66574 25596 66882 25605
rect 66574 25594 66580 25596
rect 66636 25594 66660 25596
rect 66716 25594 66740 25596
rect 66796 25594 66820 25596
rect 66876 25594 66882 25596
rect 66636 25542 66638 25594
rect 66818 25542 66820 25594
rect 66574 25540 66580 25542
rect 66636 25540 66660 25542
rect 66716 25540 66740 25542
rect 66796 25540 66820 25542
rect 66876 25540 66882 25542
rect 66574 25531 66882 25540
rect 67234 25052 67542 25061
rect 67234 25050 67240 25052
rect 67296 25050 67320 25052
rect 67376 25050 67400 25052
rect 67456 25050 67480 25052
rect 67536 25050 67542 25052
rect 67296 24998 67298 25050
rect 67478 24998 67480 25050
rect 67234 24996 67240 24998
rect 67296 24996 67320 24998
rect 67376 24996 67400 24998
rect 67456 24996 67480 24998
rect 67536 24996 67542 24998
rect 67234 24987 67542 24996
rect 66574 24508 66882 24517
rect 66574 24506 66580 24508
rect 66636 24506 66660 24508
rect 66716 24506 66740 24508
rect 66796 24506 66820 24508
rect 66876 24506 66882 24508
rect 66636 24454 66638 24506
rect 66818 24454 66820 24506
rect 66574 24452 66580 24454
rect 66636 24452 66660 24454
rect 66716 24452 66740 24454
rect 66796 24452 66820 24454
rect 66876 24452 66882 24454
rect 66574 24443 66882 24452
rect 67234 23964 67542 23973
rect 67234 23962 67240 23964
rect 67296 23962 67320 23964
rect 67376 23962 67400 23964
rect 67456 23962 67480 23964
rect 67536 23962 67542 23964
rect 67296 23910 67298 23962
rect 67478 23910 67480 23962
rect 67234 23908 67240 23910
rect 67296 23908 67320 23910
rect 67376 23908 67400 23910
rect 67456 23908 67480 23910
rect 67536 23908 67542 23910
rect 67234 23899 67542 23908
rect 66574 23420 66882 23429
rect 66574 23418 66580 23420
rect 66636 23418 66660 23420
rect 66716 23418 66740 23420
rect 66796 23418 66820 23420
rect 66876 23418 66882 23420
rect 66636 23366 66638 23418
rect 66818 23366 66820 23418
rect 66574 23364 66580 23366
rect 66636 23364 66660 23366
rect 66716 23364 66740 23366
rect 66796 23364 66820 23366
rect 66876 23364 66882 23366
rect 66574 23355 66882 23364
rect 67234 22876 67542 22885
rect 67234 22874 67240 22876
rect 67296 22874 67320 22876
rect 67376 22874 67400 22876
rect 67456 22874 67480 22876
rect 67536 22874 67542 22876
rect 67296 22822 67298 22874
rect 67478 22822 67480 22874
rect 67234 22820 67240 22822
rect 67296 22820 67320 22822
rect 67376 22820 67400 22822
rect 67456 22820 67480 22822
rect 67536 22820 67542 22822
rect 67234 22811 67542 22820
rect 66574 22332 66882 22341
rect 66574 22330 66580 22332
rect 66636 22330 66660 22332
rect 66716 22330 66740 22332
rect 66796 22330 66820 22332
rect 66876 22330 66882 22332
rect 66636 22278 66638 22330
rect 66818 22278 66820 22330
rect 66574 22276 66580 22278
rect 66636 22276 66660 22278
rect 66716 22276 66740 22278
rect 66796 22276 66820 22278
rect 66876 22276 66882 22278
rect 66574 22267 66882 22276
rect 67234 21788 67542 21797
rect 67234 21786 67240 21788
rect 67296 21786 67320 21788
rect 67376 21786 67400 21788
rect 67456 21786 67480 21788
rect 67536 21786 67542 21788
rect 67296 21734 67298 21786
rect 67478 21734 67480 21786
rect 67234 21732 67240 21734
rect 67296 21732 67320 21734
rect 67376 21732 67400 21734
rect 67456 21732 67480 21734
rect 67536 21732 67542 21734
rect 67234 21723 67542 21732
rect 66574 21244 66882 21253
rect 66574 21242 66580 21244
rect 66636 21242 66660 21244
rect 66716 21242 66740 21244
rect 66796 21242 66820 21244
rect 66876 21242 66882 21244
rect 66636 21190 66638 21242
rect 66818 21190 66820 21242
rect 66574 21188 66580 21190
rect 66636 21188 66660 21190
rect 66716 21188 66740 21190
rect 66796 21188 66820 21190
rect 66876 21188 66882 21190
rect 66574 21179 66882 21188
rect 67234 20700 67542 20709
rect 67234 20698 67240 20700
rect 67296 20698 67320 20700
rect 67376 20698 67400 20700
rect 67456 20698 67480 20700
rect 67536 20698 67542 20700
rect 67296 20646 67298 20698
rect 67478 20646 67480 20698
rect 67234 20644 67240 20646
rect 67296 20644 67320 20646
rect 67376 20644 67400 20646
rect 67456 20644 67480 20646
rect 67536 20644 67542 20646
rect 67234 20635 67542 20644
rect 66574 20156 66882 20165
rect 66574 20154 66580 20156
rect 66636 20154 66660 20156
rect 66716 20154 66740 20156
rect 66796 20154 66820 20156
rect 66876 20154 66882 20156
rect 66636 20102 66638 20154
rect 66818 20102 66820 20154
rect 66574 20100 66580 20102
rect 66636 20100 66660 20102
rect 66716 20100 66740 20102
rect 66796 20100 66820 20102
rect 66876 20100 66882 20102
rect 66574 20091 66882 20100
rect 67234 19612 67542 19621
rect 67234 19610 67240 19612
rect 67296 19610 67320 19612
rect 67376 19610 67400 19612
rect 67456 19610 67480 19612
rect 67536 19610 67542 19612
rect 67296 19558 67298 19610
rect 67478 19558 67480 19610
rect 67234 19556 67240 19558
rect 67296 19556 67320 19558
rect 67376 19556 67400 19558
rect 67456 19556 67480 19558
rect 67536 19556 67542 19558
rect 67234 19547 67542 19556
rect 66574 19068 66882 19077
rect 66574 19066 66580 19068
rect 66636 19066 66660 19068
rect 66716 19066 66740 19068
rect 66796 19066 66820 19068
rect 66876 19066 66882 19068
rect 66636 19014 66638 19066
rect 66818 19014 66820 19066
rect 66574 19012 66580 19014
rect 66636 19012 66660 19014
rect 66716 19012 66740 19014
rect 66796 19012 66820 19014
rect 66876 19012 66882 19014
rect 66574 19003 66882 19012
rect 67234 18524 67542 18533
rect 67234 18522 67240 18524
rect 67296 18522 67320 18524
rect 67376 18522 67400 18524
rect 67456 18522 67480 18524
rect 67536 18522 67542 18524
rect 67296 18470 67298 18522
rect 67478 18470 67480 18522
rect 67234 18468 67240 18470
rect 67296 18468 67320 18470
rect 67376 18468 67400 18470
rect 67456 18468 67480 18470
rect 67536 18468 67542 18470
rect 67234 18459 67542 18468
rect 66574 17980 66882 17989
rect 66574 17978 66580 17980
rect 66636 17978 66660 17980
rect 66716 17978 66740 17980
rect 66796 17978 66820 17980
rect 66876 17978 66882 17980
rect 66636 17926 66638 17978
rect 66818 17926 66820 17978
rect 66574 17924 66580 17926
rect 66636 17924 66660 17926
rect 66716 17924 66740 17926
rect 66796 17924 66820 17926
rect 66876 17924 66882 17926
rect 66574 17915 66882 17924
rect 67234 17436 67542 17445
rect 67234 17434 67240 17436
rect 67296 17434 67320 17436
rect 67376 17434 67400 17436
rect 67456 17434 67480 17436
rect 67536 17434 67542 17436
rect 67296 17382 67298 17434
rect 67478 17382 67480 17434
rect 67234 17380 67240 17382
rect 67296 17380 67320 17382
rect 67376 17380 67400 17382
rect 67456 17380 67480 17382
rect 67536 17380 67542 17382
rect 67234 17371 67542 17380
rect 66574 16892 66882 16901
rect 66574 16890 66580 16892
rect 66636 16890 66660 16892
rect 66716 16890 66740 16892
rect 66796 16890 66820 16892
rect 66876 16890 66882 16892
rect 66636 16838 66638 16890
rect 66818 16838 66820 16890
rect 66574 16836 66580 16838
rect 66636 16836 66660 16838
rect 66716 16836 66740 16838
rect 66796 16836 66820 16838
rect 66876 16836 66882 16838
rect 66574 16827 66882 16836
rect 67234 16348 67542 16357
rect 67234 16346 67240 16348
rect 67296 16346 67320 16348
rect 67376 16346 67400 16348
rect 67456 16346 67480 16348
rect 67536 16346 67542 16348
rect 67296 16294 67298 16346
rect 67478 16294 67480 16346
rect 67234 16292 67240 16294
rect 67296 16292 67320 16294
rect 67376 16292 67400 16294
rect 67456 16292 67480 16294
rect 67536 16292 67542 16294
rect 67234 16283 67542 16292
rect 66574 15804 66882 15813
rect 66574 15802 66580 15804
rect 66636 15802 66660 15804
rect 66716 15802 66740 15804
rect 66796 15802 66820 15804
rect 66876 15802 66882 15804
rect 66636 15750 66638 15802
rect 66818 15750 66820 15802
rect 66574 15748 66580 15750
rect 66636 15748 66660 15750
rect 66716 15748 66740 15750
rect 66796 15748 66820 15750
rect 66876 15748 66882 15750
rect 66574 15739 66882 15748
rect 67234 15260 67542 15269
rect 67234 15258 67240 15260
rect 67296 15258 67320 15260
rect 67376 15258 67400 15260
rect 67456 15258 67480 15260
rect 67536 15258 67542 15260
rect 67296 15206 67298 15258
rect 67478 15206 67480 15258
rect 67234 15204 67240 15206
rect 67296 15204 67320 15206
rect 67376 15204 67400 15206
rect 67456 15204 67480 15206
rect 67536 15204 67542 15206
rect 67234 15195 67542 15204
rect 66574 14716 66882 14725
rect 66574 14714 66580 14716
rect 66636 14714 66660 14716
rect 66716 14714 66740 14716
rect 66796 14714 66820 14716
rect 66876 14714 66882 14716
rect 66636 14662 66638 14714
rect 66818 14662 66820 14714
rect 66574 14660 66580 14662
rect 66636 14660 66660 14662
rect 66716 14660 66740 14662
rect 66796 14660 66820 14662
rect 66876 14660 66882 14662
rect 66574 14651 66882 14660
rect 58808 14476 58860 14482
rect 58808 14418 58860 14424
rect 36514 14172 36822 14181
rect 36514 14170 36520 14172
rect 36576 14170 36600 14172
rect 36656 14170 36680 14172
rect 36736 14170 36760 14172
rect 36816 14170 36822 14172
rect 36576 14118 36578 14170
rect 36758 14118 36760 14170
rect 36514 14116 36520 14118
rect 36576 14116 36600 14118
rect 36656 14116 36680 14118
rect 36736 14116 36760 14118
rect 36816 14116 36822 14118
rect 36514 14107 36822 14116
rect 67234 14172 67542 14181
rect 67234 14170 67240 14172
rect 67296 14170 67320 14172
rect 67376 14170 67400 14172
rect 67456 14170 67480 14172
rect 67536 14170 67542 14172
rect 67296 14118 67298 14170
rect 67478 14118 67480 14170
rect 67234 14116 67240 14118
rect 67296 14116 67320 14118
rect 67376 14116 67400 14118
rect 67456 14116 67480 14118
rect 67536 14116 67542 14118
rect 67234 14107 67542 14116
rect 35854 13628 36162 13637
rect 35854 13626 35860 13628
rect 35916 13626 35940 13628
rect 35996 13626 36020 13628
rect 36076 13626 36100 13628
rect 36156 13626 36162 13628
rect 35916 13574 35918 13626
rect 36098 13574 36100 13626
rect 35854 13572 35860 13574
rect 35916 13572 35940 13574
rect 35996 13572 36020 13574
rect 36076 13572 36100 13574
rect 36156 13572 36162 13574
rect 35854 13563 36162 13572
rect 66574 13628 66882 13637
rect 66574 13626 66580 13628
rect 66636 13626 66660 13628
rect 66716 13626 66740 13628
rect 66796 13626 66820 13628
rect 66876 13626 66882 13628
rect 66636 13574 66638 13626
rect 66818 13574 66820 13626
rect 66574 13572 66580 13574
rect 66636 13572 66660 13574
rect 66716 13572 66740 13574
rect 66796 13572 66820 13574
rect 66876 13572 66882 13574
rect 66574 13563 66882 13572
rect 36514 13084 36822 13093
rect 36514 13082 36520 13084
rect 36576 13082 36600 13084
rect 36656 13082 36680 13084
rect 36736 13082 36760 13084
rect 36816 13082 36822 13084
rect 36576 13030 36578 13082
rect 36758 13030 36760 13082
rect 36514 13028 36520 13030
rect 36576 13028 36600 13030
rect 36656 13028 36680 13030
rect 36736 13028 36760 13030
rect 36816 13028 36822 13030
rect 36514 13019 36822 13028
rect 67234 13084 67542 13093
rect 67234 13082 67240 13084
rect 67296 13082 67320 13084
rect 67376 13082 67400 13084
rect 67456 13082 67480 13084
rect 67536 13082 67542 13084
rect 67296 13030 67298 13082
rect 67478 13030 67480 13082
rect 67234 13028 67240 13030
rect 67296 13028 67320 13030
rect 67376 13028 67400 13030
rect 67456 13028 67480 13030
rect 67536 13028 67542 13030
rect 67234 13019 67542 13028
rect 35854 12540 36162 12549
rect 35854 12538 35860 12540
rect 35916 12538 35940 12540
rect 35996 12538 36020 12540
rect 36076 12538 36100 12540
rect 36156 12538 36162 12540
rect 35916 12486 35918 12538
rect 36098 12486 36100 12538
rect 35854 12484 35860 12486
rect 35916 12484 35940 12486
rect 35996 12484 36020 12486
rect 36076 12484 36100 12486
rect 36156 12484 36162 12486
rect 35854 12475 36162 12484
rect 66574 12540 66882 12549
rect 66574 12538 66580 12540
rect 66636 12538 66660 12540
rect 66716 12538 66740 12540
rect 66796 12538 66820 12540
rect 66876 12538 66882 12540
rect 66636 12486 66638 12538
rect 66818 12486 66820 12538
rect 66574 12484 66580 12486
rect 66636 12484 66660 12486
rect 66716 12484 66740 12486
rect 66796 12484 66820 12486
rect 66876 12484 66882 12486
rect 66574 12475 66882 12484
rect 36514 11996 36822 12005
rect 36514 11994 36520 11996
rect 36576 11994 36600 11996
rect 36656 11994 36680 11996
rect 36736 11994 36760 11996
rect 36816 11994 36822 11996
rect 36576 11942 36578 11994
rect 36758 11942 36760 11994
rect 36514 11940 36520 11942
rect 36576 11940 36600 11942
rect 36656 11940 36680 11942
rect 36736 11940 36760 11942
rect 36816 11940 36822 11942
rect 36514 11931 36822 11940
rect 67234 11996 67542 12005
rect 67234 11994 67240 11996
rect 67296 11994 67320 11996
rect 67376 11994 67400 11996
rect 67456 11994 67480 11996
rect 67536 11994 67542 11996
rect 67296 11942 67298 11994
rect 67478 11942 67480 11994
rect 67234 11940 67240 11942
rect 67296 11940 67320 11942
rect 67376 11940 67400 11942
rect 67456 11940 67480 11942
rect 67536 11940 67542 11942
rect 67234 11931 67542 11940
rect 35624 11552 35676 11558
rect 35624 11494 35676 11500
rect 35532 10600 35584 10606
rect 35532 10542 35584 10548
rect 35440 8560 35492 8566
rect 35440 8502 35492 8508
rect 35544 8401 35572 10542
rect 35636 9654 35664 11494
rect 35854 11452 36162 11461
rect 35854 11450 35860 11452
rect 35916 11450 35940 11452
rect 35996 11450 36020 11452
rect 36076 11450 36100 11452
rect 36156 11450 36162 11452
rect 35916 11398 35918 11450
rect 36098 11398 36100 11450
rect 35854 11396 35860 11398
rect 35916 11396 35940 11398
rect 35996 11396 36020 11398
rect 36076 11396 36100 11398
rect 36156 11396 36162 11398
rect 35854 11387 36162 11396
rect 66574 11452 66882 11461
rect 66574 11450 66580 11452
rect 66636 11450 66660 11452
rect 66716 11450 66740 11452
rect 66796 11450 66820 11452
rect 66876 11450 66882 11452
rect 66636 11398 66638 11450
rect 66818 11398 66820 11450
rect 66574 11396 66580 11398
rect 66636 11396 66660 11398
rect 66716 11396 66740 11398
rect 66796 11396 66820 11398
rect 66876 11396 66882 11398
rect 66574 11387 66882 11396
rect 38384 11348 38436 11354
rect 38384 11290 38436 11296
rect 35716 11212 35768 11218
rect 35716 11154 35768 11160
rect 35624 9648 35676 9654
rect 35624 9590 35676 9596
rect 35530 8392 35586 8401
rect 35530 8327 35586 8336
rect 35532 8288 35584 8294
rect 35532 8230 35584 8236
rect 35544 7585 35572 8230
rect 35636 7886 35664 9590
rect 35728 8430 35756 11154
rect 37832 11144 37884 11150
rect 37832 11086 37884 11092
rect 36514 10908 36822 10917
rect 36514 10906 36520 10908
rect 36576 10906 36600 10908
rect 36656 10906 36680 10908
rect 36736 10906 36760 10908
rect 36816 10906 36822 10908
rect 36576 10854 36578 10906
rect 36758 10854 36760 10906
rect 36514 10852 36520 10854
rect 36576 10852 36600 10854
rect 36656 10852 36680 10854
rect 36736 10852 36760 10854
rect 36816 10852 36822 10854
rect 36514 10843 36822 10852
rect 35854 10364 36162 10373
rect 35854 10362 35860 10364
rect 35916 10362 35940 10364
rect 35996 10362 36020 10364
rect 36076 10362 36100 10364
rect 36156 10362 36162 10364
rect 35916 10310 35918 10362
rect 36098 10310 36100 10362
rect 35854 10308 35860 10310
rect 35916 10308 35940 10310
rect 35996 10308 36020 10310
rect 36076 10308 36100 10310
rect 36156 10308 36162 10310
rect 35854 10299 36162 10308
rect 36360 10056 36412 10062
rect 36636 10056 36688 10062
rect 36360 9998 36412 10004
rect 36634 10024 36636 10033
rect 37648 10056 37700 10062
rect 36688 10024 36690 10033
rect 35900 9920 35952 9926
rect 35898 9888 35900 9897
rect 35952 9888 35954 9897
rect 35898 9823 35954 9832
rect 36372 9489 36400 9998
rect 37648 9998 37700 10004
rect 36634 9959 36690 9968
rect 36514 9820 36822 9829
rect 36514 9818 36520 9820
rect 36576 9818 36600 9820
rect 36656 9818 36680 9820
rect 36736 9818 36760 9820
rect 36816 9818 36822 9820
rect 36576 9766 36578 9818
rect 36758 9766 36760 9818
rect 36514 9764 36520 9766
rect 36576 9764 36600 9766
rect 36656 9764 36680 9766
rect 36736 9764 36760 9766
rect 36816 9764 36822 9766
rect 36514 9755 36822 9764
rect 37372 9580 37424 9586
rect 37372 9522 37424 9528
rect 36358 9480 36414 9489
rect 36358 9415 36414 9424
rect 37188 9376 37240 9382
rect 37188 9318 37240 9324
rect 35854 9276 36162 9285
rect 35854 9274 35860 9276
rect 35916 9274 35940 9276
rect 35996 9274 36020 9276
rect 36076 9274 36100 9276
rect 36156 9274 36162 9276
rect 35916 9222 35918 9274
rect 36098 9222 36100 9274
rect 35854 9220 35860 9222
rect 35916 9220 35940 9222
rect 35996 9220 36020 9222
rect 36076 9220 36100 9222
rect 36156 9220 36162 9222
rect 35854 9211 36162 9220
rect 35808 9172 35860 9178
rect 35808 9114 35860 9120
rect 35820 8974 35848 9114
rect 36176 9104 36228 9110
rect 36176 9046 36228 9052
rect 35808 8968 35860 8974
rect 35860 8916 35940 8922
rect 35808 8910 35940 8916
rect 35820 8894 35940 8910
rect 35912 8634 35940 8894
rect 35900 8628 35952 8634
rect 35900 8570 35952 8576
rect 35716 8424 35768 8430
rect 35716 8366 35768 8372
rect 36188 8242 36216 9046
rect 36360 8968 36412 8974
rect 36360 8910 36412 8916
rect 37004 8968 37056 8974
rect 37004 8910 37056 8916
rect 36266 8800 36322 8809
rect 36266 8735 36322 8744
rect 36280 8498 36308 8735
rect 36268 8492 36320 8498
rect 36268 8434 36320 8440
rect 36188 8214 36308 8242
rect 35854 8188 36162 8197
rect 35854 8186 35860 8188
rect 35916 8186 35940 8188
rect 35996 8186 36020 8188
rect 36076 8186 36100 8188
rect 36156 8186 36162 8188
rect 35916 8134 35918 8186
rect 36098 8134 36100 8186
rect 35854 8132 35860 8134
rect 35916 8132 35940 8134
rect 35996 8132 36020 8134
rect 36076 8132 36100 8134
rect 36156 8132 36162 8134
rect 35854 8123 36162 8132
rect 35624 7880 35676 7886
rect 35624 7822 35676 7828
rect 35900 7812 35952 7818
rect 35900 7754 35952 7760
rect 35530 7576 35586 7585
rect 35912 7546 35940 7754
rect 35530 7511 35532 7520
rect 35584 7511 35586 7520
rect 35900 7540 35952 7546
rect 35532 7482 35584 7488
rect 35900 7482 35952 7488
rect 35348 7404 35400 7410
rect 35348 7346 35400 7352
rect 35716 7404 35768 7410
rect 35716 7346 35768 7352
rect 35360 7290 35388 7346
rect 35360 7262 35664 7290
rect 35440 7200 35492 7206
rect 35440 7142 35492 7148
rect 35256 6792 35308 6798
rect 35256 6734 35308 6740
rect 35348 6792 35400 6798
rect 35348 6734 35400 6740
rect 35072 6656 35124 6662
rect 35072 6598 35124 6604
rect 34980 5840 35032 5846
rect 34980 5782 35032 5788
rect 35084 5710 35112 6598
rect 35164 6316 35216 6322
rect 35164 6258 35216 6264
rect 35256 6316 35308 6322
rect 35256 6258 35308 6264
rect 35072 5704 35124 5710
rect 35072 5646 35124 5652
rect 35176 5370 35204 6258
rect 35268 6118 35296 6258
rect 35256 6112 35308 6118
rect 35256 6054 35308 6060
rect 35360 5914 35388 6734
rect 35348 5908 35400 5914
rect 35348 5850 35400 5856
rect 35452 5710 35480 7142
rect 35636 6798 35664 7262
rect 35728 6934 35756 7346
rect 35854 7100 36162 7109
rect 35854 7098 35860 7100
rect 35916 7098 35940 7100
rect 35996 7098 36020 7100
rect 36076 7098 36100 7100
rect 36156 7098 36162 7100
rect 35916 7046 35918 7098
rect 36098 7046 36100 7098
rect 35854 7044 35860 7046
rect 35916 7044 35940 7046
rect 35996 7044 36020 7046
rect 36076 7044 36100 7046
rect 36156 7044 36162 7046
rect 35854 7035 36162 7044
rect 35716 6928 35768 6934
rect 35716 6870 35768 6876
rect 35624 6792 35676 6798
rect 35624 6734 35676 6740
rect 35532 6724 35584 6730
rect 35532 6666 35584 6672
rect 35256 5704 35308 5710
rect 35256 5646 35308 5652
rect 35440 5704 35492 5710
rect 35440 5646 35492 5652
rect 35164 5364 35216 5370
rect 35164 5306 35216 5312
rect 35268 5302 35296 5646
rect 35438 5536 35494 5545
rect 35438 5471 35494 5480
rect 35256 5296 35308 5302
rect 35256 5238 35308 5244
rect 35256 4616 35308 4622
rect 34978 4584 35034 4593
rect 35256 4558 35308 4564
rect 34978 4519 35034 4528
rect 34992 3670 35020 4519
rect 35268 4214 35296 4558
rect 35164 4208 35216 4214
rect 35164 4150 35216 4156
rect 35256 4208 35308 4214
rect 35256 4150 35308 4156
rect 34980 3664 35032 3670
rect 34980 3606 35032 3612
rect 34888 3528 34940 3534
rect 34888 3470 34940 3476
rect 35176 3398 35204 4150
rect 35256 4072 35308 4078
rect 35256 4014 35308 4020
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 35268 2446 35296 4014
rect 35452 2774 35480 5471
rect 35544 5234 35572 6666
rect 35636 6254 35664 6734
rect 35716 6316 35768 6322
rect 35716 6258 35768 6264
rect 35624 6248 35676 6254
rect 35624 6190 35676 6196
rect 35624 6112 35676 6118
rect 35728 6089 35756 6258
rect 35624 6054 35676 6060
rect 35714 6080 35770 6089
rect 35532 5228 35584 5234
rect 35532 5170 35584 5176
rect 35636 4706 35664 6054
rect 35714 6015 35770 6024
rect 35854 6012 36162 6021
rect 35854 6010 35860 6012
rect 35916 6010 35940 6012
rect 35996 6010 36020 6012
rect 36076 6010 36100 6012
rect 36156 6010 36162 6012
rect 35916 5958 35918 6010
rect 36098 5958 36100 6010
rect 35854 5956 35860 5958
rect 35916 5956 35940 5958
rect 35996 5956 36020 5958
rect 36076 5956 36100 5958
rect 36156 5956 36162 5958
rect 35854 5947 36162 5956
rect 35714 5808 35770 5817
rect 36280 5794 36308 8214
rect 36372 6866 36400 8910
rect 36912 8832 36964 8838
rect 36912 8774 36964 8780
rect 36514 8732 36822 8741
rect 36514 8730 36520 8732
rect 36576 8730 36600 8732
rect 36656 8730 36680 8732
rect 36736 8730 36760 8732
rect 36816 8730 36822 8732
rect 36576 8678 36578 8730
rect 36758 8678 36760 8730
rect 36514 8676 36520 8678
rect 36576 8676 36600 8678
rect 36656 8676 36680 8678
rect 36736 8676 36760 8678
rect 36816 8676 36822 8678
rect 36514 8667 36822 8676
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 36740 8294 36768 8434
rect 36728 8288 36780 8294
rect 36728 8230 36780 8236
rect 36740 7818 36768 8230
rect 36728 7812 36780 7818
rect 36728 7754 36780 7760
rect 36514 7644 36822 7653
rect 36514 7642 36520 7644
rect 36576 7642 36600 7644
rect 36656 7642 36680 7644
rect 36736 7642 36760 7644
rect 36816 7642 36822 7644
rect 36576 7590 36578 7642
rect 36758 7590 36760 7642
rect 36514 7588 36520 7590
rect 36576 7588 36600 7590
rect 36656 7588 36680 7590
rect 36736 7588 36760 7590
rect 36816 7588 36822 7590
rect 36514 7579 36822 7588
rect 36452 7540 36504 7546
rect 36452 7482 36504 7488
rect 36360 6860 36412 6866
rect 36360 6802 36412 6808
rect 36464 6644 36492 7482
rect 36544 7200 36596 7206
rect 36544 7142 36596 7148
rect 36556 6866 36584 7142
rect 36924 6905 36952 8774
rect 36910 6896 36966 6905
rect 36544 6860 36596 6866
rect 36910 6831 36966 6840
rect 36544 6802 36596 6808
rect 35714 5743 35770 5752
rect 35900 5772 35952 5778
rect 35728 4808 35756 5743
rect 35900 5714 35952 5720
rect 36096 5766 36308 5794
rect 36372 6616 36492 6644
rect 35808 5636 35860 5642
rect 35808 5578 35860 5584
rect 35820 5234 35848 5578
rect 35912 5545 35940 5714
rect 35898 5536 35954 5545
rect 35898 5471 35954 5480
rect 36096 5234 36124 5766
rect 36268 5704 36320 5710
rect 36268 5646 36320 5652
rect 36176 5568 36228 5574
rect 36176 5510 36228 5516
rect 36188 5370 36216 5510
rect 36176 5364 36228 5370
rect 36176 5306 36228 5312
rect 36188 5234 36216 5306
rect 35808 5228 35860 5234
rect 35808 5170 35860 5176
rect 36084 5228 36136 5234
rect 36084 5170 36136 5176
rect 36176 5228 36228 5234
rect 36176 5170 36228 5176
rect 35854 4924 36162 4933
rect 35854 4922 35860 4924
rect 35916 4922 35940 4924
rect 35996 4922 36020 4924
rect 36076 4922 36100 4924
rect 36156 4922 36162 4924
rect 35916 4870 35918 4922
rect 36098 4870 36100 4922
rect 35854 4868 35860 4870
rect 35916 4868 35940 4870
rect 35996 4868 36020 4870
rect 36076 4868 36100 4870
rect 36156 4868 36162 4870
rect 35854 4859 36162 4868
rect 36280 4826 36308 5646
rect 36268 4820 36320 4826
rect 35728 4780 35940 4808
rect 35636 4678 35756 4706
rect 35624 4276 35676 4282
rect 35624 4218 35676 4224
rect 35636 3126 35664 4218
rect 35728 3534 35756 4678
rect 35912 4282 35940 4780
rect 36268 4762 36320 4768
rect 36372 4570 36400 6616
rect 36514 6556 36822 6565
rect 36514 6554 36520 6556
rect 36576 6554 36600 6556
rect 36656 6554 36680 6556
rect 36736 6554 36760 6556
rect 36816 6554 36822 6556
rect 36576 6502 36578 6554
rect 36758 6502 36760 6554
rect 36514 6500 36520 6502
rect 36576 6500 36600 6502
rect 36656 6500 36680 6502
rect 36736 6500 36760 6502
rect 36816 6500 36822 6502
rect 36514 6491 36822 6500
rect 37016 6474 37044 8910
rect 37096 7268 37148 7274
rect 37096 7210 37148 7216
rect 36924 6446 37044 6474
rect 36924 6225 36952 6446
rect 37004 6316 37056 6322
rect 37004 6258 37056 6264
rect 36910 6216 36966 6225
rect 36910 6151 36966 6160
rect 36452 6112 36504 6118
rect 36452 6054 36504 6060
rect 36912 6112 36964 6118
rect 36912 6054 36964 6060
rect 36464 5846 36492 6054
rect 36820 5908 36872 5914
rect 36820 5850 36872 5856
rect 36452 5840 36504 5846
rect 36452 5782 36504 5788
rect 36450 5672 36506 5681
rect 36832 5658 36860 5850
rect 36924 5778 36952 6054
rect 36912 5772 36964 5778
rect 36912 5714 36964 5720
rect 36832 5630 36952 5658
rect 36450 5607 36452 5616
rect 36504 5607 36506 5616
rect 36452 5578 36504 5584
rect 36514 5468 36822 5477
rect 36514 5466 36520 5468
rect 36576 5466 36600 5468
rect 36656 5466 36680 5468
rect 36736 5466 36760 5468
rect 36816 5466 36822 5468
rect 36576 5414 36578 5466
rect 36758 5414 36760 5466
rect 36514 5412 36520 5414
rect 36576 5412 36600 5414
rect 36656 5412 36680 5414
rect 36736 5412 36760 5414
rect 36816 5412 36822 5414
rect 36514 5403 36822 5412
rect 36452 5364 36504 5370
rect 36452 5306 36504 5312
rect 36464 4865 36492 5306
rect 36820 5296 36872 5302
rect 36820 5238 36872 5244
rect 36544 5160 36596 5166
rect 36544 5102 36596 5108
rect 36450 4856 36506 4865
rect 36450 4791 36506 4800
rect 36188 4542 36400 4570
rect 36084 4480 36136 4486
rect 36084 4422 36136 4428
rect 35900 4276 35952 4282
rect 35900 4218 35952 4224
rect 36096 4078 36124 4422
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 36188 3890 36216 4542
rect 36268 4480 36320 4486
rect 36556 4468 36584 5102
rect 36832 4758 36860 5238
rect 36924 5234 36952 5630
rect 37016 5370 37044 6258
rect 37004 5364 37056 5370
rect 37004 5306 37056 5312
rect 36912 5228 36964 5234
rect 36912 5170 36964 5176
rect 36820 4752 36872 4758
rect 36820 4694 36872 4700
rect 37108 4672 37136 7210
rect 36268 4422 36320 4428
rect 36372 4440 36584 4468
rect 36924 4644 37136 4672
rect 36280 4185 36308 4422
rect 36266 4176 36322 4185
rect 36266 4111 36322 4120
rect 36188 3862 36308 3890
rect 35854 3836 36162 3845
rect 35854 3834 35860 3836
rect 35916 3834 35940 3836
rect 35996 3834 36020 3836
rect 36076 3834 36100 3836
rect 36156 3834 36162 3836
rect 35916 3782 35918 3834
rect 36098 3782 36100 3834
rect 35854 3780 35860 3782
rect 35916 3780 35940 3782
rect 35996 3780 36020 3782
rect 36076 3780 36100 3782
rect 36156 3780 36162 3782
rect 35854 3771 36162 3780
rect 36280 3534 36308 3862
rect 35716 3528 35768 3534
rect 35716 3470 35768 3476
rect 36268 3528 36320 3534
rect 36268 3470 36320 3476
rect 35728 3398 35756 3470
rect 35716 3392 35768 3398
rect 35716 3334 35768 3340
rect 36084 3392 36136 3398
rect 36084 3334 36136 3340
rect 36096 3194 36124 3334
rect 36084 3188 36136 3194
rect 36084 3130 36136 3136
rect 35532 3120 35584 3126
rect 35532 3062 35584 3068
rect 35624 3120 35676 3126
rect 35624 3062 35676 3068
rect 35544 2938 35572 3062
rect 35544 2910 35940 2938
rect 35912 2854 35940 2910
rect 35900 2848 35952 2854
rect 35900 2790 35952 2796
rect 36372 2774 36400 4440
rect 36514 4380 36822 4389
rect 36514 4378 36520 4380
rect 36576 4378 36600 4380
rect 36656 4378 36680 4380
rect 36736 4378 36760 4380
rect 36816 4378 36822 4380
rect 36576 4326 36578 4378
rect 36758 4326 36760 4378
rect 36514 4324 36520 4326
rect 36576 4324 36600 4326
rect 36656 4324 36680 4326
rect 36736 4324 36760 4326
rect 36816 4324 36822 4326
rect 36514 4315 36822 4324
rect 36924 4162 36952 4644
rect 36648 4146 36952 4162
rect 36636 4140 36952 4146
rect 36688 4134 36952 4140
rect 36636 4082 36688 4088
rect 36728 4072 36780 4078
rect 36728 4014 36780 4020
rect 36912 4072 36964 4078
rect 36912 4014 36964 4020
rect 36740 3942 36768 4014
rect 36728 3936 36780 3942
rect 36728 3878 36780 3884
rect 36924 3738 36952 4014
rect 36912 3732 36964 3738
rect 36912 3674 36964 3680
rect 37200 3534 37228 9318
rect 37280 8356 37332 8362
rect 37280 8298 37332 8304
rect 37292 7410 37320 8298
rect 37280 7404 37332 7410
rect 37280 7346 37332 7352
rect 37384 6866 37412 9522
rect 37464 8832 37516 8838
rect 37464 8774 37516 8780
rect 37372 6860 37424 6866
rect 37372 6802 37424 6808
rect 37280 5908 37332 5914
rect 37280 5850 37332 5856
rect 37292 5642 37320 5850
rect 37280 5636 37332 5642
rect 37280 5578 37332 5584
rect 37476 5386 37504 8774
rect 37556 8560 37608 8566
rect 37556 8502 37608 8508
rect 37384 5358 37504 5386
rect 37384 5273 37412 5358
rect 37464 5296 37516 5302
rect 37370 5264 37426 5273
rect 37464 5238 37516 5244
rect 37370 5199 37426 5208
rect 37280 5024 37332 5030
rect 37280 4966 37332 4972
rect 37372 5024 37424 5030
rect 37372 4966 37424 4972
rect 37292 4826 37320 4966
rect 37280 4820 37332 4826
rect 37280 4762 37332 4768
rect 37384 4690 37412 4966
rect 37476 4758 37504 5238
rect 37464 4752 37516 4758
rect 37464 4694 37516 4700
rect 37372 4684 37424 4690
rect 37372 4626 37424 4632
rect 37568 4570 37596 8502
rect 37476 4542 37596 4570
rect 37372 4276 37424 4282
rect 37372 4218 37424 4224
rect 37188 3528 37240 3534
rect 37188 3470 37240 3476
rect 37280 3528 37332 3534
rect 37280 3470 37332 3476
rect 37292 3346 37320 3470
rect 36924 3318 37320 3346
rect 36514 3292 36822 3301
rect 36514 3290 36520 3292
rect 36576 3290 36600 3292
rect 36656 3290 36680 3292
rect 36736 3290 36760 3292
rect 36816 3290 36822 3292
rect 36576 3238 36578 3290
rect 36758 3238 36760 3290
rect 36514 3236 36520 3238
rect 36576 3236 36600 3238
rect 36656 3236 36680 3238
rect 36736 3236 36760 3238
rect 36816 3236 36822 3238
rect 36514 3227 36822 3236
rect 35452 2746 35572 2774
rect 35544 2514 35572 2746
rect 35854 2748 36162 2757
rect 35854 2746 35860 2748
rect 35916 2746 35940 2748
rect 35996 2746 36020 2748
rect 36076 2746 36100 2748
rect 36156 2746 36162 2748
rect 35916 2694 35918 2746
rect 36098 2694 36100 2746
rect 35854 2692 35860 2694
rect 35916 2692 35940 2694
rect 35996 2692 36020 2694
rect 36076 2692 36100 2694
rect 36156 2692 36162 2694
rect 35854 2683 36162 2692
rect 36280 2746 36400 2774
rect 36280 2650 36308 2746
rect 36268 2644 36320 2650
rect 36268 2586 36320 2592
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 35532 2508 35584 2514
rect 35532 2450 35584 2456
rect 36084 2508 36136 2514
rect 36084 2450 36136 2456
rect 35256 2440 35308 2446
rect 35256 2382 35308 2388
rect 35438 1320 35494 1329
rect 35438 1255 35494 1264
rect 35452 800 35480 1255
rect 36096 800 36124 2450
rect 36372 2310 36400 2586
rect 36924 2446 36952 3318
rect 37384 2938 37412 4218
rect 37476 4146 37504 4542
rect 37556 4480 37608 4486
rect 37556 4422 37608 4428
rect 37568 4282 37596 4422
rect 37556 4276 37608 4282
rect 37556 4218 37608 4224
rect 37464 4140 37516 4146
rect 37464 4082 37516 4088
rect 37556 4140 37608 4146
rect 37556 4082 37608 4088
rect 37568 4049 37596 4082
rect 37554 4040 37610 4049
rect 37554 3975 37610 3984
rect 37384 2922 37504 2938
rect 37384 2916 37516 2922
rect 37384 2910 37464 2916
rect 37464 2858 37516 2864
rect 36912 2440 36964 2446
rect 36912 2382 36964 2388
rect 36360 2304 36412 2310
rect 36360 2246 36412 2252
rect 36514 2204 36822 2213
rect 36514 2202 36520 2204
rect 36576 2202 36600 2204
rect 36656 2202 36680 2204
rect 36736 2202 36760 2204
rect 36816 2202 36822 2204
rect 36576 2150 36578 2202
rect 36758 2150 36760 2202
rect 36514 2148 36520 2150
rect 36576 2148 36600 2150
rect 36656 2148 36680 2150
rect 36736 2148 36760 2150
rect 36816 2148 36822 2150
rect 36514 2139 36822 2148
rect 37660 1465 37688 9998
rect 37844 9586 37872 11086
rect 37832 9580 37884 9586
rect 37832 9522 37884 9528
rect 37740 9444 37792 9450
rect 37740 9386 37792 9392
rect 37752 9178 37780 9386
rect 37740 9172 37792 9178
rect 37740 9114 37792 9120
rect 37844 8106 37872 9522
rect 38016 9376 38068 9382
rect 38016 9318 38068 9324
rect 38200 9376 38252 9382
rect 38200 9318 38252 9324
rect 37844 8078 37964 8106
rect 37936 7954 37964 8078
rect 37832 7948 37884 7954
rect 37832 7890 37884 7896
rect 37924 7948 37976 7954
rect 37924 7890 37976 7896
rect 37844 6866 37872 7890
rect 37924 7812 37976 7818
rect 37924 7754 37976 7760
rect 37936 7290 37964 7754
rect 38028 7478 38056 9318
rect 38212 9081 38240 9318
rect 38198 9072 38254 9081
rect 38198 9007 38254 9016
rect 38200 8968 38252 8974
rect 38200 8910 38252 8916
rect 38016 7472 38068 7478
rect 38016 7414 38068 7420
rect 37936 7262 38056 7290
rect 37924 7200 37976 7206
rect 37924 7142 37976 7148
rect 37936 7002 37964 7142
rect 37924 6996 37976 7002
rect 37924 6938 37976 6944
rect 37832 6860 37884 6866
rect 37832 6802 37884 6808
rect 37844 6746 37872 6802
rect 37844 6718 37964 6746
rect 37936 6254 37964 6718
rect 37924 6248 37976 6254
rect 37924 6190 37976 6196
rect 37936 5574 37964 6190
rect 37832 5568 37884 5574
rect 37832 5510 37884 5516
rect 37924 5568 37976 5574
rect 37924 5510 37976 5516
rect 37740 5160 37792 5166
rect 37738 5128 37740 5137
rect 37792 5128 37794 5137
rect 37738 5063 37794 5072
rect 37738 4856 37794 4865
rect 37738 4791 37794 4800
rect 37752 4690 37780 4791
rect 37844 4690 37872 5510
rect 37740 4684 37792 4690
rect 37740 4626 37792 4632
rect 37832 4684 37884 4690
rect 37832 4626 37884 4632
rect 37936 4622 37964 5510
rect 37924 4616 37976 4622
rect 37924 4558 37976 4564
rect 37740 4072 37792 4078
rect 37738 4040 37740 4049
rect 37792 4040 37794 4049
rect 37738 3975 37794 3984
rect 37936 3194 37964 4558
rect 37924 3188 37976 3194
rect 37924 3130 37976 3136
rect 38028 3074 38056 7262
rect 38108 7268 38160 7274
rect 38108 7210 38160 7216
rect 38120 4214 38148 7210
rect 38212 6882 38240 8910
rect 38292 7744 38344 7750
rect 38292 7686 38344 7692
rect 38304 7410 38332 7686
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 38212 6854 38332 6882
rect 38200 5228 38252 5234
rect 38200 5170 38252 5176
rect 38212 4865 38240 5170
rect 38198 4856 38254 4865
rect 38198 4791 38254 4800
rect 38108 4208 38160 4214
rect 38108 4150 38160 4156
rect 38200 4208 38252 4214
rect 38200 4150 38252 4156
rect 38108 4072 38160 4078
rect 38108 4014 38160 4020
rect 37752 3046 38056 3074
rect 36726 1456 36782 1465
rect 36726 1391 36782 1400
rect 37646 1456 37702 1465
rect 37646 1391 37702 1400
rect 36740 800 36768 1391
rect 37384 870 37504 898
rect 37384 800 37412 870
rect 33416 196 33468 202
rect 33416 138 33468 144
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 37476 762 37504 870
rect 37752 762 37780 3046
rect 38120 2774 38148 4014
rect 38028 2746 38148 2774
rect 38028 800 38056 2746
rect 38108 2304 38160 2310
rect 38108 2246 38160 2252
rect 38120 2106 38148 2246
rect 38108 2100 38160 2106
rect 38108 2042 38160 2048
rect 38212 1834 38240 4150
rect 38304 1902 38332 6854
rect 38396 4214 38424 11290
rect 67234 10908 67542 10917
rect 67234 10906 67240 10908
rect 67296 10906 67320 10908
rect 67376 10906 67400 10908
rect 67456 10906 67480 10908
rect 67536 10906 67542 10908
rect 67296 10854 67298 10906
rect 67478 10854 67480 10906
rect 67234 10852 67240 10854
rect 67296 10852 67320 10854
rect 67376 10852 67400 10854
rect 67456 10852 67480 10854
rect 67536 10852 67542 10854
rect 67234 10843 67542 10852
rect 66574 10364 66882 10373
rect 66574 10362 66580 10364
rect 66636 10362 66660 10364
rect 66716 10362 66740 10364
rect 66796 10362 66820 10364
rect 66876 10362 66882 10364
rect 66636 10310 66638 10362
rect 66818 10310 66820 10362
rect 66574 10308 66580 10310
rect 66636 10308 66660 10310
rect 66716 10308 66740 10310
rect 66796 10308 66820 10310
rect 66876 10308 66882 10310
rect 66574 10299 66882 10308
rect 67234 9820 67542 9829
rect 67234 9818 67240 9820
rect 67296 9818 67320 9820
rect 67376 9818 67400 9820
rect 67456 9818 67480 9820
rect 67536 9818 67542 9820
rect 67296 9766 67298 9818
rect 67478 9766 67480 9818
rect 67234 9764 67240 9766
rect 67296 9764 67320 9766
rect 67376 9764 67400 9766
rect 67456 9764 67480 9766
rect 67536 9764 67542 9766
rect 67234 9755 67542 9764
rect 40040 9512 40092 9518
rect 40040 9454 40092 9460
rect 38752 9036 38804 9042
rect 38752 8978 38804 8984
rect 38660 8900 38712 8906
rect 38660 8842 38712 8848
rect 38672 5914 38700 8842
rect 38660 5908 38712 5914
rect 38660 5850 38712 5856
rect 38568 4480 38620 4486
rect 38620 4440 38700 4468
rect 38568 4422 38620 4428
rect 38384 4208 38436 4214
rect 38384 4150 38436 4156
rect 38568 4140 38620 4146
rect 38568 4082 38620 4088
rect 38474 3768 38530 3777
rect 38474 3703 38530 3712
rect 38488 3466 38516 3703
rect 38580 3602 38608 4082
rect 38568 3596 38620 3602
rect 38568 3538 38620 3544
rect 38476 3460 38528 3466
rect 38476 3402 38528 3408
rect 38672 3126 38700 4440
rect 38660 3120 38712 3126
rect 38660 3062 38712 3068
rect 38764 2774 38792 8978
rect 39764 8832 39816 8838
rect 39764 8774 39816 8780
rect 39776 8498 39804 8774
rect 39764 8492 39816 8498
rect 39764 8434 39816 8440
rect 39396 8424 39448 8430
rect 39396 8366 39448 8372
rect 39212 8356 39264 8362
rect 39212 8298 39264 8304
rect 39028 8288 39080 8294
rect 39028 8230 39080 8236
rect 38844 7880 38896 7886
rect 38844 7822 38896 7828
rect 38856 6458 38884 7822
rect 38936 7200 38988 7206
rect 38936 7142 38988 7148
rect 38844 6452 38896 6458
rect 38844 6394 38896 6400
rect 38948 6254 38976 7142
rect 39040 6798 39068 8230
rect 39120 7744 39172 7750
rect 39120 7686 39172 7692
rect 39028 6792 39080 6798
rect 39028 6734 39080 6740
rect 39028 6656 39080 6662
rect 39028 6598 39080 6604
rect 38936 6248 38988 6254
rect 38936 6190 38988 6196
rect 38844 5840 38896 5846
rect 38844 5782 38896 5788
rect 38672 2746 38792 2774
rect 38384 2440 38436 2446
rect 38384 2382 38436 2388
rect 38396 1970 38424 2382
rect 38384 1964 38436 1970
rect 38384 1906 38436 1912
rect 38292 1896 38344 1902
rect 38292 1838 38344 1844
rect 38200 1828 38252 1834
rect 38200 1770 38252 1776
rect 38672 800 38700 2746
rect 38856 2650 38884 5782
rect 38936 5568 38988 5574
rect 38936 5510 38988 5516
rect 38948 5370 38976 5510
rect 38936 5364 38988 5370
rect 38936 5306 38988 5312
rect 38948 4690 38976 5306
rect 38936 4684 38988 4690
rect 38936 4626 38988 4632
rect 39040 4486 39068 6598
rect 39028 4480 39080 4486
rect 39028 4422 39080 4428
rect 39132 3534 39160 7686
rect 39224 4146 39252 8298
rect 39304 6656 39356 6662
rect 39304 6598 39356 6604
rect 39316 5778 39344 6598
rect 39304 5772 39356 5778
rect 39304 5714 39356 5720
rect 39408 5284 39436 8366
rect 39856 8356 39908 8362
rect 39856 8298 39908 8304
rect 39580 6860 39632 6866
rect 39580 6802 39632 6808
rect 39672 6860 39724 6866
rect 39672 6802 39724 6808
rect 39488 6724 39540 6730
rect 39488 6666 39540 6672
rect 39500 6118 39528 6666
rect 39592 6322 39620 6802
rect 39580 6316 39632 6322
rect 39580 6258 39632 6264
rect 39488 6112 39540 6118
rect 39488 6054 39540 6060
rect 39316 5256 39436 5284
rect 39212 4140 39264 4146
rect 39212 4082 39264 4088
rect 39120 3528 39172 3534
rect 39120 3470 39172 3476
rect 38844 2644 38896 2650
rect 38844 2586 38896 2592
rect 39316 800 39344 5256
rect 39592 4554 39620 6258
rect 39684 5846 39712 6802
rect 39672 5840 39724 5846
rect 39672 5782 39724 5788
rect 39580 4548 39632 4554
rect 39632 4508 39804 4536
rect 39580 4490 39632 4496
rect 39488 4140 39540 4146
rect 39488 4082 39540 4088
rect 39396 3460 39448 3466
rect 39396 3402 39448 3408
rect 39408 2446 39436 3402
rect 39500 2514 39528 4082
rect 39776 3058 39804 4508
rect 39764 3052 39816 3058
rect 39764 2994 39816 3000
rect 39868 2961 39896 8298
rect 40052 7546 40080 9454
rect 66574 9276 66882 9285
rect 66574 9274 66580 9276
rect 66636 9274 66660 9276
rect 66716 9274 66740 9276
rect 66796 9274 66820 9276
rect 66876 9274 66882 9276
rect 66636 9222 66638 9274
rect 66818 9222 66820 9274
rect 66574 9220 66580 9222
rect 66636 9220 66660 9222
rect 66716 9220 66740 9222
rect 66796 9220 66820 9222
rect 66876 9220 66882 9222
rect 66574 9211 66882 9220
rect 67234 8732 67542 8741
rect 67234 8730 67240 8732
rect 67296 8730 67320 8732
rect 67376 8730 67400 8732
rect 67456 8730 67480 8732
rect 67536 8730 67542 8732
rect 67296 8678 67298 8730
rect 67478 8678 67480 8730
rect 67234 8676 67240 8678
rect 67296 8676 67320 8678
rect 67376 8676 67400 8678
rect 67456 8676 67480 8678
rect 67536 8676 67542 8678
rect 67234 8667 67542 8676
rect 41420 8356 41472 8362
rect 41420 8298 41472 8304
rect 40222 7984 40278 7993
rect 41432 7954 41460 8298
rect 66574 8188 66882 8197
rect 66574 8186 66580 8188
rect 66636 8186 66660 8188
rect 66716 8186 66740 8188
rect 66796 8186 66820 8188
rect 66876 8186 66882 8188
rect 66636 8134 66638 8186
rect 66818 8134 66820 8186
rect 66574 8132 66580 8134
rect 66636 8132 66660 8134
rect 66716 8132 66740 8134
rect 66796 8132 66820 8134
rect 66876 8132 66882 8134
rect 66574 8123 66882 8132
rect 40222 7919 40278 7928
rect 41420 7948 41472 7954
rect 40132 7744 40184 7750
rect 40132 7686 40184 7692
rect 40040 7540 40092 7546
rect 40040 7482 40092 7488
rect 39948 5568 40000 5574
rect 39948 5510 40000 5516
rect 39960 5234 39988 5510
rect 39948 5228 40000 5234
rect 39948 5170 40000 5176
rect 39946 5128 40002 5137
rect 39946 5063 40002 5072
rect 39960 4554 39988 5063
rect 40144 4729 40172 7686
rect 40236 6798 40264 7919
rect 41420 7890 41472 7896
rect 46480 7880 46532 7886
rect 41602 7848 41658 7857
rect 41236 7812 41288 7818
rect 46480 7822 46532 7828
rect 41602 7783 41604 7792
rect 41236 7754 41288 7760
rect 41656 7783 41658 7792
rect 41604 7754 41656 7760
rect 41248 7478 41276 7754
rect 41788 7744 41840 7750
rect 41788 7686 41840 7692
rect 41236 7472 41288 7478
rect 41236 7414 41288 7420
rect 41604 7336 41656 7342
rect 41604 7278 41656 7284
rect 40592 7200 40644 7206
rect 40592 7142 40644 7148
rect 40224 6792 40276 6798
rect 40224 6734 40276 6740
rect 40236 6390 40264 6734
rect 40408 6724 40460 6730
rect 40408 6666 40460 6672
rect 40224 6384 40276 6390
rect 40224 6326 40276 6332
rect 40130 4720 40186 4729
rect 40130 4655 40186 4664
rect 39948 4548 40000 4554
rect 39948 4490 40000 4496
rect 39960 4457 39988 4490
rect 39946 4448 40002 4457
rect 39946 4383 40002 4392
rect 40420 4146 40448 6666
rect 40498 5128 40554 5137
rect 40498 5063 40554 5072
rect 40512 4622 40540 5063
rect 40500 4616 40552 4622
rect 40500 4558 40552 4564
rect 40408 4140 40460 4146
rect 40408 4082 40460 4088
rect 40500 4140 40552 4146
rect 40500 4082 40552 4088
rect 40316 4072 40368 4078
rect 40316 4014 40368 4020
rect 39948 3936 40000 3942
rect 39948 3878 40000 3884
rect 39960 3641 39988 3878
rect 40328 3738 40356 4014
rect 40316 3732 40368 3738
rect 40316 3674 40368 3680
rect 39946 3632 40002 3641
rect 39946 3567 40002 3576
rect 39854 2952 39910 2961
rect 39854 2887 39910 2896
rect 40328 2854 40356 3674
rect 40420 2922 40448 4082
rect 40512 3641 40540 4082
rect 40498 3632 40554 3641
rect 40498 3567 40554 3576
rect 40604 3534 40632 7142
rect 41420 6656 41472 6662
rect 41420 6598 41472 6604
rect 41512 6656 41564 6662
rect 41512 6598 41564 6604
rect 41432 6322 41460 6598
rect 41420 6316 41472 6322
rect 41420 6258 41472 6264
rect 41144 6112 41196 6118
rect 41144 6054 41196 6060
rect 41156 5778 41184 6054
rect 41144 5772 41196 5778
rect 41144 5714 41196 5720
rect 40776 5568 40828 5574
rect 40776 5510 40828 5516
rect 40788 5234 40816 5510
rect 40776 5228 40828 5234
rect 40776 5170 40828 5176
rect 41328 5228 41380 5234
rect 41328 5170 41380 5176
rect 41144 4616 41196 4622
rect 41144 4558 41196 4564
rect 40776 4548 40828 4554
rect 40776 4490 40828 4496
rect 41052 4548 41104 4554
rect 41052 4490 41104 4496
rect 40788 4321 40816 4490
rect 40774 4312 40830 4321
rect 40774 4247 40830 4256
rect 40788 4060 40816 4247
rect 40696 4032 40816 4060
rect 40592 3528 40644 3534
rect 40592 3470 40644 3476
rect 40696 3398 40724 4032
rect 41064 3534 41092 4490
rect 41052 3528 41104 3534
rect 41052 3470 41104 3476
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 40776 3392 40828 3398
rect 40776 3334 40828 3340
rect 40408 2916 40460 2922
rect 40408 2858 40460 2864
rect 40316 2848 40368 2854
rect 40316 2790 40368 2796
rect 40328 2514 40356 2790
rect 39488 2508 39540 2514
rect 39488 2450 39540 2456
rect 39948 2508 40000 2514
rect 39948 2450 40000 2456
rect 40316 2508 40368 2514
rect 40316 2450 40368 2456
rect 39396 2440 39448 2446
rect 39396 2382 39448 2388
rect 39960 800 39988 2450
rect 40592 2032 40644 2038
rect 40592 1974 40644 1980
rect 40604 800 40632 1974
rect 40788 1766 40816 3334
rect 41156 2990 41184 4558
rect 41236 3936 41288 3942
rect 41236 3878 41288 3884
rect 41248 3534 41276 3878
rect 41340 3777 41368 5170
rect 41326 3768 41382 3777
rect 41524 3738 41552 6598
rect 41326 3703 41382 3712
rect 41512 3732 41564 3738
rect 41512 3674 41564 3680
rect 41236 3528 41288 3534
rect 41236 3470 41288 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41144 2984 41196 2990
rect 41144 2926 41196 2932
rect 41156 2446 41184 2926
rect 41144 2440 41196 2446
rect 41144 2382 41196 2388
rect 41052 2372 41104 2378
rect 41052 2314 41104 2320
rect 40776 1760 40828 1766
rect 40776 1702 40828 1708
rect 41064 1306 41092 2314
rect 41340 2310 41368 3470
rect 41616 2650 41644 7278
rect 41696 5160 41748 5166
rect 41696 5102 41748 5108
rect 41708 4826 41736 5102
rect 41696 4820 41748 4826
rect 41696 4762 41748 4768
rect 41696 4480 41748 4486
rect 41696 4422 41748 4428
rect 41708 3602 41736 4422
rect 41800 3913 41828 7686
rect 42156 7200 42208 7206
rect 42156 7142 42208 7148
rect 41972 6112 42024 6118
rect 41972 6054 42024 6060
rect 41880 4480 41932 4486
rect 41880 4422 41932 4428
rect 41786 3904 41842 3913
rect 41786 3839 41842 3848
rect 41892 3738 41920 4422
rect 41880 3732 41932 3738
rect 41880 3674 41932 3680
rect 41696 3596 41748 3602
rect 41696 3538 41748 3544
rect 41604 2644 41656 2650
rect 41604 2586 41656 2592
rect 41984 2446 42012 6054
rect 42064 5024 42116 5030
rect 42064 4966 42116 4972
rect 42076 4826 42104 4966
rect 42064 4820 42116 4826
rect 42064 4762 42116 4768
rect 42064 4072 42116 4078
rect 42064 4014 42116 4020
rect 42076 3194 42104 4014
rect 42064 3188 42116 3194
rect 42064 3130 42116 3136
rect 42168 2990 42196 7142
rect 43352 6384 43404 6390
rect 43352 6326 43404 6332
rect 42708 6316 42760 6322
rect 42708 6258 42760 6264
rect 42800 6316 42852 6322
rect 42800 6258 42852 6264
rect 43260 6316 43312 6322
rect 43260 6258 43312 6264
rect 42616 6112 42668 6118
rect 42616 6054 42668 6060
rect 42340 4276 42392 4282
rect 42340 4218 42392 4224
rect 42524 4276 42576 4282
rect 42524 4218 42576 4224
rect 42352 3942 42380 4218
rect 42536 4146 42564 4218
rect 42524 4140 42576 4146
rect 42524 4082 42576 4088
rect 42340 3936 42392 3942
rect 42340 3878 42392 3884
rect 42536 3670 42564 4082
rect 42524 3664 42576 3670
rect 42524 3606 42576 3612
rect 42248 3596 42300 3602
rect 42248 3538 42300 3544
rect 42260 3058 42288 3538
rect 42524 3460 42576 3466
rect 42524 3402 42576 3408
rect 42536 3369 42564 3402
rect 42522 3360 42578 3369
rect 42522 3295 42578 3304
rect 42248 3052 42300 3058
rect 42248 2994 42300 3000
rect 42156 2984 42208 2990
rect 42156 2926 42208 2932
rect 42628 2774 42656 6054
rect 42720 5370 42748 6258
rect 42812 5846 42840 6258
rect 42800 5840 42852 5846
rect 42800 5782 42852 5788
rect 42984 5772 43036 5778
rect 42984 5714 43036 5720
rect 42892 5704 42944 5710
rect 42892 5646 42944 5652
rect 42708 5364 42760 5370
rect 42708 5306 42760 5312
rect 42708 5092 42760 5098
rect 42708 5034 42760 5040
rect 42720 4593 42748 5034
rect 42904 4826 42932 5646
rect 42892 4820 42944 4826
rect 42892 4762 42944 4768
rect 42706 4584 42762 4593
rect 42706 4519 42762 4528
rect 42706 4448 42762 4457
rect 42706 4383 42762 4392
rect 42720 4146 42748 4383
rect 42890 4312 42946 4321
rect 42890 4247 42946 4256
rect 42708 4140 42760 4146
rect 42708 4082 42760 4088
rect 42904 4078 42932 4247
rect 42800 4072 42852 4078
rect 42800 4014 42852 4020
rect 42892 4072 42944 4078
rect 42892 4014 42944 4020
rect 42812 3942 42840 4014
rect 42800 3936 42852 3942
rect 42800 3878 42852 3884
rect 42996 3194 43024 5714
rect 43272 5114 43300 6258
rect 43180 5086 43300 5114
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 42984 3188 43036 3194
rect 42984 3130 43036 3136
rect 43088 2990 43116 4014
rect 43076 2984 43128 2990
rect 43076 2926 43128 2932
rect 42536 2746 42656 2774
rect 41972 2440 42024 2446
rect 41972 2382 42024 2388
rect 41880 2372 41932 2378
rect 41880 2314 41932 2320
rect 41328 2304 41380 2310
rect 41328 2246 41380 2252
rect 41064 1278 41276 1306
rect 41248 800 41276 1278
rect 41892 800 41920 2314
rect 42536 800 42564 2746
rect 43180 800 43208 5086
rect 43364 5030 43392 6326
rect 45468 6180 45520 6186
rect 45468 6122 45520 6128
rect 45192 5772 45244 5778
rect 45112 5732 45192 5760
rect 44364 5704 44416 5710
rect 44364 5646 44416 5652
rect 43720 5568 43772 5574
rect 43720 5510 43772 5516
rect 43260 5024 43312 5030
rect 43260 4966 43312 4972
rect 43352 5024 43404 5030
rect 43352 4966 43404 4972
rect 43272 4690 43300 4966
rect 43260 4684 43312 4690
rect 43260 4626 43312 4632
rect 43364 4214 43392 4966
rect 43628 4820 43680 4826
rect 43628 4762 43680 4768
rect 43640 4554 43668 4762
rect 43628 4548 43680 4554
rect 43628 4490 43680 4496
rect 43352 4208 43404 4214
rect 43352 4150 43404 4156
rect 43260 4140 43312 4146
rect 43260 4082 43312 4088
rect 43272 3641 43300 4082
rect 43258 3632 43314 3641
rect 43258 3567 43314 3576
rect 43364 3482 43392 4150
rect 43272 3454 43392 3482
rect 43272 3398 43300 3454
rect 43260 3392 43312 3398
rect 43260 3334 43312 3340
rect 43352 3392 43404 3398
rect 43352 3334 43404 3340
rect 43364 3058 43392 3334
rect 43732 3126 43760 5510
rect 44180 5228 44232 5234
rect 44180 5170 44232 5176
rect 43996 4616 44048 4622
rect 43996 4558 44048 4564
rect 44008 4282 44036 4558
rect 43996 4276 44048 4282
rect 43996 4218 44048 4224
rect 43902 4176 43958 4185
rect 43902 4111 43958 4120
rect 43812 3936 43864 3942
rect 43812 3878 43864 3884
rect 43824 3670 43852 3878
rect 43812 3664 43864 3670
rect 43812 3606 43864 3612
rect 43916 3534 43944 4111
rect 44192 4078 44220 5170
rect 44180 4072 44232 4078
rect 44180 4014 44232 4020
rect 43904 3528 43956 3534
rect 43904 3470 43956 3476
rect 44178 3360 44234 3369
rect 44178 3295 44234 3304
rect 44192 3126 44220 3295
rect 44376 3194 44404 5646
rect 44824 5092 44876 5098
rect 44824 5034 44876 5040
rect 44456 4480 44508 4486
rect 44456 4422 44508 4428
rect 44364 3188 44416 3194
rect 44364 3130 44416 3136
rect 43720 3120 43772 3126
rect 43720 3062 43772 3068
rect 44180 3120 44232 3126
rect 44180 3062 44232 3068
rect 43352 3052 43404 3058
rect 43352 2994 43404 3000
rect 44180 2984 44232 2990
rect 44180 2926 44232 2932
rect 44192 1442 44220 2926
rect 44100 1414 44220 1442
rect 43824 870 43944 898
rect 43824 800 43852 870
rect 37476 734 37780 762
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 43916 762 43944 870
rect 44100 762 44128 1414
rect 44468 800 44496 4422
rect 44732 4072 44784 4078
rect 44730 4040 44732 4049
rect 44784 4040 44786 4049
rect 44730 3975 44786 3984
rect 44836 3942 44864 5034
rect 44824 3936 44876 3942
rect 44824 3878 44876 3884
rect 44916 3936 44968 3942
rect 44916 3878 44968 3884
rect 44928 3738 44956 3878
rect 44916 3732 44968 3738
rect 44916 3674 44968 3680
rect 45112 800 45140 5732
rect 45192 5714 45244 5720
rect 45480 4690 45508 6122
rect 45836 5704 45888 5710
rect 45836 5646 45888 5652
rect 45652 5636 45704 5642
rect 45652 5578 45704 5584
rect 45560 5160 45612 5166
rect 45560 5102 45612 5108
rect 45468 4684 45520 4690
rect 45468 4626 45520 4632
rect 45284 4616 45336 4622
rect 45284 4558 45336 4564
rect 45192 3460 45244 3466
rect 45192 3402 45244 3408
rect 45204 3058 45232 3402
rect 45296 3194 45324 4558
rect 45572 3738 45600 5102
rect 45664 4078 45692 5578
rect 45744 5024 45796 5030
rect 45744 4966 45796 4972
rect 45652 4072 45704 4078
rect 45652 4014 45704 4020
rect 45756 3890 45784 4966
rect 45848 4826 45876 5646
rect 45836 4820 45888 4826
rect 45836 4762 45888 4768
rect 46492 4146 46520 7822
rect 67234 7644 67542 7653
rect 67234 7642 67240 7644
rect 67296 7642 67320 7644
rect 67376 7642 67400 7644
rect 67456 7642 67480 7644
rect 67536 7642 67542 7644
rect 67296 7590 67298 7642
rect 67478 7590 67480 7642
rect 67234 7588 67240 7590
rect 67296 7588 67320 7590
rect 67376 7588 67400 7590
rect 67456 7588 67480 7590
rect 67536 7588 67542 7590
rect 67234 7579 67542 7588
rect 66574 7100 66882 7109
rect 66574 7098 66580 7100
rect 66636 7098 66660 7100
rect 66716 7098 66740 7100
rect 66796 7098 66820 7100
rect 66876 7098 66882 7100
rect 66636 7046 66638 7098
rect 66818 7046 66820 7098
rect 66574 7044 66580 7046
rect 66636 7044 66660 7046
rect 66716 7044 66740 7046
rect 66796 7044 66820 7046
rect 66876 7044 66882 7046
rect 66574 7035 66882 7044
rect 46848 6656 46900 6662
rect 46848 6598 46900 6604
rect 46756 5228 46808 5234
rect 46756 5170 46808 5176
rect 46480 4140 46532 4146
rect 46480 4082 46532 4088
rect 46388 3936 46440 3942
rect 45756 3862 45876 3890
rect 46388 3878 46440 3884
rect 45560 3732 45612 3738
rect 45560 3674 45612 3680
rect 45284 3188 45336 3194
rect 45284 3130 45336 3136
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 45296 2854 45324 3130
rect 45744 2984 45796 2990
rect 45744 2926 45796 2932
rect 45284 2848 45336 2854
rect 45284 2790 45336 2796
rect 45756 800 45784 2926
rect 45848 2446 45876 3862
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 46400 800 46428 3878
rect 46768 3738 46796 5170
rect 46756 3732 46808 3738
rect 46756 3674 46808 3680
rect 46860 3602 46888 6598
rect 67234 6556 67542 6565
rect 67234 6554 67240 6556
rect 67296 6554 67320 6556
rect 67376 6554 67400 6556
rect 67456 6554 67480 6556
rect 67536 6554 67542 6556
rect 67296 6502 67298 6554
rect 67478 6502 67480 6554
rect 67234 6500 67240 6502
rect 67296 6500 67320 6502
rect 67376 6500 67400 6502
rect 67456 6500 67480 6502
rect 67536 6500 67542 6502
rect 67234 6491 67542 6500
rect 48872 6112 48924 6118
rect 48872 6054 48924 6060
rect 47032 5568 47084 5574
rect 47032 5510 47084 5516
rect 47044 5234 47072 5510
rect 47032 5228 47084 5234
rect 47032 5170 47084 5176
rect 46940 5160 46992 5166
rect 46940 5102 46992 5108
rect 46848 3596 46900 3602
rect 46848 3538 46900 3544
rect 46952 3194 46980 5102
rect 47952 5092 48004 5098
rect 47952 5034 48004 5040
rect 47216 5024 47268 5030
rect 47216 4966 47268 4972
rect 47228 4690 47256 4966
rect 47216 4684 47268 4690
rect 47216 4626 47268 4632
rect 47860 4480 47912 4486
rect 47860 4422 47912 4428
rect 47584 4004 47636 4010
rect 47584 3946 47636 3952
rect 47124 3528 47176 3534
rect 47124 3470 47176 3476
rect 46940 3188 46992 3194
rect 46940 3130 46992 3136
rect 46756 3052 46808 3058
rect 46756 2994 46808 3000
rect 46768 2514 46796 2994
rect 47136 2650 47164 3470
rect 47124 2644 47176 2650
rect 47124 2586 47176 2592
rect 46756 2508 46808 2514
rect 46756 2450 46808 2456
rect 47596 2310 47624 3946
rect 47872 3602 47900 4422
rect 47860 3596 47912 3602
rect 47860 3538 47912 3544
rect 47964 3534 47992 5034
rect 48320 4684 48372 4690
rect 48320 4626 48372 4632
rect 48332 4282 48360 4626
rect 48780 4616 48832 4622
rect 48780 4558 48832 4564
rect 48504 4548 48556 4554
rect 48504 4490 48556 4496
rect 48412 4480 48464 4486
rect 48412 4422 48464 4428
rect 48320 4276 48372 4282
rect 48320 4218 48372 4224
rect 48044 4140 48096 4146
rect 48044 4082 48096 4088
rect 48056 3738 48084 4082
rect 48318 3904 48374 3913
rect 48318 3839 48374 3848
rect 48044 3732 48096 3738
rect 48044 3674 48096 3680
rect 47952 3528 48004 3534
rect 47952 3470 48004 3476
rect 48136 3392 48188 3398
rect 48136 3334 48188 3340
rect 47676 2984 47728 2990
rect 47676 2926 47728 2932
rect 47584 2304 47636 2310
rect 47584 2246 47636 2252
rect 47688 800 47716 2926
rect 48148 2582 48176 3334
rect 48332 3194 48360 3839
rect 48320 3188 48372 3194
rect 48320 3130 48372 3136
rect 48136 2576 48188 2582
rect 48136 2518 48188 2524
rect 48424 2446 48452 4422
rect 48516 4146 48544 4490
rect 48792 4282 48820 4558
rect 48780 4276 48832 4282
rect 48780 4218 48832 4224
rect 48504 4140 48556 4146
rect 48504 4082 48556 4088
rect 48884 3602 48912 6054
rect 66574 6012 66882 6021
rect 66574 6010 66580 6012
rect 66636 6010 66660 6012
rect 66716 6010 66740 6012
rect 66796 6010 66820 6012
rect 66876 6010 66882 6012
rect 66636 5958 66638 6010
rect 66818 5958 66820 6010
rect 66574 5956 66580 5958
rect 66636 5956 66660 5958
rect 66716 5956 66740 5958
rect 66796 5956 66820 5958
rect 66876 5956 66882 5958
rect 66574 5947 66882 5956
rect 67234 5468 67542 5477
rect 67234 5466 67240 5468
rect 67296 5466 67320 5468
rect 67376 5466 67400 5468
rect 67456 5466 67480 5468
rect 67536 5466 67542 5468
rect 67296 5414 67298 5466
rect 67478 5414 67480 5466
rect 67234 5412 67240 5414
rect 67296 5412 67320 5414
rect 67376 5412 67400 5414
rect 67456 5412 67480 5414
rect 67536 5412 67542 5414
rect 67234 5403 67542 5412
rect 76932 5160 76984 5166
rect 76932 5102 76984 5108
rect 49608 5024 49660 5030
rect 49608 4966 49660 4972
rect 76656 5024 76708 5030
rect 76656 4966 76708 4972
rect 48872 3596 48924 3602
rect 48872 3538 48924 3544
rect 49620 2990 49648 4966
rect 66574 4924 66882 4933
rect 66574 4922 66580 4924
rect 66636 4922 66660 4924
rect 66716 4922 66740 4924
rect 66796 4922 66820 4924
rect 66876 4922 66882 4924
rect 66636 4870 66638 4922
rect 66818 4870 66820 4922
rect 66574 4868 66580 4870
rect 66636 4868 66660 4870
rect 66716 4868 66740 4870
rect 66796 4868 66820 4870
rect 66876 4868 66882 4870
rect 66574 4859 66882 4868
rect 49700 4480 49752 4486
rect 49700 4422 49752 4428
rect 49608 2984 49660 2990
rect 49608 2926 49660 2932
rect 49608 2576 49660 2582
rect 49608 2518 49660 2524
rect 47952 2440 48004 2446
rect 47952 2382 48004 2388
rect 48412 2440 48464 2446
rect 48412 2382 48464 2388
rect 47964 2106 47992 2382
rect 47952 2100 48004 2106
rect 47952 2042 48004 2048
rect 49620 800 49648 2518
rect 49712 2446 49740 4422
rect 67234 4380 67542 4389
rect 67234 4378 67240 4380
rect 67296 4378 67320 4380
rect 67376 4378 67400 4380
rect 67456 4378 67480 4380
rect 67536 4378 67542 4380
rect 67296 4326 67298 4378
rect 67478 4326 67480 4378
rect 67234 4324 67240 4326
rect 67296 4324 67320 4326
rect 67376 4324 67400 4326
rect 67456 4324 67480 4326
rect 67536 4324 67542 4326
rect 67234 4315 67542 4324
rect 74632 4140 74684 4146
rect 74632 4082 74684 4088
rect 53196 4072 53248 4078
rect 53196 4014 53248 4020
rect 53840 4072 53892 4078
rect 53840 4014 53892 4020
rect 65432 4072 65484 4078
rect 65432 4014 65484 4020
rect 68652 4072 68704 4078
rect 68652 4014 68704 4020
rect 69296 4072 69348 4078
rect 69296 4014 69348 4020
rect 71688 4072 71740 4078
rect 71688 4014 71740 4020
rect 74264 4072 74316 4078
rect 74264 4014 74316 4020
rect 51356 3936 51408 3942
rect 51356 3878 51408 3884
rect 52828 3936 52880 3942
rect 52828 3878 52880 3884
rect 50804 3528 50856 3534
rect 50804 3470 50856 3476
rect 50528 3460 50580 3466
rect 50528 3402 50580 3408
rect 49976 3392 50028 3398
rect 49976 3334 50028 3340
rect 49792 3052 49844 3058
rect 49792 2994 49844 3000
rect 49804 2514 49832 2994
rect 49988 2650 50016 3334
rect 49976 2644 50028 2650
rect 49976 2586 50028 2592
rect 50540 2514 50568 3402
rect 50816 3194 50844 3470
rect 50804 3188 50856 3194
rect 50804 3130 50856 3136
rect 51368 3058 51396 3878
rect 51356 3052 51408 3058
rect 51356 2994 51408 3000
rect 52092 3052 52144 3058
rect 52092 2994 52144 3000
rect 51540 2916 51592 2922
rect 51540 2858 51592 2864
rect 49792 2508 49844 2514
rect 49792 2450 49844 2456
rect 50528 2508 50580 2514
rect 50528 2450 50580 2456
rect 49700 2440 49752 2446
rect 49700 2382 49752 2388
rect 51552 800 51580 2858
rect 52104 2514 52132 2994
rect 52092 2508 52144 2514
rect 52092 2450 52144 2456
rect 52840 2446 52868 3878
rect 53208 3738 53236 4014
rect 53196 3732 53248 3738
rect 53196 3674 53248 3680
rect 53012 3528 53064 3534
rect 53012 3470 53064 3476
rect 53024 3194 53052 3470
rect 53852 3194 53880 4014
rect 54024 3936 54076 3942
rect 54024 3878 54076 3884
rect 54036 3602 54064 3878
rect 54024 3596 54076 3602
rect 54024 3538 54076 3544
rect 59452 3528 59504 3534
rect 59452 3470 59504 3476
rect 63408 3528 63460 3534
rect 63408 3470 63460 3476
rect 64512 3528 64564 3534
rect 64512 3470 64564 3476
rect 57336 3460 57388 3466
rect 57336 3402 57388 3408
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 53012 3188 53064 3194
rect 53012 3130 53064 3136
rect 53840 3188 53892 3194
rect 53840 3130 53892 3136
rect 56060 3058 56088 3334
rect 57348 3194 57376 3402
rect 57428 3392 57480 3398
rect 57428 3334 57480 3340
rect 58624 3392 58676 3398
rect 58624 3334 58676 3340
rect 57336 3188 57388 3194
rect 57336 3130 57388 3136
rect 57440 3058 57468 3334
rect 54024 3052 54076 3058
rect 54024 2994 54076 3000
rect 56048 3052 56100 3058
rect 56048 2994 56100 3000
rect 57428 3052 57480 3058
rect 57428 2994 57480 3000
rect 53472 2984 53524 2990
rect 53472 2926 53524 2932
rect 52828 2440 52880 2446
rect 52828 2382 52880 2388
rect 53484 800 53512 2926
rect 54036 2514 54064 2994
rect 55312 2848 55364 2854
rect 55312 2790 55364 2796
rect 54024 2508 54076 2514
rect 54024 2450 54076 2456
rect 55324 2446 55352 2790
rect 58636 2446 58664 3334
rect 59464 3194 59492 3470
rect 60924 3460 60976 3466
rect 60924 3402 60976 3408
rect 60936 3194 60964 3402
rect 61108 3392 61160 3398
rect 61108 3334 61160 3340
rect 62764 3392 62816 3398
rect 62764 3334 62816 3340
rect 59452 3188 59504 3194
rect 59452 3130 59504 3136
rect 60924 3188 60976 3194
rect 60924 3130 60976 3136
rect 61120 3058 61148 3334
rect 61108 3052 61160 3058
rect 61108 2994 61160 3000
rect 61752 3052 61804 3058
rect 61752 2994 61804 3000
rect 61200 2984 61252 2990
rect 61200 2926 61252 2932
rect 59268 2848 59320 2854
rect 59268 2790 59320 2796
rect 55312 2440 55364 2446
rect 55312 2382 55364 2388
rect 55404 2440 55456 2446
rect 55404 2382 55456 2388
rect 58624 2440 58676 2446
rect 58624 2382 58676 2388
rect 55416 800 55444 2382
rect 57336 2372 57388 2378
rect 57336 2314 57388 2320
rect 57348 800 57376 2314
rect 59280 800 59308 2790
rect 61212 800 61240 2926
rect 61764 2514 61792 2994
rect 61752 2508 61804 2514
rect 61752 2450 61804 2456
rect 62776 2446 62804 3334
rect 63420 3194 63448 3470
rect 64524 3194 64552 3470
rect 64880 3392 64932 3398
rect 64880 3334 64932 3340
rect 63408 3188 63460 3194
rect 63408 3130 63460 3136
rect 64512 3188 64564 3194
rect 64512 3130 64564 3136
rect 64892 3058 64920 3334
rect 65444 3194 65472 4014
rect 66260 3936 66312 3942
rect 66260 3878 66312 3884
rect 68284 3936 68336 3942
rect 68284 3878 68336 3884
rect 65432 3188 65484 3194
rect 65432 3130 65484 3136
rect 64880 3052 64932 3058
rect 64880 2994 64932 3000
rect 65524 3052 65576 3058
rect 65524 2994 65576 3000
rect 65064 2984 65116 2990
rect 65064 2926 65116 2932
rect 62764 2440 62816 2446
rect 62764 2382 62816 2388
rect 63132 2440 63184 2446
rect 63132 2382 63184 2388
rect 63144 800 63172 2382
rect 65076 800 65104 2926
rect 65536 2514 65564 2994
rect 65524 2508 65576 2514
rect 65524 2450 65576 2456
rect 66272 2446 66300 3878
rect 66574 3836 66882 3845
rect 66574 3834 66580 3836
rect 66636 3834 66660 3836
rect 66716 3834 66740 3836
rect 66796 3834 66820 3836
rect 66876 3834 66882 3836
rect 66636 3782 66638 3834
rect 66818 3782 66820 3834
rect 66574 3780 66580 3782
rect 66636 3780 66660 3782
rect 66716 3780 66740 3782
rect 66796 3780 66820 3782
rect 66876 3780 66882 3782
rect 66574 3771 66882 3780
rect 67234 3292 67542 3301
rect 67234 3290 67240 3292
rect 67296 3290 67320 3292
rect 67376 3290 67400 3292
rect 67456 3290 67480 3292
rect 67536 3290 67542 3292
rect 67296 3238 67298 3290
rect 67478 3238 67480 3290
rect 67234 3236 67240 3238
rect 67296 3236 67320 3238
rect 67376 3236 67400 3238
rect 67456 3236 67480 3238
rect 67536 3236 67542 3238
rect 67234 3227 67542 3236
rect 67640 3052 67692 3058
rect 67640 2994 67692 3000
rect 66996 2916 67048 2922
rect 66996 2858 67048 2864
rect 66574 2748 66882 2757
rect 66574 2746 66580 2748
rect 66636 2746 66660 2748
rect 66716 2746 66740 2748
rect 66796 2746 66820 2748
rect 66876 2746 66882 2748
rect 66636 2694 66638 2746
rect 66818 2694 66820 2746
rect 66574 2692 66580 2694
rect 66636 2692 66660 2694
rect 66716 2692 66740 2694
rect 66796 2692 66820 2694
rect 66876 2692 66882 2694
rect 66574 2683 66882 2692
rect 66260 2440 66312 2446
rect 66260 2382 66312 2388
rect 67008 800 67036 2858
rect 67652 2514 67680 2994
rect 67640 2508 67692 2514
rect 67640 2450 67692 2456
rect 68296 2446 68324 3878
rect 68664 3738 68692 4014
rect 68652 3732 68704 3738
rect 68652 3674 68704 3680
rect 68468 3528 68520 3534
rect 68468 3470 68520 3476
rect 68480 3194 68508 3470
rect 69308 3194 69336 4014
rect 69480 3936 69532 3942
rect 69480 3878 69532 3884
rect 69492 3602 69520 3878
rect 71700 3738 71728 4014
rect 73712 3936 73764 3942
rect 73712 3878 73764 3884
rect 71688 3732 71740 3738
rect 71688 3674 71740 3680
rect 73724 3602 73752 3878
rect 69480 3596 69532 3602
rect 69480 3538 69532 3544
rect 73712 3596 73764 3602
rect 73712 3538 73764 3544
rect 72976 3528 73028 3534
rect 72976 3470 73028 3476
rect 71504 3392 71556 3398
rect 71504 3334 71556 3340
rect 68468 3188 68520 3194
rect 68468 3130 68520 3136
rect 69296 3188 69348 3194
rect 69296 3130 69348 3136
rect 70308 3120 70360 3126
rect 70308 3062 70360 3068
rect 69480 3052 69532 3058
rect 69480 2994 69532 3000
rect 68928 2984 68980 2990
rect 68928 2926 68980 2932
rect 68284 2440 68336 2446
rect 68284 2382 68336 2388
rect 67234 2204 67542 2213
rect 67234 2202 67240 2204
rect 67296 2202 67320 2204
rect 67376 2202 67400 2204
rect 67456 2202 67480 2204
rect 67536 2202 67542 2204
rect 67296 2150 67298 2202
rect 67478 2150 67480 2202
rect 67234 2148 67240 2150
rect 67296 2148 67320 2150
rect 67376 2148 67400 2150
rect 67456 2148 67480 2150
rect 67536 2148 67542 2150
rect 67234 2139 67542 2148
rect 68940 800 68968 2926
rect 69492 2514 69520 2994
rect 70320 2514 70348 3062
rect 71516 3058 71544 3334
rect 71504 3052 71556 3058
rect 71504 2994 71556 3000
rect 72608 3052 72660 3058
rect 72608 2994 72660 3000
rect 70860 2984 70912 2990
rect 70860 2926 70912 2932
rect 70492 2848 70544 2854
rect 70492 2790 70544 2796
rect 69480 2508 69532 2514
rect 69480 2450 69532 2456
rect 70308 2508 70360 2514
rect 70308 2450 70360 2456
rect 70504 2446 70532 2790
rect 70492 2440 70544 2446
rect 70492 2382 70544 2388
rect 70872 800 70900 2926
rect 72620 2514 72648 2994
rect 72988 2650 73016 3470
rect 73252 3392 73304 3398
rect 73252 3334 73304 3340
rect 72976 2644 73028 2650
rect 72976 2586 73028 2592
rect 72608 2508 72660 2514
rect 72608 2450 72660 2456
rect 72792 2508 72844 2514
rect 72792 2450 72844 2456
rect 72804 800 72832 2450
rect 73264 2446 73292 3334
rect 74276 3058 74304 4014
rect 74448 3528 74500 3534
rect 74448 3470 74500 3476
rect 74460 3194 74488 3470
rect 74540 3392 74592 3398
rect 74540 3334 74592 3340
rect 74448 3188 74500 3194
rect 74448 3130 74500 3136
rect 74552 3058 74580 3334
rect 74264 3052 74316 3058
rect 74264 2994 74316 3000
rect 74540 3052 74592 3058
rect 74540 2994 74592 3000
rect 73252 2440 73304 2446
rect 73252 2382 73304 2388
rect 74276 1873 74304 2994
rect 74644 2650 74672 4082
rect 76564 4072 76616 4078
rect 76564 4014 76616 4020
rect 75460 3460 75512 3466
rect 75460 3402 75512 3408
rect 74724 2984 74776 2990
rect 74724 2926 74776 2932
rect 74632 2644 74684 2650
rect 74632 2586 74684 2592
rect 74262 1864 74318 1873
rect 74262 1799 74318 1808
rect 74736 800 74764 2926
rect 75472 2514 75500 3402
rect 76196 2848 76248 2854
rect 76196 2790 76248 2796
rect 75460 2508 75512 2514
rect 75460 2450 75512 2456
rect 76208 2446 76236 2790
rect 76196 2440 76248 2446
rect 76196 2382 76248 2388
rect 76576 2122 76604 4014
rect 76668 3534 76696 4966
rect 76944 4826 76972 5102
rect 76932 4820 76984 4826
rect 76932 4762 76984 4768
rect 77576 4616 77628 4622
rect 77576 4558 77628 4564
rect 77024 4072 77076 4078
rect 77024 4014 77076 4020
rect 77036 3602 77064 4014
rect 77588 3738 77616 4558
rect 77576 3732 77628 3738
rect 77576 3674 77628 3680
rect 77024 3596 77076 3602
rect 77024 3538 77076 3544
rect 76656 3528 76708 3534
rect 76656 3470 76708 3476
rect 76656 3052 76708 3058
rect 76656 2994 76708 3000
rect 76668 2650 76696 2994
rect 76656 2644 76708 2650
rect 76656 2586 76708 2592
rect 76576 2094 76696 2122
rect 76668 800 76696 2094
rect 43916 734 44128 762
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 77298 0 77354 800
<< via2 >>
rect 5140 37562 5196 37564
rect 5220 37562 5276 37564
rect 5300 37562 5356 37564
rect 5380 37562 5436 37564
rect 5140 37510 5186 37562
rect 5186 37510 5196 37562
rect 5220 37510 5250 37562
rect 5250 37510 5262 37562
rect 5262 37510 5276 37562
rect 5300 37510 5314 37562
rect 5314 37510 5326 37562
rect 5326 37510 5356 37562
rect 5380 37510 5390 37562
rect 5390 37510 5436 37562
rect 5140 37508 5196 37510
rect 5220 37508 5276 37510
rect 5300 37508 5356 37510
rect 5380 37508 5436 37510
rect 5800 37018 5856 37020
rect 5880 37018 5936 37020
rect 5960 37018 6016 37020
rect 6040 37018 6096 37020
rect 5800 36966 5846 37018
rect 5846 36966 5856 37018
rect 5880 36966 5910 37018
rect 5910 36966 5922 37018
rect 5922 36966 5936 37018
rect 5960 36966 5974 37018
rect 5974 36966 5986 37018
rect 5986 36966 6016 37018
rect 6040 36966 6050 37018
rect 6050 36966 6096 37018
rect 5800 36964 5856 36966
rect 5880 36964 5936 36966
rect 5960 36964 6016 36966
rect 6040 36964 6096 36966
rect 5140 36474 5196 36476
rect 5220 36474 5276 36476
rect 5300 36474 5356 36476
rect 5380 36474 5436 36476
rect 5140 36422 5186 36474
rect 5186 36422 5196 36474
rect 5220 36422 5250 36474
rect 5250 36422 5262 36474
rect 5262 36422 5276 36474
rect 5300 36422 5314 36474
rect 5314 36422 5326 36474
rect 5326 36422 5356 36474
rect 5380 36422 5390 36474
rect 5390 36422 5436 36474
rect 5140 36420 5196 36422
rect 5220 36420 5276 36422
rect 5300 36420 5356 36422
rect 5380 36420 5436 36422
rect 5800 35930 5856 35932
rect 5880 35930 5936 35932
rect 5960 35930 6016 35932
rect 6040 35930 6096 35932
rect 5800 35878 5846 35930
rect 5846 35878 5856 35930
rect 5880 35878 5910 35930
rect 5910 35878 5922 35930
rect 5922 35878 5936 35930
rect 5960 35878 5974 35930
rect 5974 35878 5986 35930
rect 5986 35878 6016 35930
rect 6040 35878 6050 35930
rect 6050 35878 6096 35930
rect 5800 35876 5856 35878
rect 5880 35876 5936 35878
rect 5960 35876 6016 35878
rect 6040 35876 6096 35878
rect 5140 35386 5196 35388
rect 5220 35386 5276 35388
rect 5300 35386 5356 35388
rect 5380 35386 5436 35388
rect 5140 35334 5186 35386
rect 5186 35334 5196 35386
rect 5220 35334 5250 35386
rect 5250 35334 5262 35386
rect 5262 35334 5276 35386
rect 5300 35334 5314 35386
rect 5314 35334 5326 35386
rect 5326 35334 5356 35386
rect 5380 35334 5390 35386
rect 5390 35334 5436 35386
rect 5140 35332 5196 35334
rect 5220 35332 5276 35334
rect 5300 35332 5356 35334
rect 5380 35332 5436 35334
rect 5800 34842 5856 34844
rect 5880 34842 5936 34844
rect 5960 34842 6016 34844
rect 6040 34842 6096 34844
rect 5800 34790 5846 34842
rect 5846 34790 5856 34842
rect 5880 34790 5910 34842
rect 5910 34790 5922 34842
rect 5922 34790 5936 34842
rect 5960 34790 5974 34842
rect 5974 34790 5986 34842
rect 5986 34790 6016 34842
rect 6040 34790 6050 34842
rect 6050 34790 6096 34842
rect 5800 34788 5856 34790
rect 5880 34788 5936 34790
rect 5960 34788 6016 34790
rect 6040 34788 6096 34790
rect 5140 34298 5196 34300
rect 5220 34298 5276 34300
rect 5300 34298 5356 34300
rect 5380 34298 5436 34300
rect 5140 34246 5186 34298
rect 5186 34246 5196 34298
rect 5220 34246 5250 34298
rect 5250 34246 5262 34298
rect 5262 34246 5276 34298
rect 5300 34246 5314 34298
rect 5314 34246 5326 34298
rect 5326 34246 5356 34298
rect 5380 34246 5390 34298
rect 5390 34246 5436 34298
rect 5140 34244 5196 34246
rect 5220 34244 5276 34246
rect 5300 34244 5356 34246
rect 5380 34244 5436 34246
rect 5800 33754 5856 33756
rect 5880 33754 5936 33756
rect 5960 33754 6016 33756
rect 6040 33754 6096 33756
rect 5800 33702 5846 33754
rect 5846 33702 5856 33754
rect 5880 33702 5910 33754
rect 5910 33702 5922 33754
rect 5922 33702 5936 33754
rect 5960 33702 5974 33754
rect 5974 33702 5986 33754
rect 5986 33702 6016 33754
rect 6040 33702 6050 33754
rect 6050 33702 6096 33754
rect 5800 33700 5856 33702
rect 5880 33700 5936 33702
rect 5960 33700 6016 33702
rect 6040 33700 6096 33702
rect 5140 33210 5196 33212
rect 5220 33210 5276 33212
rect 5300 33210 5356 33212
rect 5380 33210 5436 33212
rect 5140 33158 5186 33210
rect 5186 33158 5196 33210
rect 5220 33158 5250 33210
rect 5250 33158 5262 33210
rect 5262 33158 5276 33210
rect 5300 33158 5314 33210
rect 5314 33158 5326 33210
rect 5326 33158 5356 33210
rect 5380 33158 5390 33210
rect 5390 33158 5436 33210
rect 5140 33156 5196 33158
rect 5220 33156 5276 33158
rect 5300 33156 5356 33158
rect 5380 33156 5436 33158
rect 5800 32666 5856 32668
rect 5880 32666 5936 32668
rect 5960 32666 6016 32668
rect 6040 32666 6096 32668
rect 5800 32614 5846 32666
rect 5846 32614 5856 32666
rect 5880 32614 5910 32666
rect 5910 32614 5922 32666
rect 5922 32614 5936 32666
rect 5960 32614 5974 32666
rect 5974 32614 5986 32666
rect 5986 32614 6016 32666
rect 6040 32614 6050 32666
rect 6050 32614 6096 32666
rect 5800 32612 5856 32614
rect 5880 32612 5936 32614
rect 5960 32612 6016 32614
rect 6040 32612 6096 32614
rect 7102 32408 7158 32464
rect 5140 32122 5196 32124
rect 5220 32122 5276 32124
rect 5300 32122 5356 32124
rect 5380 32122 5436 32124
rect 5140 32070 5186 32122
rect 5186 32070 5196 32122
rect 5220 32070 5250 32122
rect 5250 32070 5262 32122
rect 5262 32070 5276 32122
rect 5300 32070 5314 32122
rect 5314 32070 5326 32122
rect 5326 32070 5356 32122
rect 5380 32070 5390 32122
rect 5390 32070 5436 32122
rect 5140 32068 5196 32070
rect 5220 32068 5276 32070
rect 5300 32068 5356 32070
rect 5380 32068 5436 32070
rect 5800 31578 5856 31580
rect 5880 31578 5936 31580
rect 5960 31578 6016 31580
rect 6040 31578 6096 31580
rect 5800 31526 5846 31578
rect 5846 31526 5856 31578
rect 5880 31526 5910 31578
rect 5910 31526 5922 31578
rect 5922 31526 5936 31578
rect 5960 31526 5974 31578
rect 5974 31526 5986 31578
rect 5986 31526 6016 31578
rect 6040 31526 6050 31578
rect 6050 31526 6096 31578
rect 5800 31524 5856 31526
rect 5880 31524 5936 31526
rect 5960 31524 6016 31526
rect 6040 31524 6096 31526
rect 5140 31034 5196 31036
rect 5220 31034 5276 31036
rect 5300 31034 5356 31036
rect 5380 31034 5436 31036
rect 5140 30982 5186 31034
rect 5186 30982 5196 31034
rect 5220 30982 5250 31034
rect 5250 30982 5262 31034
rect 5262 30982 5276 31034
rect 5300 30982 5314 31034
rect 5314 30982 5326 31034
rect 5326 30982 5356 31034
rect 5380 30982 5390 31034
rect 5390 30982 5436 31034
rect 5140 30980 5196 30982
rect 5220 30980 5276 30982
rect 5300 30980 5356 30982
rect 5380 30980 5436 30982
rect 5800 30490 5856 30492
rect 5880 30490 5936 30492
rect 5960 30490 6016 30492
rect 6040 30490 6096 30492
rect 5800 30438 5846 30490
rect 5846 30438 5856 30490
rect 5880 30438 5910 30490
rect 5910 30438 5922 30490
rect 5922 30438 5936 30490
rect 5960 30438 5974 30490
rect 5974 30438 5986 30490
rect 5986 30438 6016 30490
rect 6040 30438 6050 30490
rect 6050 30438 6096 30490
rect 5800 30436 5856 30438
rect 5880 30436 5936 30438
rect 5960 30436 6016 30438
rect 6040 30436 6096 30438
rect 5140 29946 5196 29948
rect 5220 29946 5276 29948
rect 5300 29946 5356 29948
rect 5380 29946 5436 29948
rect 5140 29894 5186 29946
rect 5186 29894 5196 29946
rect 5220 29894 5250 29946
rect 5250 29894 5262 29946
rect 5262 29894 5276 29946
rect 5300 29894 5314 29946
rect 5314 29894 5326 29946
rect 5326 29894 5356 29946
rect 5380 29894 5390 29946
rect 5390 29894 5436 29946
rect 5140 29892 5196 29894
rect 5220 29892 5276 29894
rect 5300 29892 5356 29894
rect 5380 29892 5436 29894
rect 10966 29552 11022 29608
rect 5800 29402 5856 29404
rect 5880 29402 5936 29404
rect 5960 29402 6016 29404
rect 6040 29402 6096 29404
rect 5800 29350 5846 29402
rect 5846 29350 5856 29402
rect 5880 29350 5910 29402
rect 5910 29350 5922 29402
rect 5922 29350 5936 29402
rect 5960 29350 5974 29402
rect 5974 29350 5986 29402
rect 5986 29350 6016 29402
rect 6040 29350 6050 29402
rect 6050 29350 6096 29402
rect 5800 29348 5856 29350
rect 5880 29348 5936 29350
rect 5960 29348 6016 29350
rect 6040 29348 6096 29350
rect 5140 28858 5196 28860
rect 5220 28858 5276 28860
rect 5300 28858 5356 28860
rect 5380 28858 5436 28860
rect 5140 28806 5186 28858
rect 5186 28806 5196 28858
rect 5220 28806 5250 28858
rect 5250 28806 5262 28858
rect 5262 28806 5276 28858
rect 5300 28806 5314 28858
rect 5314 28806 5326 28858
rect 5326 28806 5356 28858
rect 5380 28806 5390 28858
rect 5390 28806 5436 28858
rect 5140 28804 5196 28806
rect 5220 28804 5276 28806
rect 5300 28804 5356 28806
rect 5380 28804 5436 28806
rect 5800 28314 5856 28316
rect 5880 28314 5936 28316
rect 5960 28314 6016 28316
rect 6040 28314 6096 28316
rect 5800 28262 5846 28314
rect 5846 28262 5856 28314
rect 5880 28262 5910 28314
rect 5910 28262 5922 28314
rect 5922 28262 5936 28314
rect 5960 28262 5974 28314
rect 5974 28262 5986 28314
rect 5986 28262 6016 28314
rect 6040 28262 6050 28314
rect 6050 28262 6096 28314
rect 5800 28260 5856 28262
rect 5880 28260 5936 28262
rect 5960 28260 6016 28262
rect 6040 28260 6096 28262
rect 5140 27770 5196 27772
rect 5220 27770 5276 27772
rect 5300 27770 5356 27772
rect 5380 27770 5436 27772
rect 5140 27718 5186 27770
rect 5186 27718 5196 27770
rect 5220 27718 5250 27770
rect 5250 27718 5262 27770
rect 5262 27718 5276 27770
rect 5300 27718 5314 27770
rect 5314 27718 5326 27770
rect 5326 27718 5356 27770
rect 5380 27718 5390 27770
rect 5390 27718 5436 27770
rect 5140 27716 5196 27718
rect 5220 27716 5276 27718
rect 5300 27716 5356 27718
rect 5380 27716 5436 27718
rect 5800 27226 5856 27228
rect 5880 27226 5936 27228
rect 5960 27226 6016 27228
rect 6040 27226 6096 27228
rect 5800 27174 5846 27226
rect 5846 27174 5856 27226
rect 5880 27174 5910 27226
rect 5910 27174 5922 27226
rect 5922 27174 5936 27226
rect 5960 27174 5974 27226
rect 5974 27174 5986 27226
rect 5986 27174 6016 27226
rect 6040 27174 6050 27226
rect 6050 27174 6096 27226
rect 5800 27172 5856 27174
rect 5880 27172 5936 27174
rect 5960 27172 6016 27174
rect 6040 27172 6096 27174
rect 5140 26682 5196 26684
rect 5220 26682 5276 26684
rect 5300 26682 5356 26684
rect 5380 26682 5436 26684
rect 5140 26630 5186 26682
rect 5186 26630 5196 26682
rect 5220 26630 5250 26682
rect 5250 26630 5262 26682
rect 5262 26630 5276 26682
rect 5300 26630 5314 26682
rect 5314 26630 5326 26682
rect 5326 26630 5356 26682
rect 5380 26630 5390 26682
rect 5390 26630 5436 26682
rect 5140 26628 5196 26630
rect 5220 26628 5276 26630
rect 5300 26628 5356 26630
rect 5380 26628 5436 26630
rect 14554 36488 14610 36544
rect 5800 26138 5856 26140
rect 5880 26138 5936 26140
rect 5960 26138 6016 26140
rect 6040 26138 6096 26140
rect 5800 26086 5846 26138
rect 5846 26086 5856 26138
rect 5880 26086 5910 26138
rect 5910 26086 5922 26138
rect 5922 26086 5936 26138
rect 5960 26086 5974 26138
rect 5974 26086 5986 26138
rect 5986 26086 6016 26138
rect 6040 26086 6050 26138
rect 6050 26086 6096 26138
rect 5800 26084 5856 26086
rect 5880 26084 5936 26086
rect 5960 26084 6016 26086
rect 6040 26084 6096 26086
rect 5140 25594 5196 25596
rect 5220 25594 5276 25596
rect 5300 25594 5356 25596
rect 5380 25594 5436 25596
rect 5140 25542 5186 25594
rect 5186 25542 5196 25594
rect 5220 25542 5250 25594
rect 5250 25542 5262 25594
rect 5262 25542 5276 25594
rect 5300 25542 5314 25594
rect 5314 25542 5326 25594
rect 5326 25542 5356 25594
rect 5380 25542 5390 25594
rect 5390 25542 5436 25594
rect 5140 25540 5196 25542
rect 5220 25540 5276 25542
rect 5300 25540 5356 25542
rect 5380 25540 5436 25542
rect 5800 25050 5856 25052
rect 5880 25050 5936 25052
rect 5960 25050 6016 25052
rect 6040 25050 6096 25052
rect 5800 24998 5846 25050
rect 5846 24998 5856 25050
rect 5880 24998 5910 25050
rect 5910 24998 5922 25050
rect 5922 24998 5936 25050
rect 5960 24998 5974 25050
rect 5974 24998 5986 25050
rect 5986 24998 6016 25050
rect 6040 24998 6050 25050
rect 6050 24998 6096 25050
rect 5800 24996 5856 24998
rect 5880 24996 5936 24998
rect 5960 24996 6016 24998
rect 6040 24996 6096 24998
rect 5140 24506 5196 24508
rect 5220 24506 5276 24508
rect 5300 24506 5356 24508
rect 5380 24506 5436 24508
rect 5140 24454 5186 24506
rect 5186 24454 5196 24506
rect 5220 24454 5250 24506
rect 5250 24454 5262 24506
rect 5262 24454 5276 24506
rect 5300 24454 5314 24506
rect 5314 24454 5326 24506
rect 5326 24454 5356 24506
rect 5380 24454 5390 24506
rect 5390 24454 5436 24506
rect 5140 24452 5196 24454
rect 5220 24452 5276 24454
rect 5300 24452 5356 24454
rect 5380 24452 5436 24454
rect 5800 23962 5856 23964
rect 5880 23962 5936 23964
rect 5960 23962 6016 23964
rect 6040 23962 6096 23964
rect 5800 23910 5846 23962
rect 5846 23910 5856 23962
rect 5880 23910 5910 23962
rect 5910 23910 5922 23962
rect 5922 23910 5936 23962
rect 5960 23910 5974 23962
rect 5974 23910 5986 23962
rect 5986 23910 6016 23962
rect 6040 23910 6050 23962
rect 6050 23910 6096 23962
rect 5800 23908 5856 23910
rect 5880 23908 5936 23910
rect 5960 23908 6016 23910
rect 6040 23908 6096 23910
rect 5140 23418 5196 23420
rect 5220 23418 5276 23420
rect 5300 23418 5356 23420
rect 5380 23418 5436 23420
rect 5140 23366 5186 23418
rect 5186 23366 5196 23418
rect 5220 23366 5250 23418
rect 5250 23366 5262 23418
rect 5262 23366 5276 23418
rect 5300 23366 5314 23418
rect 5314 23366 5326 23418
rect 5326 23366 5356 23418
rect 5380 23366 5390 23418
rect 5390 23366 5436 23418
rect 5140 23364 5196 23366
rect 5220 23364 5276 23366
rect 5300 23364 5356 23366
rect 5380 23364 5436 23366
rect 5800 22874 5856 22876
rect 5880 22874 5936 22876
rect 5960 22874 6016 22876
rect 6040 22874 6096 22876
rect 5800 22822 5846 22874
rect 5846 22822 5856 22874
rect 5880 22822 5910 22874
rect 5910 22822 5922 22874
rect 5922 22822 5936 22874
rect 5960 22822 5974 22874
rect 5974 22822 5986 22874
rect 5986 22822 6016 22874
rect 6040 22822 6050 22874
rect 6050 22822 6096 22874
rect 5800 22820 5856 22822
rect 5880 22820 5936 22822
rect 5960 22820 6016 22822
rect 6040 22820 6096 22822
rect 5140 22330 5196 22332
rect 5220 22330 5276 22332
rect 5300 22330 5356 22332
rect 5380 22330 5436 22332
rect 5140 22278 5186 22330
rect 5186 22278 5196 22330
rect 5220 22278 5250 22330
rect 5250 22278 5262 22330
rect 5262 22278 5276 22330
rect 5300 22278 5314 22330
rect 5314 22278 5326 22330
rect 5326 22278 5356 22330
rect 5380 22278 5390 22330
rect 5390 22278 5436 22330
rect 5140 22276 5196 22278
rect 5220 22276 5276 22278
rect 5300 22276 5356 22278
rect 5380 22276 5436 22278
rect 5800 21786 5856 21788
rect 5880 21786 5936 21788
rect 5960 21786 6016 21788
rect 6040 21786 6096 21788
rect 5800 21734 5846 21786
rect 5846 21734 5856 21786
rect 5880 21734 5910 21786
rect 5910 21734 5922 21786
rect 5922 21734 5936 21786
rect 5960 21734 5974 21786
rect 5974 21734 5986 21786
rect 5986 21734 6016 21786
rect 6040 21734 6050 21786
rect 6050 21734 6096 21786
rect 5800 21732 5856 21734
rect 5880 21732 5936 21734
rect 5960 21732 6016 21734
rect 6040 21732 6096 21734
rect 5140 21242 5196 21244
rect 5220 21242 5276 21244
rect 5300 21242 5356 21244
rect 5380 21242 5436 21244
rect 5140 21190 5186 21242
rect 5186 21190 5196 21242
rect 5220 21190 5250 21242
rect 5250 21190 5262 21242
rect 5262 21190 5276 21242
rect 5300 21190 5314 21242
rect 5314 21190 5326 21242
rect 5326 21190 5356 21242
rect 5380 21190 5390 21242
rect 5390 21190 5436 21242
rect 5140 21188 5196 21190
rect 5220 21188 5276 21190
rect 5300 21188 5356 21190
rect 5380 21188 5436 21190
rect 5800 20698 5856 20700
rect 5880 20698 5936 20700
rect 5960 20698 6016 20700
rect 6040 20698 6096 20700
rect 5800 20646 5846 20698
rect 5846 20646 5856 20698
rect 5880 20646 5910 20698
rect 5910 20646 5922 20698
rect 5922 20646 5936 20698
rect 5960 20646 5974 20698
rect 5974 20646 5986 20698
rect 5986 20646 6016 20698
rect 6040 20646 6050 20698
rect 6050 20646 6096 20698
rect 5800 20644 5856 20646
rect 5880 20644 5936 20646
rect 5960 20644 6016 20646
rect 6040 20644 6096 20646
rect 5140 20154 5196 20156
rect 5220 20154 5276 20156
rect 5300 20154 5356 20156
rect 5380 20154 5436 20156
rect 5140 20102 5186 20154
rect 5186 20102 5196 20154
rect 5220 20102 5250 20154
rect 5250 20102 5262 20154
rect 5262 20102 5276 20154
rect 5300 20102 5314 20154
rect 5314 20102 5326 20154
rect 5326 20102 5356 20154
rect 5380 20102 5390 20154
rect 5390 20102 5436 20154
rect 5140 20100 5196 20102
rect 5220 20100 5276 20102
rect 5300 20100 5356 20102
rect 5380 20100 5436 20102
rect 5800 19610 5856 19612
rect 5880 19610 5936 19612
rect 5960 19610 6016 19612
rect 6040 19610 6096 19612
rect 5800 19558 5846 19610
rect 5846 19558 5856 19610
rect 5880 19558 5910 19610
rect 5910 19558 5922 19610
rect 5922 19558 5936 19610
rect 5960 19558 5974 19610
rect 5974 19558 5986 19610
rect 5986 19558 6016 19610
rect 6040 19558 6050 19610
rect 6050 19558 6096 19610
rect 5800 19556 5856 19558
rect 5880 19556 5936 19558
rect 5960 19556 6016 19558
rect 6040 19556 6096 19558
rect 5140 19066 5196 19068
rect 5220 19066 5276 19068
rect 5300 19066 5356 19068
rect 5380 19066 5436 19068
rect 5140 19014 5186 19066
rect 5186 19014 5196 19066
rect 5220 19014 5250 19066
rect 5250 19014 5262 19066
rect 5262 19014 5276 19066
rect 5300 19014 5314 19066
rect 5314 19014 5326 19066
rect 5326 19014 5356 19066
rect 5380 19014 5390 19066
rect 5390 19014 5436 19066
rect 5140 19012 5196 19014
rect 5220 19012 5276 19014
rect 5300 19012 5356 19014
rect 5380 19012 5436 19014
rect 5800 18522 5856 18524
rect 5880 18522 5936 18524
rect 5960 18522 6016 18524
rect 6040 18522 6096 18524
rect 5800 18470 5846 18522
rect 5846 18470 5856 18522
rect 5880 18470 5910 18522
rect 5910 18470 5922 18522
rect 5922 18470 5936 18522
rect 5960 18470 5974 18522
rect 5974 18470 5986 18522
rect 5986 18470 6016 18522
rect 6040 18470 6050 18522
rect 6050 18470 6096 18522
rect 5800 18468 5856 18470
rect 5880 18468 5936 18470
rect 5960 18468 6016 18470
rect 6040 18468 6096 18470
rect 5140 17978 5196 17980
rect 5220 17978 5276 17980
rect 5300 17978 5356 17980
rect 5380 17978 5436 17980
rect 5140 17926 5186 17978
rect 5186 17926 5196 17978
rect 5220 17926 5250 17978
rect 5250 17926 5262 17978
rect 5262 17926 5276 17978
rect 5300 17926 5314 17978
rect 5314 17926 5326 17978
rect 5326 17926 5356 17978
rect 5380 17926 5390 17978
rect 5390 17926 5436 17978
rect 5140 17924 5196 17926
rect 5220 17924 5276 17926
rect 5300 17924 5356 17926
rect 5380 17924 5436 17926
rect 5800 17434 5856 17436
rect 5880 17434 5936 17436
rect 5960 17434 6016 17436
rect 6040 17434 6096 17436
rect 5800 17382 5846 17434
rect 5846 17382 5856 17434
rect 5880 17382 5910 17434
rect 5910 17382 5922 17434
rect 5922 17382 5936 17434
rect 5960 17382 5974 17434
rect 5974 17382 5986 17434
rect 5986 17382 6016 17434
rect 6040 17382 6050 17434
rect 6050 17382 6096 17434
rect 5800 17380 5856 17382
rect 5880 17380 5936 17382
rect 5960 17380 6016 17382
rect 6040 17380 6096 17382
rect 5140 16890 5196 16892
rect 5220 16890 5276 16892
rect 5300 16890 5356 16892
rect 5380 16890 5436 16892
rect 5140 16838 5186 16890
rect 5186 16838 5196 16890
rect 5220 16838 5250 16890
rect 5250 16838 5262 16890
rect 5262 16838 5276 16890
rect 5300 16838 5314 16890
rect 5314 16838 5326 16890
rect 5326 16838 5356 16890
rect 5380 16838 5390 16890
rect 5390 16838 5436 16890
rect 5140 16836 5196 16838
rect 5220 16836 5276 16838
rect 5300 16836 5356 16838
rect 5380 16836 5436 16838
rect 5800 16346 5856 16348
rect 5880 16346 5936 16348
rect 5960 16346 6016 16348
rect 6040 16346 6096 16348
rect 5800 16294 5846 16346
rect 5846 16294 5856 16346
rect 5880 16294 5910 16346
rect 5910 16294 5922 16346
rect 5922 16294 5936 16346
rect 5960 16294 5974 16346
rect 5974 16294 5986 16346
rect 5986 16294 6016 16346
rect 6040 16294 6050 16346
rect 6050 16294 6096 16346
rect 5800 16292 5856 16294
rect 5880 16292 5936 16294
rect 5960 16292 6016 16294
rect 6040 16292 6096 16294
rect 5140 15802 5196 15804
rect 5220 15802 5276 15804
rect 5300 15802 5356 15804
rect 5380 15802 5436 15804
rect 5140 15750 5186 15802
rect 5186 15750 5196 15802
rect 5220 15750 5250 15802
rect 5250 15750 5262 15802
rect 5262 15750 5276 15802
rect 5300 15750 5314 15802
rect 5314 15750 5326 15802
rect 5326 15750 5356 15802
rect 5380 15750 5390 15802
rect 5390 15750 5436 15802
rect 5140 15748 5196 15750
rect 5220 15748 5276 15750
rect 5300 15748 5356 15750
rect 5380 15748 5436 15750
rect 5800 15258 5856 15260
rect 5880 15258 5936 15260
rect 5960 15258 6016 15260
rect 6040 15258 6096 15260
rect 5800 15206 5846 15258
rect 5846 15206 5856 15258
rect 5880 15206 5910 15258
rect 5910 15206 5922 15258
rect 5922 15206 5936 15258
rect 5960 15206 5974 15258
rect 5974 15206 5986 15258
rect 5986 15206 6016 15258
rect 6040 15206 6050 15258
rect 6050 15206 6096 15258
rect 5800 15204 5856 15206
rect 5880 15204 5936 15206
rect 5960 15204 6016 15206
rect 6040 15204 6096 15206
rect 5140 14714 5196 14716
rect 5220 14714 5276 14716
rect 5300 14714 5356 14716
rect 5380 14714 5436 14716
rect 5140 14662 5186 14714
rect 5186 14662 5196 14714
rect 5220 14662 5250 14714
rect 5250 14662 5262 14714
rect 5262 14662 5276 14714
rect 5300 14662 5314 14714
rect 5314 14662 5326 14714
rect 5326 14662 5356 14714
rect 5380 14662 5390 14714
rect 5390 14662 5436 14714
rect 5140 14660 5196 14662
rect 5220 14660 5276 14662
rect 5300 14660 5356 14662
rect 5380 14660 5436 14662
rect 5800 14170 5856 14172
rect 5880 14170 5936 14172
rect 5960 14170 6016 14172
rect 6040 14170 6096 14172
rect 5800 14118 5846 14170
rect 5846 14118 5856 14170
rect 5880 14118 5910 14170
rect 5910 14118 5922 14170
rect 5922 14118 5936 14170
rect 5960 14118 5974 14170
rect 5974 14118 5986 14170
rect 5986 14118 6016 14170
rect 6040 14118 6050 14170
rect 6050 14118 6096 14170
rect 5800 14116 5856 14118
rect 5880 14116 5936 14118
rect 5960 14116 6016 14118
rect 6040 14116 6096 14118
rect 5140 13626 5196 13628
rect 5220 13626 5276 13628
rect 5300 13626 5356 13628
rect 5380 13626 5436 13628
rect 5140 13574 5186 13626
rect 5186 13574 5196 13626
rect 5220 13574 5250 13626
rect 5250 13574 5262 13626
rect 5262 13574 5276 13626
rect 5300 13574 5314 13626
rect 5314 13574 5326 13626
rect 5326 13574 5356 13626
rect 5380 13574 5390 13626
rect 5390 13574 5436 13626
rect 5140 13572 5196 13574
rect 5220 13572 5276 13574
rect 5300 13572 5356 13574
rect 5380 13572 5436 13574
rect 5800 13082 5856 13084
rect 5880 13082 5936 13084
rect 5960 13082 6016 13084
rect 6040 13082 6096 13084
rect 5800 13030 5846 13082
rect 5846 13030 5856 13082
rect 5880 13030 5910 13082
rect 5910 13030 5922 13082
rect 5922 13030 5936 13082
rect 5960 13030 5974 13082
rect 5974 13030 5986 13082
rect 5986 13030 6016 13082
rect 6040 13030 6050 13082
rect 6050 13030 6096 13082
rect 5800 13028 5856 13030
rect 5880 13028 5936 13030
rect 5960 13028 6016 13030
rect 6040 13028 6096 13030
rect 5140 12538 5196 12540
rect 5220 12538 5276 12540
rect 5300 12538 5356 12540
rect 5380 12538 5436 12540
rect 5140 12486 5186 12538
rect 5186 12486 5196 12538
rect 5220 12486 5250 12538
rect 5250 12486 5262 12538
rect 5262 12486 5276 12538
rect 5300 12486 5314 12538
rect 5314 12486 5326 12538
rect 5326 12486 5356 12538
rect 5380 12486 5390 12538
rect 5390 12486 5436 12538
rect 5140 12484 5196 12486
rect 5220 12484 5276 12486
rect 5300 12484 5356 12486
rect 5380 12484 5436 12486
rect 5800 11994 5856 11996
rect 5880 11994 5936 11996
rect 5960 11994 6016 11996
rect 6040 11994 6096 11996
rect 5800 11942 5846 11994
rect 5846 11942 5856 11994
rect 5880 11942 5910 11994
rect 5910 11942 5922 11994
rect 5922 11942 5936 11994
rect 5960 11942 5974 11994
rect 5974 11942 5986 11994
rect 5986 11942 6016 11994
rect 6040 11942 6050 11994
rect 6050 11942 6096 11994
rect 5800 11940 5856 11942
rect 5880 11940 5936 11942
rect 5960 11940 6016 11942
rect 6040 11940 6096 11942
rect 5140 11450 5196 11452
rect 5220 11450 5276 11452
rect 5300 11450 5356 11452
rect 5380 11450 5436 11452
rect 5140 11398 5186 11450
rect 5186 11398 5196 11450
rect 5220 11398 5250 11450
rect 5250 11398 5262 11450
rect 5262 11398 5276 11450
rect 5300 11398 5314 11450
rect 5314 11398 5326 11450
rect 5326 11398 5356 11450
rect 5380 11398 5390 11450
rect 5390 11398 5436 11450
rect 5140 11396 5196 11398
rect 5220 11396 5276 11398
rect 5300 11396 5356 11398
rect 5380 11396 5436 11398
rect 5800 10906 5856 10908
rect 5880 10906 5936 10908
rect 5960 10906 6016 10908
rect 6040 10906 6096 10908
rect 5800 10854 5846 10906
rect 5846 10854 5856 10906
rect 5880 10854 5910 10906
rect 5910 10854 5922 10906
rect 5922 10854 5936 10906
rect 5960 10854 5974 10906
rect 5974 10854 5986 10906
rect 5986 10854 6016 10906
rect 6040 10854 6050 10906
rect 6050 10854 6096 10906
rect 5800 10852 5856 10854
rect 5880 10852 5936 10854
rect 5960 10852 6016 10854
rect 6040 10852 6096 10854
rect 5140 10362 5196 10364
rect 5220 10362 5276 10364
rect 5300 10362 5356 10364
rect 5380 10362 5436 10364
rect 5140 10310 5186 10362
rect 5186 10310 5196 10362
rect 5220 10310 5250 10362
rect 5250 10310 5262 10362
rect 5262 10310 5276 10362
rect 5300 10310 5314 10362
rect 5314 10310 5326 10362
rect 5326 10310 5356 10362
rect 5380 10310 5390 10362
rect 5390 10310 5436 10362
rect 5140 10308 5196 10310
rect 5220 10308 5276 10310
rect 5300 10308 5356 10310
rect 5380 10308 5436 10310
rect 5800 9818 5856 9820
rect 5880 9818 5936 9820
rect 5960 9818 6016 9820
rect 6040 9818 6096 9820
rect 5800 9766 5846 9818
rect 5846 9766 5856 9818
rect 5880 9766 5910 9818
rect 5910 9766 5922 9818
rect 5922 9766 5936 9818
rect 5960 9766 5974 9818
rect 5974 9766 5986 9818
rect 5986 9766 6016 9818
rect 6040 9766 6050 9818
rect 6050 9766 6096 9818
rect 5800 9764 5856 9766
rect 5880 9764 5936 9766
rect 5960 9764 6016 9766
rect 6040 9764 6096 9766
rect 5140 9274 5196 9276
rect 5220 9274 5276 9276
rect 5300 9274 5356 9276
rect 5380 9274 5436 9276
rect 5140 9222 5186 9274
rect 5186 9222 5196 9274
rect 5220 9222 5250 9274
rect 5250 9222 5262 9274
rect 5262 9222 5276 9274
rect 5300 9222 5314 9274
rect 5314 9222 5326 9274
rect 5326 9222 5356 9274
rect 5380 9222 5390 9274
rect 5390 9222 5436 9274
rect 5140 9220 5196 9222
rect 5220 9220 5276 9222
rect 5300 9220 5356 9222
rect 5380 9220 5436 9222
rect 5800 8730 5856 8732
rect 5880 8730 5936 8732
rect 5960 8730 6016 8732
rect 6040 8730 6096 8732
rect 5800 8678 5846 8730
rect 5846 8678 5856 8730
rect 5880 8678 5910 8730
rect 5910 8678 5922 8730
rect 5922 8678 5936 8730
rect 5960 8678 5974 8730
rect 5974 8678 5986 8730
rect 5986 8678 6016 8730
rect 6040 8678 6050 8730
rect 6050 8678 6096 8730
rect 5800 8676 5856 8678
rect 5880 8676 5936 8678
rect 5960 8676 6016 8678
rect 6040 8676 6096 8678
rect 5140 8186 5196 8188
rect 5220 8186 5276 8188
rect 5300 8186 5356 8188
rect 5380 8186 5436 8188
rect 5140 8134 5186 8186
rect 5186 8134 5196 8186
rect 5220 8134 5250 8186
rect 5250 8134 5262 8186
rect 5262 8134 5276 8186
rect 5300 8134 5314 8186
rect 5314 8134 5326 8186
rect 5326 8134 5356 8186
rect 5380 8134 5390 8186
rect 5390 8134 5436 8186
rect 5140 8132 5196 8134
rect 5220 8132 5276 8134
rect 5300 8132 5356 8134
rect 5380 8132 5436 8134
rect 5800 7642 5856 7644
rect 5880 7642 5936 7644
rect 5960 7642 6016 7644
rect 6040 7642 6096 7644
rect 5800 7590 5846 7642
rect 5846 7590 5856 7642
rect 5880 7590 5910 7642
rect 5910 7590 5922 7642
rect 5922 7590 5936 7642
rect 5960 7590 5974 7642
rect 5974 7590 5986 7642
rect 5986 7590 6016 7642
rect 6040 7590 6050 7642
rect 6050 7590 6096 7642
rect 5800 7588 5856 7590
rect 5880 7588 5936 7590
rect 5960 7588 6016 7590
rect 6040 7588 6096 7590
rect 5140 7098 5196 7100
rect 5220 7098 5276 7100
rect 5300 7098 5356 7100
rect 5380 7098 5436 7100
rect 5140 7046 5186 7098
rect 5186 7046 5196 7098
rect 5220 7046 5250 7098
rect 5250 7046 5262 7098
rect 5262 7046 5276 7098
rect 5300 7046 5314 7098
rect 5314 7046 5326 7098
rect 5326 7046 5356 7098
rect 5380 7046 5390 7098
rect 5390 7046 5436 7098
rect 5140 7044 5196 7046
rect 5220 7044 5276 7046
rect 5300 7044 5356 7046
rect 5380 7044 5436 7046
rect 5800 6554 5856 6556
rect 5880 6554 5936 6556
rect 5960 6554 6016 6556
rect 6040 6554 6096 6556
rect 5800 6502 5846 6554
rect 5846 6502 5856 6554
rect 5880 6502 5910 6554
rect 5910 6502 5922 6554
rect 5922 6502 5936 6554
rect 5960 6502 5974 6554
rect 5974 6502 5986 6554
rect 5986 6502 6016 6554
rect 6040 6502 6050 6554
rect 6050 6502 6096 6554
rect 5800 6500 5856 6502
rect 5880 6500 5936 6502
rect 5960 6500 6016 6502
rect 6040 6500 6096 6502
rect 5140 6010 5196 6012
rect 5220 6010 5276 6012
rect 5300 6010 5356 6012
rect 5380 6010 5436 6012
rect 5140 5958 5186 6010
rect 5186 5958 5196 6010
rect 5220 5958 5250 6010
rect 5250 5958 5262 6010
rect 5262 5958 5276 6010
rect 5300 5958 5314 6010
rect 5314 5958 5326 6010
rect 5326 5958 5356 6010
rect 5380 5958 5390 6010
rect 5390 5958 5436 6010
rect 5140 5956 5196 5958
rect 5220 5956 5276 5958
rect 5300 5956 5356 5958
rect 5380 5956 5436 5958
rect 5140 4922 5196 4924
rect 5220 4922 5276 4924
rect 5300 4922 5356 4924
rect 5380 4922 5436 4924
rect 5140 4870 5186 4922
rect 5186 4870 5196 4922
rect 5220 4870 5250 4922
rect 5250 4870 5262 4922
rect 5262 4870 5276 4922
rect 5300 4870 5314 4922
rect 5314 4870 5326 4922
rect 5326 4870 5356 4922
rect 5380 4870 5390 4922
rect 5390 4870 5436 4922
rect 5140 4868 5196 4870
rect 5220 4868 5276 4870
rect 5300 4868 5356 4870
rect 5380 4868 5436 4870
rect 5140 3834 5196 3836
rect 5220 3834 5276 3836
rect 5300 3834 5356 3836
rect 5380 3834 5436 3836
rect 5140 3782 5186 3834
rect 5186 3782 5196 3834
rect 5220 3782 5250 3834
rect 5250 3782 5262 3834
rect 5262 3782 5276 3834
rect 5300 3782 5314 3834
rect 5314 3782 5326 3834
rect 5326 3782 5356 3834
rect 5380 3782 5390 3834
rect 5390 3782 5436 3834
rect 5140 3780 5196 3782
rect 5220 3780 5276 3782
rect 5300 3780 5356 3782
rect 5380 3780 5436 3782
rect 5800 5466 5856 5468
rect 5880 5466 5936 5468
rect 5960 5466 6016 5468
rect 6040 5466 6096 5468
rect 5800 5414 5846 5466
rect 5846 5414 5856 5466
rect 5880 5414 5910 5466
rect 5910 5414 5922 5466
rect 5922 5414 5936 5466
rect 5960 5414 5974 5466
rect 5974 5414 5986 5466
rect 5986 5414 6016 5466
rect 6040 5414 6050 5466
rect 6050 5414 6096 5466
rect 5800 5412 5856 5414
rect 5880 5412 5936 5414
rect 5960 5412 6016 5414
rect 6040 5412 6096 5414
rect 5800 4378 5856 4380
rect 5880 4378 5936 4380
rect 5960 4378 6016 4380
rect 6040 4378 6096 4380
rect 5800 4326 5846 4378
rect 5846 4326 5856 4378
rect 5880 4326 5910 4378
rect 5910 4326 5922 4378
rect 5922 4326 5936 4378
rect 5960 4326 5974 4378
rect 5974 4326 5986 4378
rect 5986 4326 6016 4378
rect 6040 4326 6050 4378
rect 6050 4326 6096 4378
rect 5800 4324 5856 4326
rect 5880 4324 5936 4326
rect 5960 4324 6016 4326
rect 6040 4324 6096 4326
rect 5800 3290 5856 3292
rect 5880 3290 5936 3292
rect 5960 3290 6016 3292
rect 6040 3290 6096 3292
rect 5800 3238 5846 3290
rect 5846 3238 5856 3290
rect 5880 3238 5910 3290
rect 5910 3238 5922 3290
rect 5922 3238 5936 3290
rect 5960 3238 5974 3290
rect 5974 3238 5986 3290
rect 5986 3238 6016 3290
rect 6040 3238 6050 3290
rect 6050 3238 6096 3290
rect 5800 3236 5856 3238
rect 5880 3236 5936 3238
rect 5960 3236 6016 3238
rect 6040 3236 6096 3238
rect 5140 2746 5196 2748
rect 5220 2746 5276 2748
rect 5300 2746 5356 2748
rect 5380 2746 5436 2748
rect 5140 2694 5186 2746
rect 5186 2694 5196 2746
rect 5220 2694 5250 2746
rect 5250 2694 5262 2746
rect 5262 2694 5276 2746
rect 5300 2694 5314 2746
rect 5314 2694 5326 2746
rect 5326 2694 5356 2746
rect 5380 2694 5390 2746
rect 5390 2694 5436 2746
rect 5140 2692 5196 2694
rect 5220 2692 5276 2694
rect 5300 2692 5356 2694
rect 5380 2692 5436 2694
rect 4894 2352 4950 2408
rect 5630 2488 5686 2544
rect 6550 2624 6606 2680
rect 5800 2202 5856 2204
rect 5880 2202 5936 2204
rect 5960 2202 6016 2204
rect 6040 2202 6096 2204
rect 5800 2150 5846 2202
rect 5846 2150 5856 2202
rect 5880 2150 5910 2202
rect 5910 2150 5922 2202
rect 5922 2150 5936 2202
rect 5960 2150 5974 2202
rect 5974 2150 5986 2202
rect 5986 2150 6016 2202
rect 6040 2150 6050 2202
rect 6050 2150 6096 2202
rect 5800 2148 5856 2150
rect 5880 2148 5936 2150
rect 5960 2148 6016 2150
rect 6040 2148 6096 2150
rect 7838 4936 7894 4992
rect 8206 3188 8262 3224
rect 8206 3168 8208 3188
rect 8208 3168 8260 3188
rect 8260 3168 8262 3188
rect 11610 10648 11666 10704
rect 10414 8880 10470 8936
rect 9310 5344 9366 5400
rect 9494 3848 9550 3904
rect 10138 5208 10194 5264
rect 10046 4020 10048 4040
rect 10048 4020 10100 4040
rect 10100 4020 10102 4040
rect 10046 3984 10102 4020
rect 9954 3052 10010 3088
rect 9954 3032 9956 3052
rect 9956 3032 10008 3052
rect 10008 3032 10010 3052
rect 9034 1944 9090 2000
rect 6734 1264 6790 1320
rect 10598 4664 10654 4720
rect 10598 2216 10654 2272
rect 9126 40 9182 96
rect 10966 5616 11022 5672
rect 10966 3440 11022 3496
rect 11334 4664 11390 4720
rect 11242 3304 11298 3360
rect 32678 36352 32734 36408
rect 12254 8608 12310 8664
rect 12070 7268 12126 7304
rect 12070 7248 12072 7268
rect 12072 7248 12124 7268
rect 12124 7248 12126 7268
rect 11886 5888 11942 5944
rect 11518 3712 11574 3768
rect 11978 4664 12034 4720
rect 11978 4120 12034 4176
rect 12990 9288 13046 9344
rect 12254 4256 12310 4312
rect 12346 3304 12402 3360
rect 12622 3168 12678 3224
rect 12806 3712 12862 3768
rect 10966 1264 11022 1320
rect 13542 4684 13598 4720
rect 13542 4664 13544 4684
rect 13544 4664 13596 4684
rect 13596 4664 13598 4684
rect 13818 3068 13820 3088
rect 13820 3068 13872 3088
rect 13872 3068 13874 3088
rect 13818 3032 13874 3068
rect 14278 7112 14334 7168
rect 14278 5208 14334 5264
rect 14830 5772 14886 5808
rect 14830 5752 14832 5772
rect 14832 5752 14884 5772
rect 14884 5752 14886 5772
rect 15014 7792 15070 7848
rect 15014 5208 15070 5264
rect 14646 5108 14648 5128
rect 14648 5108 14700 5128
rect 14700 5108 14702 5128
rect 14646 5072 14702 5108
rect 15014 4392 15070 4448
rect 14738 4140 14794 4176
rect 14738 4120 14740 4140
rect 14740 4120 14792 4140
rect 14792 4120 14794 4140
rect 14646 3576 14702 3632
rect 15106 3576 15162 3632
rect 15382 6976 15438 7032
rect 15382 3848 15438 3904
rect 15106 3068 15108 3088
rect 15108 3068 15160 3088
rect 15160 3068 15162 3088
rect 15106 3032 15162 3068
rect 15566 5480 15622 5536
rect 15842 5480 15898 5536
rect 15842 5072 15898 5128
rect 15750 3884 15752 3904
rect 15752 3884 15804 3904
rect 15804 3884 15806 3904
rect 15750 3848 15806 3884
rect 17222 10104 17278 10160
rect 16302 5888 16358 5944
rect 16762 7268 16818 7304
rect 16762 7248 16764 7268
rect 16764 7248 16816 7268
rect 16816 7248 16818 7268
rect 16578 5616 16634 5672
rect 16486 4664 16542 4720
rect 16394 4256 16450 4312
rect 16302 3576 16358 3632
rect 16762 3984 16818 4040
rect 17130 5888 17186 5944
rect 17314 4120 17370 4176
rect 17314 3848 17370 3904
rect 17314 3304 17370 3360
rect 17314 3032 17370 3088
rect 17314 2080 17370 2136
rect 21730 11328 21786 11384
rect 22466 11328 22522 11384
rect 21822 10784 21878 10840
rect 17958 10512 18014 10568
rect 17958 9152 18014 9208
rect 18142 8508 18144 8528
rect 18144 8508 18196 8528
rect 18196 8508 18198 8528
rect 18142 8472 18198 8508
rect 17774 8200 17830 8256
rect 18142 8356 18198 8392
rect 18142 8336 18144 8356
rect 18144 8336 18196 8356
rect 18196 8336 18198 8356
rect 18050 6160 18106 6216
rect 17774 5752 17830 5808
rect 17498 5480 17554 5536
rect 17590 4664 17646 4720
rect 17866 4800 17922 4856
rect 17774 4664 17830 4720
rect 17682 4392 17738 4448
rect 17590 3984 17646 4040
rect 17774 4120 17830 4176
rect 17682 3304 17738 3360
rect 17498 2760 17554 2816
rect 18326 5344 18382 5400
rect 18142 4936 18198 4992
rect 18142 4664 18198 4720
rect 18602 8744 18658 8800
rect 18510 6568 18566 6624
rect 18510 6024 18566 6080
rect 18510 5480 18566 5536
rect 18142 3848 18198 3904
rect 19246 9152 19302 9208
rect 20442 10004 20444 10024
rect 20444 10004 20496 10024
rect 20496 10004 20498 10024
rect 19430 9288 19486 9344
rect 19430 8744 19486 8800
rect 19614 9696 19670 9752
rect 19246 6432 19302 6488
rect 19154 6024 19210 6080
rect 19338 6024 19394 6080
rect 19246 5616 19302 5672
rect 18694 1944 18750 2000
rect 19062 5344 19118 5400
rect 19154 5072 19210 5128
rect 20442 9968 20498 10004
rect 19522 3848 19578 3904
rect 19890 8336 19946 8392
rect 20350 8608 20406 8664
rect 20166 7520 20222 7576
rect 19890 6024 19946 6080
rect 20258 7112 20314 7168
rect 20534 8336 20590 8392
rect 19982 4276 20038 4312
rect 19982 4256 19984 4276
rect 19984 4256 20036 4276
rect 20036 4256 20038 4276
rect 19890 3984 19946 4040
rect 20442 5888 20498 5944
rect 20258 3712 20314 3768
rect 20166 3168 20222 3224
rect 20810 9868 20812 9888
rect 20812 9868 20864 9888
rect 20864 9868 20866 9888
rect 20810 9832 20866 9868
rect 21178 10240 21234 10296
rect 21178 8200 21234 8256
rect 22190 10376 22246 10432
rect 21822 9696 21878 9752
rect 20994 7656 21050 7712
rect 20810 5752 20866 5808
rect 20810 5616 20866 5672
rect 20902 5344 20958 5400
rect 20902 4392 20958 4448
rect 21178 7284 21180 7304
rect 21180 7284 21232 7304
rect 21232 7284 21234 7304
rect 21178 7248 21234 7284
rect 21454 7520 21510 7576
rect 21454 6568 21510 6624
rect 21362 6452 21418 6488
rect 21362 6432 21364 6452
rect 21364 6432 21416 6452
rect 21416 6432 21418 6452
rect 20718 2644 20774 2680
rect 20718 2624 20720 2644
rect 20720 2624 20772 2644
rect 20772 2624 20774 2644
rect 21086 2252 21088 2272
rect 21088 2252 21140 2272
rect 21140 2252 21142 2272
rect 21086 2216 21142 2252
rect 21362 5208 21418 5264
rect 21914 7112 21970 7168
rect 21822 5072 21878 5128
rect 21270 4800 21326 4856
rect 21362 4020 21364 4040
rect 21364 4020 21416 4040
rect 21416 4020 21418 4040
rect 21362 3984 21418 4020
rect 21730 4528 21786 4584
rect 21638 3848 21694 3904
rect 22742 11212 22798 11248
rect 22742 11192 22744 11212
rect 22744 11192 22796 11212
rect 22796 11192 22798 11212
rect 23202 11192 23258 11248
rect 22466 7420 22468 7440
rect 22468 7420 22520 7440
rect 22520 7420 22522 7440
rect 22466 7384 22522 7420
rect 22282 6976 22338 7032
rect 22190 6704 22246 6760
rect 22742 7928 22798 7984
rect 22558 6840 22614 6896
rect 22466 5480 22522 5536
rect 22190 4256 22246 4312
rect 22006 2488 22062 2544
rect 23386 11076 23442 11112
rect 23386 11056 23388 11076
rect 23388 11056 23440 11076
rect 23440 11056 23442 11076
rect 23018 8900 23074 8936
rect 23018 8880 23020 8900
rect 23020 8880 23072 8900
rect 23072 8880 23074 8900
rect 23018 5616 23074 5672
rect 23478 9968 23534 10024
rect 23294 6452 23350 6488
rect 23294 6432 23296 6452
rect 23296 6432 23348 6452
rect 23348 6432 23350 6452
rect 23202 4276 23258 4312
rect 23202 4256 23204 4276
rect 23204 4256 23256 4276
rect 23256 4256 23258 4276
rect 23386 5480 23442 5536
rect 23570 4800 23626 4856
rect 23754 7656 23810 7712
rect 23846 6976 23902 7032
rect 23754 6432 23810 6488
rect 24030 7248 24086 7304
rect 24030 6296 24086 6352
rect 24030 5888 24086 5944
rect 24214 9560 24270 9616
rect 25226 11500 25228 11520
rect 25228 11500 25280 11520
rect 25280 11500 25282 11520
rect 25226 11464 25282 11500
rect 24306 8744 24362 8800
rect 24398 8608 24454 8664
rect 22926 2624 22982 2680
rect 24306 7656 24362 7712
rect 24398 6452 24454 6488
rect 24398 6432 24400 6452
rect 24400 6432 24452 6452
rect 24452 6432 24454 6452
rect 24122 5616 24178 5672
rect 22834 1944 22890 2000
rect 24306 4936 24362 4992
rect 24306 4528 24362 4584
rect 24674 9696 24730 9752
rect 24858 9968 24914 10024
rect 24766 8200 24822 8256
rect 24766 7792 24822 7848
rect 25318 10784 25374 10840
rect 25042 7656 25098 7712
rect 24950 7520 25006 7576
rect 24674 6432 24730 6488
rect 24674 5344 24730 5400
rect 25134 5616 25190 5672
rect 24858 5228 24914 5264
rect 24858 5208 24860 5228
rect 24860 5208 24912 5228
rect 24912 5208 24914 5228
rect 24582 4120 24638 4176
rect 24950 3848 25006 3904
rect 24766 3576 24822 3632
rect 26054 11348 26110 11384
rect 26054 11328 26056 11348
rect 26056 11328 26108 11348
rect 26108 11328 26110 11348
rect 26238 11212 26294 11248
rect 26238 11192 26240 11212
rect 26240 11192 26292 11212
rect 26292 11192 26294 11212
rect 26054 10668 26110 10704
rect 26054 10648 26056 10668
rect 26056 10648 26108 10668
rect 26108 10648 26110 10668
rect 26330 9696 26386 9752
rect 25318 8336 25374 8392
rect 25502 6740 25504 6760
rect 25504 6740 25556 6760
rect 25556 6740 25558 6760
rect 25502 6704 25558 6740
rect 25502 5616 25558 5672
rect 25962 9460 25964 9480
rect 25964 9460 26016 9480
rect 26016 9460 26018 9480
rect 25962 9424 26018 9460
rect 25870 8880 25926 8936
rect 25870 8064 25926 8120
rect 25686 7656 25742 7712
rect 25778 6840 25834 6896
rect 25686 6024 25742 6080
rect 26146 7112 26202 7168
rect 25502 5364 25558 5400
rect 25502 5344 25504 5364
rect 25504 5344 25556 5364
rect 25556 5344 25558 5364
rect 25594 4256 25650 4312
rect 25594 3712 25650 3768
rect 25870 4392 25926 4448
rect 25686 3340 25688 3360
rect 25688 3340 25740 3360
rect 25740 3340 25742 3360
rect 25686 3304 25742 3340
rect 26606 6840 26662 6896
rect 26422 4684 26478 4720
rect 26422 4664 26424 4684
rect 26424 4664 26476 4684
rect 26476 4664 26478 4684
rect 26146 3848 26202 3904
rect 26146 3460 26202 3496
rect 26146 3440 26148 3460
rect 26148 3440 26200 3460
rect 26200 3440 26202 3460
rect 26330 3848 26386 3904
rect 27618 10104 27674 10160
rect 27710 9968 27766 10024
rect 27066 7928 27122 7984
rect 26974 3304 27030 3360
rect 27434 8608 27490 8664
rect 27434 8200 27490 8256
rect 28446 11636 28448 11656
rect 28448 11636 28500 11656
rect 28500 11636 28502 11656
rect 28446 11600 28502 11636
rect 27342 5772 27398 5808
rect 27342 5752 27344 5772
rect 27344 5752 27396 5772
rect 27396 5752 27398 5772
rect 27434 5616 27490 5672
rect 27618 5480 27674 5536
rect 27526 5072 27582 5128
rect 27618 4936 27674 4992
rect 27342 4256 27398 4312
rect 27342 2896 27398 2952
rect 27894 5480 27950 5536
rect 27986 4564 27988 4584
rect 27988 4564 28040 4584
rect 28040 4564 28042 4584
rect 27986 4528 28042 4564
rect 28446 8472 28502 8528
rect 28814 11872 28870 11928
rect 28814 10548 28816 10568
rect 28816 10548 28868 10568
rect 28868 10548 28870 10568
rect 28814 10512 28870 10548
rect 28446 8064 28502 8120
rect 28262 7248 28318 7304
rect 28538 6704 28594 6760
rect 28446 6296 28502 6352
rect 28630 6296 28686 6352
rect 28354 5208 28410 5264
rect 28262 2388 28264 2408
rect 28264 2388 28316 2408
rect 28316 2388 28318 2408
rect 28262 2352 28318 2388
rect 28998 9560 29054 9616
rect 28722 3476 28724 3496
rect 28724 3476 28776 3496
rect 28776 3476 28778 3496
rect 28722 3440 28778 3476
rect 28722 3168 28778 3224
rect 28538 2896 28594 2952
rect 28906 4936 28962 4992
rect 29090 5752 29146 5808
rect 28998 4528 29054 4584
rect 28906 3168 28962 3224
rect 29274 7520 29330 7576
rect 29550 10784 29606 10840
rect 29274 5072 29330 5128
rect 29734 6976 29790 7032
rect 29734 6704 29790 6760
rect 29550 5888 29606 5944
rect 29458 5772 29514 5808
rect 29458 5752 29460 5772
rect 29460 5752 29512 5772
rect 29512 5752 29514 5772
rect 29642 5616 29698 5672
rect 29642 4528 29698 4584
rect 29642 4120 29698 4176
rect 29918 7112 29974 7168
rect 29918 6024 29974 6080
rect 29458 3576 29514 3632
rect 27710 1536 27766 1592
rect 28354 1400 28410 1456
rect 29918 3304 29974 3360
rect 30470 11056 30526 11112
rect 30470 10376 30526 10432
rect 30378 10104 30434 10160
rect 30562 9868 30564 9888
rect 30564 9868 30616 9888
rect 30616 9868 30618 9888
rect 30562 9832 30618 9868
rect 30102 7384 30158 7440
rect 30102 5072 30158 5128
rect 30562 7928 30618 7984
rect 30470 7828 30472 7848
rect 30472 7828 30524 7848
rect 30524 7828 30526 7848
rect 30470 7792 30526 7828
rect 30378 7112 30434 7168
rect 30746 6840 30802 6896
rect 29366 1400 29422 1456
rect 31114 9424 31170 9480
rect 30930 6568 30986 6624
rect 30838 5208 30894 5264
rect 30930 3848 30986 3904
rect 30930 3712 30986 3768
rect 31298 9152 31354 9208
rect 31298 6976 31354 7032
rect 31206 3712 31262 3768
rect 31574 9560 31630 9616
rect 31758 7520 31814 7576
rect 31574 6976 31630 7032
rect 31666 6432 31722 6488
rect 31758 6024 31814 6080
rect 31666 5752 31722 5808
rect 31666 5480 31722 5536
rect 31942 8064 31998 8120
rect 31942 7792 31998 7848
rect 31942 7112 31998 7168
rect 31942 6160 31998 6216
rect 35860 37562 35916 37564
rect 35940 37562 35996 37564
rect 36020 37562 36076 37564
rect 36100 37562 36156 37564
rect 35860 37510 35906 37562
rect 35906 37510 35916 37562
rect 35940 37510 35970 37562
rect 35970 37510 35982 37562
rect 35982 37510 35996 37562
rect 36020 37510 36034 37562
rect 36034 37510 36046 37562
rect 36046 37510 36076 37562
rect 36100 37510 36110 37562
rect 36110 37510 36156 37562
rect 35860 37508 35916 37510
rect 35940 37508 35996 37510
rect 36020 37508 36076 37510
rect 36100 37508 36156 37510
rect 36520 37018 36576 37020
rect 36600 37018 36656 37020
rect 36680 37018 36736 37020
rect 36760 37018 36816 37020
rect 36520 36966 36566 37018
rect 36566 36966 36576 37018
rect 36600 36966 36630 37018
rect 36630 36966 36642 37018
rect 36642 36966 36656 37018
rect 36680 36966 36694 37018
rect 36694 36966 36706 37018
rect 36706 36966 36736 37018
rect 36760 36966 36770 37018
rect 36770 36966 36816 37018
rect 36520 36964 36576 36966
rect 36600 36964 36656 36966
rect 36680 36964 36736 36966
rect 36760 36964 36816 36966
rect 32218 8628 32274 8664
rect 32218 8608 32220 8628
rect 32220 8608 32272 8628
rect 32272 8608 32274 8628
rect 32218 7404 32274 7440
rect 32218 7384 32220 7404
rect 32220 7384 32272 7404
rect 32272 7384 32274 7404
rect 32218 7112 32274 7168
rect 32034 5480 32090 5536
rect 30746 2896 30802 2952
rect 31390 2760 31446 2816
rect 25042 176 25098 232
rect 32494 8336 32550 8392
rect 32770 9696 32826 9752
rect 32402 6976 32458 7032
rect 32586 5652 32588 5672
rect 32588 5652 32640 5672
rect 32640 5652 32642 5672
rect 32586 5616 32642 5652
rect 33322 10920 33378 10976
rect 33230 9560 33286 9616
rect 33138 8880 33194 8936
rect 33046 8472 33102 8528
rect 33230 8472 33286 8528
rect 33046 7112 33102 7168
rect 32954 5480 33010 5536
rect 33598 10140 33600 10160
rect 33600 10140 33652 10160
rect 33652 10140 33654 10160
rect 33598 10104 33654 10140
rect 33690 9152 33746 9208
rect 33414 8336 33470 8392
rect 33414 7384 33470 7440
rect 33322 7112 33378 7168
rect 32770 2896 32826 2952
rect 33138 4548 33194 4584
rect 33138 4528 33140 4548
rect 33140 4528 33192 4548
rect 33192 4528 33194 4548
rect 33046 2896 33102 2952
rect 34242 9696 34298 9752
rect 33966 9152 34022 9208
rect 33874 7520 33930 7576
rect 33874 7112 33930 7168
rect 34242 8064 34298 8120
rect 34334 7928 34390 7984
rect 34610 9036 34666 9072
rect 34610 9016 34612 9036
rect 34612 9016 34664 9036
rect 34664 9016 34666 9036
rect 34334 6976 34390 7032
rect 34150 6568 34206 6624
rect 34518 6296 34574 6352
rect 34426 5788 34428 5808
rect 34428 5788 34480 5808
rect 34480 5788 34482 5808
rect 34426 5752 34482 5788
rect 33874 3304 33930 3360
rect 34978 10532 35034 10568
rect 34978 10512 34980 10532
rect 34980 10512 35032 10532
rect 35032 10512 35034 10532
rect 34794 8200 34850 8256
rect 34794 7792 34850 7848
rect 34978 9288 35034 9344
rect 35162 9152 35218 9208
rect 35254 8916 35256 8936
rect 35256 8916 35308 8936
rect 35308 8916 35310 8936
rect 35254 8880 35310 8916
rect 35070 8608 35126 8664
rect 34978 7928 35034 7984
rect 34886 7248 34942 7304
rect 34794 5072 34850 5128
rect 34702 4936 34758 4992
rect 34702 4256 34758 4312
rect 34610 3576 34666 3632
rect 35860 36474 35916 36476
rect 35940 36474 35996 36476
rect 36020 36474 36076 36476
rect 36100 36474 36156 36476
rect 35860 36422 35906 36474
rect 35906 36422 35916 36474
rect 35940 36422 35970 36474
rect 35970 36422 35982 36474
rect 35982 36422 35996 36474
rect 36020 36422 36034 36474
rect 36034 36422 36046 36474
rect 36046 36422 36076 36474
rect 36100 36422 36110 36474
rect 36110 36422 36156 36474
rect 35860 36420 35916 36422
rect 35940 36420 35996 36422
rect 36020 36420 36076 36422
rect 36100 36420 36156 36422
rect 36520 35930 36576 35932
rect 36600 35930 36656 35932
rect 36680 35930 36736 35932
rect 36760 35930 36816 35932
rect 36520 35878 36566 35930
rect 36566 35878 36576 35930
rect 36600 35878 36630 35930
rect 36630 35878 36642 35930
rect 36642 35878 36656 35930
rect 36680 35878 36694 35930
rect 36694 35878 36706 35930
rect 36706 35878 36736 35930
rect 36760 35878 36770 35930
rect 36770 35878 36816 35930
rect 36520 35876 36576 35878
rect 36600 35876 36656 35878
rect 36680 35876 36736 35878
rect 36760 35876 36816 35878
rect 35860 35386 35916 35388
rect 35940 35386 35996 35388
rect 36020 35386 36076 35388
rect 36100 35386 36156 35388
rect 35860 35334 35906 35386
rect 35906 35334 35916 35386
rect 35940 35334 35970 35386
rect 35970 35334 35982 35386
rect 35982 35334 35996 35386
rect 36020 35334 36034 35386
rect 36034 35334 36046 35386
rect 36046 35334 36076 35386
rect 36100 35334 36110 35386
rect 36110 35334 36156 35386
rect 35860 35332 35916 35334
rect 35940 35332 35996 35334
rect 36020 35332 36076 35334
rect 36100 35332 36156 35334
rect 36520 34842 36576 34844
rect 36600 34842 36656 34844
rect 36680 34842 36736 34844
rect 36760 34842 36816 34844
rect 36520 34790 36566 34842
rect 36566 34790 36576 34842
rect 36600 34790 36630 34842
rect 36630 34790 36642 34842
rect 36642 34790 36656 34842
rect 36680 34790 36694 34842
rect 36694 34790 36706 34842
rect 36706 34790 36736 34842
rect 36760 34790 36770 34842
rect 36770 34790 36816 34842
rect 36520 34788 36576 34790
rect 36600 34788 36656 34790
rect 36680 34788 36736 34790
rect 36760 34788 36816 34790
rect 35860 34298 35916 34300
rect 35940 34298 35996 34300
rect 36020 34298 36076 34300
rect 36100 34298 36156 34300
rect 35860 34246 35906 34298
rect 35906 34246 35916 34298
rect 35940 34246 35970 34298
rect 35970 34246 35982 34298
rect 35982 34246 35996 34298
rect 36020 34246 36034 34298
rect 36034 34246 36046 34298
rect 36046 34246 36076 34298
rect 36100 34246 36110 34298
rect 36110 34246 36156 34298
rect 35860 34244 35916 34246
rect 35940 34244 35996 34246
rect 36020 34244 36076 34246
rect 36100 34244 36156 34246
rect 36520 33754 36576 33756
rect 36600 33754 36656 33756
rect 36680 33754 36736 33756
rect 36760 33754 36816 33756
rect 36520 33702 36566 33754
rect 36566 33702 36576 33754
rect 36600 33702 36630 33754
rect 36630 33702 36642 33754
rect 36642 33702 36656 33754
rect 36680 33702 36694 33754
rect 36694 33702 36706 33754
rect 36706 33702 36736 33754
rect 36760 33702 36770 33754
rect 36770 33702 36816 33754
rect 36520 33700 36576 33702
rect 36600 33700 36656 33702
rect 36680 33700 36736 33702
rect 36760 33700 36816 33702
rect 35860 33210 35916 33212
rect 35940 33210 35996 33212
rect 36020 33210 36076 33212
rect 36100 33210 36156 33212
rect 35860 33158 35906 33210
rect 35906 33158 35916 33210
rect 35940 33158 35970 33210
rect 35970 33158 35982 33210
rect 35982 33158 35996 33210
rect 36020 33158 36034 33210
rect 36034 33158 36046 33210
rect 36046 33158 36076 33210
rect 36100 33158 36110 33210
rect 36110 33158 36156 33210
rect 35860 33156 35916 33158
rect 35940 33156 35996 33158
rect 36020 33156 36076 33158
rect 36100 33156 36156 33158
rect 36520 32666 36576 32668
rect 36600 32666 36656 32668
rect 36680 32666 36736 32668
rect 36760 32666 36816 32668
rect 36520 32614 36566 32666
rect 36566 32614 36576 32666
rect 36600 32614 36630 32666
rect 36630 32614 36642 32666
rect 36642 32614 36656 32666
rect 36680 32614 36694 32666
rect 36694 32614 36706 32666
rect 36706 32614 36736 32666
rect 36760 32614 36770 32666
rect 36770 32614 36816 32666
rect 36520 32612 36576 32614
rect 36600 32612 36656 32614
rect 36680 32612 36736 32614
rect 36760 32612 36816 32614
rect 35860 32122 35916 32124
rect 35940 32122 35996 32124
rect 36020 32122 36076 32124
rect 36100 32122 36156 32124
rect 35860 32070 35906 32122
rect 35906 32070 35916 32122
rect 35940 32070 35970 32122
rect 35970 32070 35982 32122
rect 35982 32070 35996 32122
rect 36020 32070 36034 32122
rect 36034 32070 36046 32122
rect 36046 32070 36076 32122
rect 36100 32070 36110 32122
rect 36110 32070 36156 32122
rect 35860 32068 35916 32070
rect 35940 32068 35996 32070
rect 36020 32068 36076 32070
rect 36100 32068 36156 32070
rect 36520 31578 36576 31580
rect 36600 31578 36656 31580
rect 36680 31578 36736 31580
rect 36760 31578 36816 31580
rect 36520 31526 36566 31578
rect 36566 31526 36576 31578
rect 36600 31526 36630 31578
rect 36630 31526 36642 31578
rect 36642 31526 36656 31578
rect 36680 31526 36694 31578
rect 36694 31526 36706 31578
rect 36706 31526 36736 31578
rect 36760 31526 36770 31578
rect 36770 31526 36816 31578
rect 36520 31524 36576 31526
rect 36600 31524 36656 31526
rect 36680 31524 36736 31526
rect 36760 31524 36816 31526
rect 35860 31034 35916 31036
rect 35940 31034 35996 31036
rect 36020 31034 36076 31036
rect 36100 31034 36156 31036
rect 35860 30982 35906 31034
rect 35906 30982 35916 31034
rect 35940 30982 35970 31034
rect 35970 30982 35982 31034
rect 35982 30982 35996 31034
rect 36020 30982 36034 31034
rect 36034 30982 36046 31034
rect 36046 30982 36076 31034
rect 36100 30982 36110 31034
rect 36110 30982 36156 31034
rect 35860 30980 35916 30982
rect 35940 30980 35996 30982
rect 36020 30980 36076 30982
rect 36100 30980 36156 30982
rect 36520 30490 36576 30492
rect 36600 30490 36656 30492
rect 36680 30490 36736 30492
rect 36760 30490 36816 30492
rect 36520 30438 36566 30490
rect 36566 30438 36576 30490
rect 36600 30438 36630 30490
rect 36630 30438 36642 30490
rect 36642 30438 36656 30490
rect 36680 30438 36694 30490
rect 36694 30438 36706 30490
rect 36706 30438 36736 30490
rect 36760 30438 36770 30490
rect 36770 30438 36816 30490
rect 36520 30436 36576 30438
rect 36600 30436 36656 30438
rect 36680 30436 36736 30438
rect 36760 30436 36816 30438
rect 35860 29946 35916 29948
rect 35940 29946 35996 29948
rect 36020 29946 36076 29948
rect 36100 29946 36156 29948
rect 35860 29894 35906 29946
rect 35906 29894 35916 29946
rect 35940 29894 35970 29946
rect 35970 29894 35982 29946
rect 35982 29894 35996 29946
rect 36020 29894 36034 29946
rect 36034 29894 36046 29946
rect 36046 29894 36076 29946
rect 36100 29894 36110 29946
rect 36110 29894 36156 29946
rect 35860 29892 35916 29894
rect 35940 29892 35996 29894
rect 36020 29892 36076 29894
rect 36100 29892 36156 29894
rect 36520 29402 36576 29404
rect 36600 29402 36656 29404
rect 36680 29402 36736 29404
rect 36760 29402 36816 29404
rect 36520 29350 36566 29402
rect 36566 29350 36576 29402
rect 36600 29350 36630 29402
rect 36630 29350 36642 29402
rect 36642 29350 36656 29402
rect 36680 29350 36694 29402
rect 36694 29350 36706 29402
rect 36706 29350 36736 29402
rect 36760 29350 36770 29402
rect 36770 29350 36816 29402
rect 36520 29348 36576 29350
rect 36600 29348 36656 29350
rect 36680 29348 36736 29350
rect 36760 29348 36816 29350
rect 35860 28858 35916 28860
rect 35940 28858 35996 28860
rect 36020 28858 36076 28860
rect 36100 28858 36156 28860
rect 35860 28806 35906 28858
rect 35906 28806 35916 28858
rect 35940 28806 35970 28858
rect 35970 28806 35982 28858
rect 35982 28806 35996 28858
rect 36020 28806 36034 28858
rect 36034 28806 36046 28858
rect 36046 28806 36076 28858
rect 36100 28806 36110 28858
rect 36110 28806 36156 28858
rect 35860 28804 35916 28806
rect 35940 28804 35996 28806
rect 36020 28804 36076 28806
rect 36100 28804 36156 28806
rect 36520 28314 36576 28316
rect 36600 28314 36656 28316
rect 36680 28314 36736 28316
rect 36760 28314 36816 28316
rect 36520 28262 36566 28314
rect 36566 28262 36576 28314
rect 36600 28262 36630 28314
rect 36630 28262 36642 28314
rect 36642 28262 36656 28314
rect 36680 28262 36694 28314
rect 36694 28262 36706 28314
rect 36706 28262 36736 28314
rect 36760 28262 36770 28314
rect 36770 28262 36816 28314
rect 36520 28260 36576 28262
rect 36600 28260 36656 28262
rect 36680 28260 36736 28262
rect 36760 28260 36816 28262
rect 35860 27770 35916 27772
rect 35940 27770 35996 27772
rect 36020 27770 36076 27772
rect 36100 27770 36156 27772
rect 35860 27718 35906 27770
rect 35906 27718 35916 27770
rect 35940 27718 35970 27770
rect 35970 27718 35982 27770
rect 35982 27718 35996 27770
rect 36020 27718 36034 27770
rect 36034 27718 36046 27770
rect 36046 27718 36076 27770
rect 36100 27718 36110 27770
rect 36110 27718 36156 27770
rect 35860 27716 35916 27718
rect 35940 27716 35996 27718
rect 36020 27716 36076 27718
rect 36100 27716 36156 27718
rect 36520 27226 36576 27228
rect 36600 27226 36656 27228
rect 36680 27226 36736 27228
rect 36760 27226 36816 27228
rect 36520 27174 36566 27226
rect 36566 27174 36576 27226
rect 36600 27174 36630 27226
rect 36630 27174 36642 27226
rect 36642 27174 36656 27226
rect 36680 27174 36694 27226
rect 36694 27174 36706 27226
rect 36706 27174 36736 27226
rect 36760 27174 36770 27226
rect 36770 27174 36816 27226
rect 36520 27172 36576 27174
rect 36600 27172 36656 27174
rect 36680 27172 36736 27174
rect 36760 27172 36816 27174
rect 35860 26682 35916 26684
rect 35940 26682 35996 26684
rect 36020 26682 36076 26684
rect 36100 26682 36156 26684
rect 35860 26630 35906 26682
rect 35906 26630 35916 26682
rect 35940 26630 35970 26682
rect 35970 26630 35982 26682
rect 35982 26630 35996 26682
rect 36020 26630 36034 26682
rect 36034 26630 36046 26682
rect 36046 26630 36076 26682
rect 36100 26630 36110 26682
rect 36110 26630 36156 26682
rect 35860 26628 35916 26630
rect 35940 26628 35996 26630
rect 36020 26628 36076 26630
rect 36100 26628 36156 26630
rect 36520 26138 36576 26140
rect 36600 26138 36656 26140
rect 36680 26138 36736 26140
rect 36760 26138 36816 26140
rect 36520 26086 36566 26138
rect 36566 26086 36576 26138
rect 36600 26086 36630 26138
rect 36630 26086 36642 26138
rect 36642 26086 36656 26138
rect 36680 26086 36694 26138
rect 36694 26086 36706 26138
rect 36706 26086 36736 26138
rect 36760 26086 36770 26138
rect 36770 26086 36816 26138
rect 36520 26084 36576 26086
rect 36600 26084 36656 26086
rect 36680 26084 36736 26086
rect 36760 26084 36816 26086
rect 35860 25594 35916 25596
rect 35940 25594 35996 25596
rect 36020 25594 36076 25596
rect 36100 25594 36156 25596
rect 35860 25542 35906 25594
rect 35906 25542 35916 25594
rect 35940 25542 35970 25594
rect 35970 25542 35982 25594
rect 35982 25542 35996 25594
rect 36020 25542 36034 25594
rect 36034 25542 36046 25594
rect 36046 25542 36076 25594
rect 36100 25542 36110 25594
rect 36110 25542 36156 25594
rect 35860 25540 35916 25542
rect 35940 25540 35996 25542
rect 36020 25540 36076 25542
rect 36100 25540 36156 25542
rect 36520 25050 36576 25052
rect 36600 25050 36656 25052
rect 36680 25050 36736 25052
rect 36760 25050 36816 25052
rect 36520 24998 36566 25050
rect 36566 24998 36576 25050
rect 36600 24998 36630 25050
rect 36630 24998 36642 25050
rect 36642 24998 36656 25050
rect 36680 24998 36694 25050
rect 36694 24998 36706 25050
rect 36706 24998 36736 25050
rect 36760 24998 36770 25050
rect 36770 24998 36816 25050
rect 36520 24996 36576 24998
rect 36600 24996 36656 24998
rect 36680 24996 36736 24998
rect 36760 24996 36816 24998
rect 35860 24506 35916 24508
rect 35940 24506 35996 24508
rect 36020 24506 36076 24508
rect 36100 24506 36156 24508
rect 35860 24454 35906 24506
rect 35906 24454 35916 24506
rect 35940 24454 35970 24506
rect 35970 24454 35982 24506
rect 35982 24454 35996 24506
rect 36020 24454 36034 24506
rect 36034 24454 36046 24506
rect 36046 24454 36076 24506
rect 36100 24454 36110 24506
rect 36110 24454 36156 24506
rect 35860 24452 35916 24454
rect 35940 24452 35996 24454
rect 36020 24452 36076 24454
rect 36100 24452 36156 24454
rect 36520 23962 36576 23964
rect 36600 23962 36656 23964
rect 36680 23962 36736 23964
rect 36760 23962 36816 23964
rect 36520 23910 36566 23962
rect 36566 23910 36576 23962
rect 36600 23910 36630 23962
rect 36630 23910 36642 23962
rect 36642 23910 36656 23962
rect 36680 23910 36694 23962
rect 36694 23910 36706 23962
rect 36706 23910 36736 23962
rect 36760 23910 36770 23962
rect 36770 23910 36816 23962
rect 36520 23908 36576 23910
rect 36600 23908 36656 23910
rect 36680 23908 36736 23910
rect 36760 23908 36816 23910
rect 35860 23418 35916 23420
rect 35940 23418 35996 23420
rect 36020 23418 36076 23420
rect 36100 23418 36156 23420
rect 35860 23366 35906 23418
rect 35906 23366 35916 23418
rect 35940 23366 35970 23418
rect 35970 23366 35982 23418
rect 35982 23366 35996 23418
rect 36020 23366 36034 23418
rect 36034 23366 36046 23418
rect 36046 23366 36076 23418
rect 36100 23366 36110 23418
rect 36110 23366 36156 23418
rect 35860 23364 35916 23366
rect 35940 23364 35996 23366
rect 36020 23364 36076 23366
rect 36100 23364 36156 23366
rect 36520 22874 36576 22876
rect 36600 22874 36656 22876
rect 36680 22874 36736 22876
rect 36760 22874 36816 22876
rect 36520 22822 36566 22874
rect 36566 22822 36576 22874
rect 36600 22822 36630 22874
rect 36630 22822 36642 22874
rect 36642 22822 36656 22874
rect 36680 22822 36694 22874
rect 36694 22822 36706 22874
rect 36706 22822 36736 22874
rect 36760 22822 36770 22874
rect 36770 22822 36816 22874
rect 36520 22820 36576 22822
rect 36600 22820 36656 22822
rect 36680 22820 36736 22822
rect 36760 22820 36816 22822
rect 35860 22330 35916 22332
rect 35940 22330 35996 22332
rect 36020 22330 36076 22332
rect 36100 22330 36156 22332
rect 35860 22278 35906 22330
rect 35906 22278 35916 22330
rect 35940 22278 35970 22330
rect 35970 22278 35982 22330
rect 35982 22278 35996 22330
rect 36020 22278 36034 22330
rect 36034 22278 36046 22330
rect 36046 22278 36076 22330
rect 36100 22278 36110 22330
rect 36110 22278 36156 22330
rect 35860 22276 35916 22278
rect 35940 22276 35996 22278
rect 36020 22276 36076 22278
rect 36100 22276 36156 22278
rect 36520 21786 36576 21788
rect 36600 21786 36656 21788
rect 36680 21786 36736 21788
rect 36760 21786 36816 21788
rect 36520 21734 36566 21786
rect 36566 21734 36576 21786
rect 36600 21734 36630 21786
rect 36630 21734 36642 21786
rect 36642 21734 36656 21786
rect 36680 21734 36694 21786
rect 36694 21734 36706 21786
rect 36706 21734 36736 21786
rect 36760 21734 36770 21786
rect 36770 21734 36816 21786
rect 36520 21732 36576 21734
rect 36600 21732 36656 21734
rect 36680 21732 36736 21734
rect 36760 21732 36816 21734
rect 35860 21242 35916 21244
rect 35940 21242 35996 21244
rect 36020 21242 36076 21244
rect 36100 21242 36156 21244
rect 35860 21190 35906 21242
rect 35906 21190 35916 21242
rect 35940 21190 35970 21242
rect 35970 21190 35982 21242
rect 35982 21190 35996 21242
rect 36020 21190 36034 21242
rect 36034 21190 36046 21242
rect 36046 21190 36076 21242
rect 36100 21190 36110 21242
rect 36110 21190 36156 21242
rect 35860 21188 35916 21190
rect 35940 21188 35996 21190
rect 36020 21188 36076 21190
rect 36100 21188 36156 21190
rect 36520 20698 36576 20700
rect 36600 20698 36656 20700
rect 36680 20698 36736 20700
rect 36760 20698 36816 20700
rect 36520 20646 36566 20698
rect 36566 20646 36576 20698
rect 36600 20646 36630 20698
rect 36630 20646 36642 20698
rect 36642 20646 36656 20698
rect 36680 20646 36694 20698
rect 36694 20646 36706 20698
rect 36706 20646 36736 20698
rect 36760 20646 36770 20698
rect 36770 20646 36816 20698
rect 36520 20644 36576 20646
rect 36600 20644 36656 20646
rect 36680 20644 36736 20646
rect 36760 20644 36816 20646
rect 35860 20154 35916 20156
rect 35940 20154 35996 20156
rect 36020 20154 36076 20156
rect 36100 20154 36156 20156
rect 35860 20102 35906 20154
rect 35906 20102 35916 20154
rect 35940 20102 35970 20154
rect 35970 20102 35982 20154
rect 35982 20102 35996 20154
rect 36020 20102 36034 20154
rect 36034 20102 36046 20154
rect 36046 20102 36076 20154
rect 36100 20102 36110 20154
rect 36110 20102 36156 20154
rect 35860 20100 35916 20102
rect 35940 20100 35996 20102
rect 36020 20100 36076 20102
rect 36100 20100 36156 20102
rect 36520 19610 36576 19612
rect 36600 19610 36656 19612
rect 36680 19610 36736 19612
rect 36760 19610 36816 19612
rect 36520 19558 36566 19610
rect 36566 19558 36576 19610
rect 36600 19558 36630 19610
rect 36630 19558 36642 19610
rect 36642 19558 36656 19610
rect 36680 19558 36694 19610
rect 36694 19558 36706 19610
rect 36706 19558 36736 19610
rect 36760 19558 36770 19610
rect 36770 19558 36816 19610
rect 36520 19556 36576 19558
rect 36600 19556 36656 19558
rect 36680 19556 36736 19558
rect 36760 19556 36816 19558
rect 35860 19066 35916 19068
rect 35940 19066 35996 19068
rect 36020 19066 36076 19068
rect 36100 19066 36156 19068
rect 35860 19014 35906 19066
rect 35906 19014 35916 19066
rect 35940 19014 35970 19066
rect 35970 19014 35982 19066
rect 35982 19014 35996 19066
rect 36020 19014 36034 19066
rect 36034 19014 36046 19066
rect 36046 19014 36076 19066
rect 36100 19014 36110 19066
rect 36110 19014 36156 19066
rect 35860 19012 35916 19014
rect 35940 19012 35996 19014
rect 36020 19012 36076 19014
rect 36100 19012 36156 19014
rect 36520 18522 36576 18524
rect 36600 18522 36656 18524
rect 36680 18522 36736 18524
rect 36760 18522 36816 18524
rect 36520 18470 36566 18522
rect 36566 18470 36576 18522
rect 36600 18470 36630 18522
rect 36630 18470 36642 18522
rect 36642 18470 36656 18522
rect 36680 18470 36694 18522
rect 36694 18470 36706 18522
rect 36706 18470 36736 18522
rect 36760 18470 36770 18522
rect 36770 18470 36816 18522
rect 36520 18468 36576 18470
rect 36600 18468 36656 18470
rect 36680 18468 36736 18470
rect 36760 18468 36816 18470
rect 35860 17978 35916 17980
rect 35940 17978 35996 17980
rect 36020 17978 36076 17980
rect 36100 17978 36156 17980
rect 35860 17926 35906 17978
rect 35906 17926 35916 17978
rect 35940 17926 35970 17978
rect 35970 17926 35982 17978
rect 35982 17926 35996 17978
rect 36020 17926 36034 17978
rect 36034 17926 36046 17978
rect 36046 17926 36076 17978
rect 36100 17926 36110 17978
rect 36110 17926 36156 17978
rect 35860 17924 35916 17926
rect 35940 17924 35996 17926
rect 36020 17924 36076 17926
rect 36100 17924 36156 17926
rect 36520 17434 36576 17436
rect 36600 17434 36656 17436
rect 36680 17434 36736 17436
rect 36760 17434 36816 17436
rect 36520 17382 36566 17434
rect 36566 17382 36576 17434
rect 36600 17382 36630 17434
rect 36630 17382 36642 17434
rect 36642 17382 36656 17434
rect 36680 17382 36694 17434
rect 36694 17382 36706 17434
rect 36706 17382 36736 17434
rect 36760 17382 36770 17434
rect 36770 17382 36816 17434
rect 36520 17380 36576 17382
rect 36600 17380 36656 17382
rect 36680 17380 36736 17382
rect 36760 17380 36816 17382
rect 35860 16890 35916 16892
rect 35940 16890 35996 16892
rect 36020 16890 36076 16892
rect 36100 16890 36156 16892
rect 35860 16838 35906 16890
rect 35906 16838 35916 16890
rect 35940 16838 35970 16890
rect 35970 16838 35982 16890
rect 35982 16838 35996 16890
rect 36020 16838 36034 16890
rect 36034 16838 36046 16890
rect 36046 16838 36076 16890
rect 36100 16838 36110 16890
rect 36110 16838 36156 16890
rect 35860 16836 35916 16838
rect 35940 16836 35996 16838
rect 36020 16836 36076 16838
rect 36100 16836 36156 16838
rect 36520 16346 36576 16348
rect 36600 16346 36656 16348
rect 36680 16346 36736 16348
rect 36760 16346 36816 16348
rect 36520 16294 36566 16346
rect 36566 16294 36576 16346
rect 36600 16294 36630 16346
rect 36630 16294 36642 16346
rect 36642 16294 36656 16346
rect 36680 16294 36694 16346
rect 36694 16294 36706 16346
rect 36706 16294 36736 16346
rect 36760 16294 36770 16346
rect 36770 16294 36816 16346
rect 36520 16292 36576 16294
rect 36600 16292 36656 16294
rect 36680 16292 36736 16294
rect 36760 16292 36816 16294
rect 35860 15802 35916 15804
rect 35940 15802 35996 15804
rect 36020 15802 36076 15804
rect 36100 15802 36156 15804
rect 35860 15750 35906 15802
rect 35906 15750 35916 15802
rect 35940 15750 35970 15802
rect 35970 15750 35982 15802
rect 35982 15750 35996 15802
rect 36020 15750 36034 15802
rect 36034 15750 36046 15802
rect 36046 15750 36076 15802
rect 36100 15750 36110 15802
rect 36110 15750 36156 15802
rect 35860 15748 35916 15750
rect 35940 15748 35996 15750
rect 36020 15748 36076 15750
rect 36100 15748 36156 15750
rect 36520 15258 36576 15260
rect 36600 15258 36656 15260
rect 36680 15258 36736 15260
rect 36760 15258 36816 15260
rect 36520 15206 36566 15258
rect 36566 15206 36576 15258
rect 36600 15206 36630 15258
rect 36630 15206 36642 15258
rect 36642 15206 36656 15258
rect 36680 15206 36694 15258
rect 36694 15206 36706 15258
rect 36706 15206 36736 15258
rect 36760 15206 36770 15258
rect 36770 15206 36816 15258
rect 36520 15204 36576 15206
rect 36600 15204 36656 15206
rect 36680 15204 36736 15206
rect 36760 15204 36816 15206
rect 35860 14714 35916 14716
rect 35940 14714 35996 14716
rect 36020 14714 36076 14716
rect 36100 14714 36156 14716
rect 35860 14662 35906 14714
rect 35906 14662 35916 14714
rect 35940 14662 35970 14714
rect 35970 14662 35982 14714
rect 35982 14662 35996 14714
rect 36020 14662 36034 14714
rect 36034 14662 36046 14714
rect 36046 14662 36076 14714
rect 36100 14662 36110 14714
rect 36110 14662 36156 14714
rect 35860 14660 35916 14662
rect 35940 14660 35996 14662
rect 36020 14660 36076 14662
rect 36100 14660 36156 14662
rect 66580 37562 66636 37564
rect 66660 37562 66716 37564
rect 66740 37562 66796 37564
rect 66820 37562 66876 37564
rect 66580 37510 66626 37562
rect 66626 37510 66636 37562
rect 66660 37510 66690 37562
rect 66690 37510 66702 37562
rect 66702 37510 66716 37562
rect 66740 37510 66754 37562
rect 66754 37510 66766 37562
rect 66766 37510 66796 37562
rect 66820 37510 66830 37562
rect 66830 37510 66876 37562
rect 66580 37508 66636 37510
rect 66660 37508 66716 37510
rect 66740 37508 66796 37510
rect 66820 37508 66876 37510
rect 67240 37018 67296 37020
rect 67320 37018 67376 37020
rect 67400 37018 67456 37020
rect 67480 37018 67536 37020
rect 67240 36966 67286 37018
rect 67286 36966 67296 37018
rect 67320 36966 67350 37018
rect 67350 36966 67362 37018
rect 67362 36966 67376 37018
rect 67400 36966 67414 37018
rect 67414 36966 67426 37018
rect 67426 36966 67456 37018
rect 67480 36966 67490 37018
rect 67490 36966 67536 37018
rect 67240 36964 67296 36966
rect 67320 36964 67376 36966
rect 67400 36964 67456 36966
rect 67480 36964 67536 36966
rect 66580 36474 66636 36476
rect 66660 36474 66716 36476
rect 66740 36474 66796 36476
rect 66820 36474 66876 36476
rect 66580 36422 66626 36474
rect 66626 36422 66636 36474
rect 66660 36422 66690 36474
rect 66690 36422 66702 36474
rect 66702 36422 66716 36474
rect 66740 36422 66754 36474
rect 66754 36422 66766 36474
rect 66766 36422 66796 36474
rect 66820 36422 66830 36474
rect 66830 36422 66876 36474
rect 66580 36420 66636 36422
rect 66660 36420 66716 36422
rect 66740 36420 66796 36422
rect 66820 36420 66876 36422
rect 67240 35930 67296 35932
rect 67320 35930 67376 35932
rect 67400 35930 67456 35932
rect 67480 35930 67536 35932
rect 67240 35878 67286 35930
rect 67286 35878 67296 35930
rect 67320 35878 67350 35930
rect 67350 35878 67362 35930
rect 67362 35878 67376 35930
rect 67400 35878 67414 35930
rect 67414 35878 67426 35930
rect 67426 35878 67456 35930
rect 67480 35878 67490 35930
rect 67490 35878 67536 35930
rect 67240 35876 67296 35878
rect 67320 35876 67376 35878
rect 67400 35876 67456 35878
rect 67480 35876 67536 35878
rect 66580 35386 66636 35388
rect 66660 35386 66716 35388
rect 66740 35386 66796 35388
rect 66820 35386 66876 35388
rect 66580 35334 66626 35386
rect 66626 35334 66636 35386
rect 66660 35334 66690 35386
rect 66690 35334 66702 35386
rect 66702 35334 66716 35386
rect 66740 35334 66754 35386
rect 66754 35334 66766 35386
rect 66766 35334 66796 35386
rect 66820 35334 66830 35386
rect 66830 35334 66876 35386
rect 66580 35332 66636 35334
rect 66660 35332 66716 35334
rect 66740 35332 66796 35334
rect 66820 35332 66876 35334
rect 67240 34842 67296 34844
rect 67320 34842 67376 34844
rect 67400 34842 67456 34844
rect 67480 34842 67536 34844
rect 67240 34790 67286 34842
rect 67286 34790 67296 34842
rect 67320 34790 67350 34842
rect 67350 34790 67362 34842
rect 67362 34790 67376 34842
rect 67400 34790 67414 34842
rect 67414 34790 67426 34842
rect 67426 34790 67456 34842
rect 67480 34790 67490 34842
rect 67490 34790 67536 34842
rect 67240 34788 67296 34790
rect 67320 34788 67376 34790
rect 67400 34788 67456 34790
rect 67480 34788 67536 34790
rect 66580 34298 66636 34300
rect 66660 34298 66716 34300
rect 66740 34298 66796 34300
rect 66820 34298 66876 34300
rect 66580 34246 66626 34298
rect 66626 34246 66636 34298
rect 66660 34246 66690 34298
rect 66690 34246 66702 34298
rect 66702 34246 66716 34298
rect 66740 34246 66754 34298
rect 66754 34246 66766 34298
rect 66766 34246 66796 34298
rect 66820 34246 66830 34298
rect 66830 34246 66876 34298
rect 66580 34244 66636 34246
rect 66660 34244 66716 34246
rect 66740 34244 66796 34246
rect 66820 34244 66876 34246
rect 67240 33754 67296 33756
rect 67320 33754 67376 33756
rect 67400 33754 67456 33756
rect 67480 33754 67536 33756
rect 67240 33702 67286 33754
rect 67286 33702 67296 33754
rect 67320 33702 67350 33754
rect 67350 33702 67362 33754
rect 67362 33702 67376 33754
rect 67400 33702 67414 33754
rect 67414 33702 67426 33754
rect 67426 33702 67456 33754
rect 67480 33702 67490 33754
rect 67490 33702 67536 33754
rect 67240 33700 67296 33702
rect 67320 33700 67376 33702
rect 67400 33700 67456 33702
rect 67480 33700 67536 33702
rect 66580 33210 66636 33212
rect 66660 33210 66716 33212
rect 66740 33210 66796 33212
rect 66820 33210 66876 33212
rect 66580 33158 66626 33210
rect 66626 33158 66636 33210
rect 66660 33158 66690 33210
rect 66690 33158 66702 33210
rect 66702 33158 66716 33210
rect 66740 33158 66754 33210
rect 66754 33158 66766 33210
rect 66766 33158 66796 33210
rect 66820 33158 66830 33210
rect 66830 33158 66876 33210
rect 66580 33156 66636 33158
rect 66660 33156 66716 33158
rect 66740 33156 66796 33158
rect 66820 33156 66876 33158
rect 67240 32666 67296 32668
rect 67320 32666 67376 32668
rect 67400 32666 67456 32668
rect 67480 32666 67536 32668
rect 67240 32614 67286 32666
rect 67286 32614 67296 32666
rect 67320 32614 67350 32666
rect 67350 32614 67362 32666
rect 67362 32614 67376 32666
rect 67400 32614 67414 32666
rect 67414 32614 67426 32666
rect 67426 32614 67456 32666
rect 67480 32614 67490 32666
rect 67490 32614 67536 32666
rect 67240 32612 67296 32614
rect 67320 32612 67376 32614
rect 67400 32612 67456 32614
rect 67480 32612 67536 32614
rect 66580 32122 66636 32124
rect 66660 32122 66716 32124
rect 66740 32122 66796 32124
rect 66820 32122 66876 32124
rect 66580 32070 66626 32122
rect 66626 32070 66636 32122
rect 66660 32070 66690 32122
rect 66690 32070 66702 32122
rect 66702 32070 66716 32122
rect 66740 32070 66754 32122
rect 66754 32070 66766 32122
rect 66766 32070 66796 32122
rect 66820 32070 66830 32122
rect 66830 32070 66876 32122
rect 66580 32068 66636 32070
rect 66660 32068 66716 32070
rect 66740 32068 66796 32070
rect 66820 32068 66876 32070
rect 67240 31578 67296 31580
rect 67320 31578 67376 31580
rect 67400 31578 67456 31580
rect 67480 31578 67536 31580
rect 67240 31526 67286 31578
rect 67286 31526 67296 31578
rect 67320 31526 67350 31578
rect 67350 31526 67362 31578
rect 67362 31526 67376 31578
rect 67400 31526 67414 31578
rect 67414 31526 67426 31578
rect 67426 31526 67456 31578
rect 67480 31526 67490 31578
rect 67490 31526 67536 31578
rect 67240 31524 67296 31526
rect 67320 31524 67376 31526
rect 67400 31524 67456 31526
rect 67480 31524 67536 31526
rect 66580 31034 66636 31036
rect 66660 31034 66716 31036
rect 66740 31034 66796 31036
rect 66820 31034 66876 31036
rect 66580 30982 66626 31034
rect 66626 30982 66636 31034
rect 66660 30982 66690 31034
rect 66690 30982 66702 31034
rect 66702 30982 66716 31034
rect 66740 30982 66754 31034
rect 66754 30982 66766 31034
rect 66766 30982 66796 31034
rect 66820 30982 66830 31034
rect 66830 30982 66876 31034
rect 66580 30980 66636 30982
rect 66660 30980 66716 30982
rect 66740 30980 66796 30982
rect 66820 30980 66876 30982
rect 67240 30490 67296 30492
rect 67320 30490 67376 30492
rect 67400 30490 67456 30492
rect 67480 30490 67536 30492
rect 67240 30438 67286 30490
rect 67286 30438 67296 30490
rect 67320 30438 67350 30490
rect 67350 30438 67362 30490
rect 67362 30438 67376 30490
rect 67400 30438 67414 30490
rect 67414 30438 67426 30490
rect 67426 30438 67456 30490
rect 67480 30438 67490 30490
rect 67490 30438 67536 30490
rect 67240 30436 67296 30438
rect 67320 30436 67376 30438
rect 67400 30436 67456 30438
rect 67480 30436 67536 30438
rect 66580 29946 66636 29948
rect 66660 29946 66716 29948
rect 66740 29946 66796 29948
rect 66820 29946 66876 29948
rect 66580 29894 66626 29946
rect 66626 29894 66636 29946
rect 66660 29894 66690 29946
rect 66690 29894 66702 29946
rect 66702 29894 66716 29946
rect 66740 29894 66754 29946
rect 66754 29894 66766 29946
rect 66766 29894 66796 29946
rect 66820 29894 66830 29946
rect 66830 29894 66876 29946
rect 66580 29892 66636 29894
rect 66660 29892 66716 29894
rect 66740 29892 66796 29894
rect 66820 29892 66876 29894
rect 67240 29402 67296 29404
rect 67320 29402 67376 29404
rect 67400 29402 67456 29404
rect 67480 29402 67536 29404
rect 67240 29350 67286 29402
rect 67286 29350 67296 29402
rect 67320 29350 67350 29402
rect 67350 29350 67362 29402
rect 67362 29350 67376 29402
rect 67400 29350 67414 29402
rect 67414 29350 67426 29402
rect 67426 29350 67456 29402
rect 67480 29350 67490 29402
rect 67490 29350 67536 29402
rect 67240 29348 67296 29350
rect 67320 29348 67376 29350
rect 67400 29348 67456 29350
rect 67480 29348 67536 29350
rect 66580 28858 66636 28860
rect 66660 28858 66716 28860
rect 66740 28858 66796 28860
rect 66820 28858 66876 28860
rect 66580 28806 66626 28858
rect 66626 28806 66636 28858
rect 66660 28806 66690 28858
rect 66690 28806 66702 28858
rect 66702 28806 66716 28858
rect 66740 28806 66754 28858
rect 66754 28806 66766 28858
rect 66766 28806 66796 28858
rect 66820 28806 66830 28858
rect 66830 28806 66876 28858
rect 66580 28804 66636 28806
rect 66660 28804 66716 28806
rect 66740 28804 66796 28806
rect 66820 28804 66876 28806
rect 67240 28314 67296 28316
rect 67320 28314 67376 28316
rect 67400 28314 67456 28316
rect 67480 28314 67536 28316
rect 67240 28262 67286 28314
rect 67286 28262 67296 28314
rect 67320 28262 67350 28314
rect 67350 28262 67362 28314
rect 67362 28262 67376 28314
rect 67400 28262 67414 28314
rect 67414 28262 67426 28314
rect 67426 28262 67456 28314
rect 67480 28262 67490 28314
rect 67490 28262 67536 28314
rect 67240 28260 67296 28262
rect 67320 28260 67376 28262
rect 67400 28260 67456 28262
rect 67480 28260 67536 28262
rect 66580 27770 66636 27772
rect 66660 27770 66716 27772
rect 66740 27770 66796 27772
rect 66820 27770 66876 27772
rect 66580 27718 66626 27770
rect 66626 27718 66636 27770
rect 66660 27718 66690 27770
rect 66690 27718 66702 27770
rect 66702 27718 66716 27770
rect 66740 27718 66754 27770
rect 66754 27718 66766 27770
rect 66766 27718 66796 27770
rect 66820 27718 66830 27770
rect 66830 27718 66876 27770
rect 66580 27716 66636 27718
rect 66660 27716 66716 27718
rect 66740 27716 66796 27718
rect 66820 27716 66876 27718
rect 67240 27226 67296 27228
rect 67320 27226 67376 27228
rect 67400 27226 67456 27228
rect 67480 27226 67536 27228
rect 67240 27174 67286 27226
rect 67286 27174 67296 27226
rect 67320 27174 67350 27226
rect 67350 27174 67362 27226
rect 67362 27174 67376 27226
rect 67400 27174 67414 27226
rect 67414 27174 67426 27226
rect 67426 27174 67456 27226
rect 67480 27174 67490 27226
rect 67490 27174 67536 27226
rect 67240 27172 67296 27174
rect 67320 27172 67376 27174
rect 67400 27172 67456 27174
rect 67480 27172 67536 27174
rect 66580 26682 66636 26684
rect 66660 26682 66716 26684
rect 66740 26682 66796 26684
rect 66820 26682 66876 26684
rect 66580 26630 66626 26682
rect 66626 26630 66636 26682
rect 66660 26630 66690 26682
rect 66690 26630 66702 26682
rect 66702 26630 66716 26682
rect 66740 26630 66754 26682
rect 66754 26630 66766 26682
rect 66766 26630 66796 26682
rect 66820 26630 66830 26682
rect 66830 26630 66876 26682
rect 66580 26628 66636 26630
rect 66660 26628 66716 26630
rect 66740 26628 66796 26630
rect 66820 26628 66876 26630
rect 67240 26138 67296 26140
rect 67320 26138 67376 26140
rect 67400 26138 67456 26140
rect 67480 26138 67536 26140
rect 67240 26086 67286 26138
rect 67286 26086 67296 26138
rect 67320 26086 67350 26138
rect 67350 26086 67362 26138
rect 67362 26086 67376 26138
rect 67400 26086 67414 26138
rect 67414 26086 67426 26138
rect 67426 26086 67456 26138
rect 67480 26086 67490 26138
rect 67490 26086 67536 26138
rect 67240 26084 67296 26086
rect 67320 26084 67376 26086
rect 67400 26084 67456 26086
rect 67480 26084 67536 26086
rect 66580 25594 66636 25596
rect 66660 25594 66716 25596
rect 66740 25594 66796 25596
rect 66820 25594 66876 25596
rect 66580 25542 66626 25594
rect 66626 25542 66636 25594
rect 66660 25542 66690 25594
rect 66690 25542 66702 25594
rect 66702 25542 66716 25594
rect 66740 25542 66754 25594
rect 66754 25542 66766 25594
rect 66766 25542 66796 25594
rect 66820 25542 66830 25594
rect 66830 25542 66876 25594
rect 66580 25540 66636 25542
rect 66660 25540 66716 25542
rect 66740 25540 66796 25542
rect 66820 25540 66876 25542
rect 67240 25050 67296 25052
rect 67320 25050 67376 25052
rect 67400 25050 67456 25052
rect 67480 25050 67536 25052
rect 67240 24998 67286 25050
rect 67286 24998 67296 25050
rect 67320 24998 67350 25050
rect 67350 24998 67362 25050
rect 67362 24998 67376 25050
rect 67400 24998 67414 25050
rect 67414 24998 67426 25050
rect 67426 24998 67456 25050
rect 67480 24998 67490 25050
rect 67490 24998 67536 25050
rect 67240 24996 67296 24998
rect 67320 24996 67376 24998
rect 67400 24996 67456 24998
rect 67480 24996 67536 24998
rect 66580 24506 66636 24508
rect 66660 24506 66716 24508
rect 66740 24506 66796 24508
rect 66820 24506 66876 24508
rect 66580 24454 66626 24506
rect 66626 24454 66636 24506
rect 66660 24454 66690 24506
rect 66690 24454 66702 24506
rect 66702 24454 66716 24506
rect 66740 24454 66754 24506
rect 66754 24454 66766 24506
rect 66766 24454 66796 24506
rect 66820 24454 66830 24506
rect 66830 24454 66876 24506
rect 66580 24452 66636 24454
rect 66660 24452 66716 24454
rect 66740 24452 66796 24454
rect 66820 24452 66876 24454
rect 67240 23962 67296 23964
rect 67320 23962 67376 23964
rect 67400 23962 67456 23964
rect 67480 23962 67536 23964
rect 67240 23910 67286 23962
rect 67286 23910 67296 23962
rect 67320 23910 67350 23962
rect 67350 23910 67362 23962
rect 67362 23910 67376 23962
rect 67400 23910 67414 23962
rect 67414 23910 67426 23962
rect 67426 23910 67456 23962
rect 67480 23910 67490 23962
rect 67490 23910 67536 23962
rect 67240 23908 67296 23910
rect 67320 23908 67376 23910
rect 67400 23908 67456 23910
rect 67480 23908 67536 23910
rect 66580 23418 66636 23420
rect 66660 23418 66716 23420
rect 66740 23418 66796 23420
rect 66820 23418 66876 23420
rect 66580 23366 66626 23418
rect 66626 23366 66636 23418
rect 66660 23366 66690 23418
rect 66690 23366 66702 23418
rect 66702 23366 66716 23418
rect 66740 23366 66754 23418
rect 66754 23366 66766 23418
rect 66766 23366 66796 23418
rect 66820 23366 66830 23418
rect 66830 23366 66876 23418
rect 66580 23364 66636 23366
rect 66660 23364 66716 23366
rect 66740 23364 66796 23366
rect 66820 23364 66876 23366
rect 67240 22874 67296 22876
rect 67320 22874 67376 22876
rect 67400 22874 67456 22876
rect 67480 22874 67536 22876
rect 67240 22822 67286 22874
rect 67286 22822 67296 22874
rect 67320 22822 67350 22874
rect 67350 22822 67362 22874
rect 67362 22822 67376 22874
rect 67400 22822 67414 22874
rect 67414 22822 67426 22874
rect 67426 22822 67456 22874
rect 67480 22822 67490 22874
rect 67490 22822 67536 22874
rect 67240 22820 67296 22822
rect 67320 22820 67376 22822
rect 67400 22820 67456 22822
rect 67480 22820 67536 22822
rect 66580 22330 66636 22332
rect 66660 22330 66716 22332
rect 66740 22330 66796 22332
rect 66820 22330 66876 22332
rect 66580 22278 66626 22330
rect 66626 22278 66636 22330
rect 66660 22278 66690 22330
rect 66690 22278 66702 22330
rect 66702 22278 66716 22330
rect 66740 22278 66754 22330
rect 66754 22278 66766 22330
rect 66766 22278 66796 22330
rect 66820 22278 66830 22330
rect 66830 22278 66876 22330
rect 66580 22276 66636 22278
rect 66660 22276 66716 22278
rect 66740 22276 66796 22278
rect 66820 22276 66876 22278
rect 67240 21786 67296 21788
rect 67320 21786 67376 21788
rect 67400 21786 67456 21788
rect 67480 21786 67536 21788
rect 67240 21734 67286 21786
rect 67286 21734 67296 21786
rect 67320 21734 67350 21786
rect 67350 21734 67362 21786
rect 67362 21734 67376 21786
rect 67400 21734 67414 21786
rect 67414 21734 67426 21786
rect 67426 21734 67456 21786
rect 67480 21734 67490 21786
rect 67490 21734 67536 21786
rect 67240 21732 67296 21734
rect 67320 21732 67376 21734
rect 67400 21732 67456 21734
rect 67480 21732 67536 21734
rect 66580 21242 66636 21244
rect 66660 21242 66716 21244
rect 66740 21242 66796 21244
rect 66820 21242 66876 21244
rect 66580 21190 66626 21242
rect 66626 21190 66636 21242
rect 66660 21190 66690 21242
rect 66690 21190 66702 21242
rect 66702 21190 66716 21242
rect 66740 21190 66754 21242
rect 66754 21190 66766 21242
rect 66766 21190 66796 21242
rect 66820 21190 66830 21242
rect 66830 21190 66876 21242
rect 66580 21188 66636 21190
rect 66660 21188 66716 21190
rect 66740 21188 66796 21190
rect 66820 21188 66876 21190
rect 67240 20698 67296 20700
rect 67320 20698 67376 20700
rect 67400 20698 67456 20700
rect 67480 20698 67536 20700
rect 67240 20646 67286 20698
rect 67286 20646 67296 20698
rect 67320 20646 67350 20698
rect 67350 20646 67362 20698
rect 67362 20646 67376 20698
rect 67400 20646 67414 20698
rect 67414 20646 67426 20698
rect 67426 20646 67456 20698
rect 67480 20646 67490 20698
rect 67490 20646 67536 20698
rect 67240 20644 67296 20646
rect 67320 20644 67376 20646
rect 67400 20644 67456 20646
rect 67480 20644 67536 20646
rect 66580 20154 66636 20156
rect 66660 20154 66716 20156
rect 66740 20154 66796 20156
rect 66820 20154 66876 20156
rect 66580 20102 66626 20154
rect 66626 20102 66636 20154
rect 66660 20102 66690 20154
rect 66690 20102 66702 20154
rect 66702 20102 66716 20154
rect 66740 20102 66754 20154
rect 66754 20102 66766 20154
rect 66766 20102 66796 20154
rect 66820 20102 66830 20154
rect 66830 20102 66876 20154
rect 66580 20100 66636 20102
rect 66660 20100 66716 20102
rect 66740 20100 66796 20102
rect 66820 20100 66876 20102
rect 67240 19610 67296 19612
rect 67320 19610 67376 19612
rect 67400 19610 67456 19612
rect 67480 19610 67536 19612
rect 67240 19558 67286 19610
rect 67286 19558 67296 19610
rect 67320 19558 67350 19610
rect 67350 19558 67362 19610
rect 67362 19558 67376 19610
rect 67400 19558 67414 19610
rect 67414 19558 67426 19610
rect 67426 19558 67456 19610
rect 67480 19558 67490 19610
rect 67490 19558 67536 19610
rect 67240 19556 67296 19558
rect 67320 19556 67376 19558
rect 67400 19556 67456 19558
rect 67480 19556 67536 19558
rect 66580 19066 66636 19068
rect 66660 19066 66716 19068
rect 66740 19066 66796 19068
rect 66820 19066 66876 19068
rect 66580 19014 66626 19066
rect 66626 19014 66636 19066
rect 66660 19014 66690 19066
rect 66690 19014 66702 19066
rect 66702 19014 66716 19066
rect 66740 19014 66754 19066
rect 66754 19014 66766 19066
rect 66766 19014 66796 19066
rect 66820 19014 66830 19066
rect 66830 19014 66876 19066
rect 66580 19012 66636 19014
rect 66660 19012 66716 19014
rect 66740 19012 66796 19014
rect 66820 19012 66876 19014
rect 67240 18522 67296 18524
rect 67320 18522 67376 18524
rect 67400 18522 67456 18524
rect 67480 18522 67536 18524
rect 67240 18470 67286 18522
rect 67286 18470 67296 18522
rect 67320 18470 67350 18522
rect 67350 18470 67362 18522
rect 67362 18470 67376 18522
rect 67400 18470 67414 18522
rect 67414 18470 67426 18522
rect 67426 18470 67456 18522
rect 67480 18470 67490 18522
rect 67490 18470 67536 18522
rect 67240 18468 67296 18470
rect 67320 18468 67376 18470
rect 67400 18468 67456 18470
rect 67480 18468 67536 18470
rect 66580 17978 66636 17980
rect 66660 17978 66716 17980
rect 66740 17978 66796 17980
rect 66820 17978 66876 17980
rect 66580 17926 66626 17978
rect 66626 17926 66636 17978
rect 66660 17926 66690 17978
rect 66690 17926 66702 17978
rect 66702 17926 66716 17978
rect 66740 17926 66754 17978
rect 66754 17926 66766 17978
rect 66766 17926 66796 17978
rect 66820 17926 66830 17978
rect 66830 17926 66876 17978
rect 66580 17924 66636 17926
rect 66660 17924 66716 17926
rect 66740 17924 66796 17926
rect 66820 17924 66876 17926
rect 67240 17434 67296 17436
rect 67320 17434 67376 17436
rect 67400 17434 67456 17436
rect 67480 17434 67536 17436
rect 67240 17382 67286 17434
rect 67286 17382 67296 17434
rect 67320 17382 67350 17434
rect 67350 17382 67362 17434
rect 67362 17382 67376 17434
rect 67400 17382 67414 17434
rect 67414 17382 67426 17434
rect 67426 17382 67456 17434
rect 67480 17382 67490 17434
rect 67490 17382 67536 17434
rect 67240 17380 67296 17382
rect 67320 17380 67376 17382
rect 67400 17380 67456 17382
rect 67480 17380 67536 17382
rect 66580 16890 66636 16892
rect 66660 16890 66716 16892
rect 66740 16890 66796 16892
rect 66820 16890 66876 16892
rect 66580 16838 66626 16890
rect 66626 16838 66636 16890
rect 66660 16838 66690 16890
rect 66690 16838 66702 16890
rect 66702 16838 66716 16890
rect 66740 16838 66754 16890
rect 66754 16838 66766 16890
rect 66766 16838 66796 16890
rect 66820 16838 66830 16890
rect 66830 16838 66876 16890
rect 66580 16836 66636 16838
rect 66660 16836 66716 16838
rect 66740 16836 66796 16838
rect 66820 16836 66876 16838
rect 67240 16346 67296 16348
rect 67320 16346 67376 16348
rect 67400 16346 67456 16348
rect 67480 16346 67536 16348
rect 67240 16294 67286 16346
rect 67286 16294 67296 16346
rect 67320 16294 67350 16346
rect 67350 16294 67362 16346
rect 67362 16294 67376 16346
rect 67400 16294 67414 16346
rect 67414 16294 67426 16346
rect 67426 16294 67456 16346
rect 67480 16294 67490 16346
rect 67490 16294 67536 16346
rect 67240 16292 67296 16294
rect 67320 16292 67376 16294
rect 67400 16292 67456 16294
rect 67480 16292 67536 16294
rect 66580 15802 66636 15804
rect 66660 15802 66716 15804
rect 66740 15802 66796 15804
rect 66820 15802 66876 15804
rect 66580 15750 66626 15802
rect 66626 15750 66636 15802
rect 66660 15750 66690 15802
rect 66690 15750 66702 15802
rect 66702 15750 66716 15802
rect 66740 15750 66754 15802
rect 66754 15750 66766 15802
rect 66766 15750 66796 15802
rect 66820 15750 66830 15802
rect 66830 15750 66876 15802
rect 66580 15748 66636 15750
rect 66660 15748 66716 15750
rect 66740 15748 66796 15750
rect 66820 15748 66876 15750
rect 67240 15258 67296 15260
rect 67320 15258 67376 15260
rect 67400 15258 67456 15260
rect 67480 15258 67536 15260
rect 67240 15206 67286 15258
rect 67286 15206 67296 15258
rect 67320 15206 67350 15258
rect 67350 15206 67362 15258
rect 67362 15206 67376 15258
rect 67400 15206 67414 15258
rect 67414 15206 67426 15258
rect 67426 15206 67456 15258
rect 67480 15206 67490 15258
rect 67490 15206 67536 15258
rect 67240 15204 67296 15206
rect 67320 15204 67376 15206
rect 67400 15204 67456 15206
rect 67480 15204 67536 15206
rect 66580 14714 66636 14716
rect 66660 14714 66716 14716
rect 66740 14714 66796 14716
rect 66820 14714 66876 14716
rect 66580 14662 66626 14714
rect 66626 14662 66636 14714
rect 66660 14662 66690 14714
rect 66690 14662 66702 14714
rect 66702 14662 66716 14714
rect 66740 14662 66754 14714
rect 66754 14662 66766 14714
rect 66766 14662 66796 14714
rect 66820 14662 66830 14714
rect 66830 14662 66876 14714
rect 66580 14660 66636 14662
rect 66660 14660 66716 14662
rect 66740 14660 66796 14662
rect 66820 14660 66876 14662
rect 36520 14170 36576 14172
rect 36600 14170 36656 14172
rect 36680 14170 36736 14172
rect 36760 14170 36816 14172
rect 36520 14118 36566 14170
rect 36566 14118 36576 14170
rect 36600 14118 36630 14170
rect 36630 14118 36642 14170
rect 36642 14118 36656 14170
rect 36680 14118 36694 14170
rect 36694 14118 36706 14170
rect 36706 14118 36736 14170
rect 36760 14118 36770 14170
rect 36770 14118 36816 14170
rect 36520 14116 36576 14118
rect 36600 14116 36656 14118
rect 36680 14116 36736 14118
rect 36760 14116 36816 14118
rect 67240 14170 67296 14172
rect 67320 14170 67376 14172
rect 67400 14170 67456 14172
rect 67480 14170 67536 14172
rect 67240 14118 67286 14170
rect 67286 14118 67296 14170
rect 67320 14118 67350 14170
rect 67350 14118 67362 14170
rect 67362 14118 67376 14170
rect 67400 14118 67414 14170
rect 67414 14118 67426 14170
rect 67426 14118 67456 14170
rect 67480 14118 67490 14170
rect 67490 14118 67536 14170
rect 67240 14116 67296 14118
rect 67320 14116 67376 14118
rect 67400 14116 67456 14118
rect 67480 14116 67536 14118
rect 35860 13626 35916 13628
rect 35940 13626 35996 13628
rect 36020 13626 36076 13628
rect 36100 13626 36156 13628
rect 35860 13574 35906 13626
rect 35906 13574 35916 13626
rect 35940 13574 35970 13626
rect 35970 13574 35982 13626
rect 35982 13574 35996 13626
rect 36020 13574 36034 13626
rect 36034 13574 36046 13626
rect 36046 13574 36076 13626
rect 36100 13574 36110 13626
rect 36110 13574 36156 13626
rect 35860 13572 35916 13574
rect 35940 13572 35996 13574
rect 36020 13572 36076 13574
rect 36100 13572 36156 13574
rect 66580 13626 66636 13628
rect 66660 13626 66716 13628
rect 66740 13626 66796 13628
rect 66820 13626 66876 13628
rect 66580 13574 66626 13626
rect 66626 13574 66636 13626
rect 66660 13574 66690 13626
rect 66690 13574 66702 13626
rect 66702 13574 66716 13626
rect 66740 13574 66754 13626
rect 66754 13574 66766 13626
rect 66766 13574 66796 13626
rect 66820 13574 66830 13626
rect 66830 13574 66876 13626
rect 66580 13572 66636 13574
rect 66660 13572 66716 13574
rect 66740 13572 66796 13574
rect 66820 13572 66876 13574
rect 36520 13082 36576 13084
rect 36600 13082 36656 13084
rect 36680 13082 36736 13084
rect 36760 13082 36816 13084
rect 36520 13030 36566 13082
rect 36566 13030 36576 13082
rect 36600 13030 36630 13082
rect 36630 13030 36642 13082
rect 36642 13030 36656 13082
rect 36680 13030 36694 13082
rect 36694 13030 36706 13082
rect 36706 13030 36736 13082
rect 36760 13030 36770 13082
rect 36770 13030 36816 13082
rect 36520 13028 36576 13030
rect 36600 13028 36656 13030
rect 36680 13028 36736 13030
rect 36760 13028 36816 13030
rect 67240 13082 67296 13084
rect 67320 13082 67376 13084
rect 67400 13082 67456 13084
rect 67480 13082 67536 13084
rect 67240 13030 67286 13082
rect 67286 13030 67296 13082
rect 67320 13030 67350 13082
rect 67350 13030 67362 13082
rect 67362 13030 67376 13082
rect 67400 13030 67414 13082
rect 67414 13030 67426 13082
rect 67426 13030 67456 13082
rect 67480 13030 67490 13082
rect 67490 13030 67536 13082
rect 67240 13028 67296 13030
rect 67320 13028 67376 13030
rect 67400 13028 67456 13030
rect 67480 13028 67536 13030
rect 35860 12538 35916 12540
rect 35940 12538 35996 12540
rect 36020 12538 36076 12540
rect 36100 12538 36156 12540
rect 35860 12486 35906 12538
rect 35906 12486 35916 12538
rect 35940 12486 35970 12538
rect 35970 12486 35982 12538
rect 35982 12486 35996 12538
rect 36020 12486 36034 12538
rect 36034 12486 36046 12538
rect 36046 12486 36076 12538
rect 36100 12486 36110 12538
rect 36110 12486 36156 12538
rect 35860 12484 35916 12486
rect 35940 12484 35996 12486
rect 36020 12484 36076 12486
rect 36100 12484 36156 12486
rect 66580 12538 66636 12540
rect 66660 12538 66716 12540
rect 66740 12538 66796 12540
rect 66820 12538 66876 12540
rect 66580 12486 66626 12538
rect 66626 12486 66636 12538
rect 66660 12486 66690 12538
rect 66690 12486 66702 12538
rect 66702 12486 66716 12538
rect 66740 12486 66754 12538
rect 66754 12486 66766 12538
rect 66766 12486 66796 12538
rect 66820 12486 66830 12538
rect 66830 12486 66876 12538
rect 66580 12484 66636 12486
rect 66660 12484 66716 12486
rect 66740 12484 66796 12486
rect 66820 12484 66876 12486
rect 36520 11994 36576 11996
rect 36600 11994 36656 11996
rect 36680 11994 36736 11996
rect 36760 11994 36816 11996
rect 36520 11942 36566 11994
rect 36566 11942 36576 11994
rect 36600 11942 36630 11994
rect 36630 11942 36642 11994
rect 36642 11942 36656 11994
rect 36680 11942 36694 11994
rect 36694 11942 36706 11994
rect 36706 11942 36736 11994
rect 36760 11942 36770 11994
rect 36770 11942 36816 11994
rect 36520 11940 36576 11942
rect 36600 11940 36656 11942
rect 36680 11940 36736 11942
rect 36760 11940 36816 11942
rect 67240 11994 67296 11996
rect 67320 11994 67376 11996
rect 67400 11994 67456 11996
rect 67480 11994 67536 11996
rect 67240 11942 67286 11994
rect 67286 11942 67296 11994
rect 67320 11942 67350 11994
rect 67350 11942 67362 11994
rect 67362 11942 67376 11994
rect 67400 11942 67414 11994
rect 67414 11942 67426 11994
rect 67426 11942 67456 11994
rect 67480 11942 67490 11994
rect 67490 11942 67536 11994
rect 67240 11940 67296 11942
rect 67320 11940 67376 11942
rect 67400 11940 67456 11942
rect 67480 11940 67536 11942
rect 35860 11450 35916 11452
rect 35940 11450 35996 11452
rect 36020 11450 36076 11452
rect 36100 11450 36156 11452
rect 35860 11398 35906 11450
rect 35906 11398 35916 11450
rect 35940 11398 35970 11450
rect 35970 11398 35982 11450
rect 35982 11398 35996 11450
rect 36020 11398 36034 11450
rect 36034 11398 36046 11450
rect 36046 11398 36076 11450
rect 36100 11398 36110 11450
rect 36110 11398 36156 11450
rect 35860 11396 35916 11398
rect 35940 11396 35996 11398
rect 36020 11396 36076 11398
rect 36100 11396 36156 11398
rect 66580 11450 66636 11452
rect 66660 11450 66716 11452
rect 66740 11450 66796 11452
rect 66820 11450 66876 11452
rect 66580 11398 66626 11450
rect 66626 11398 66636 11450
rect 66660 11398 66690 11450
rect 66690 11398 66702 11450
rect 66702 11398 66716 11450
rect 66740 11398 66754 11450
rect 66754 11398 66766 11450
rect 66766 11398 66796 11450
rect 66820 11398 66830 11450
rect 66830 11398 66876 11450
rect 66580 11396 66636 11398
rect 66660 11396 66716 11398
rect 66740 11396 66796 11398
rect 66820 11396 66876 11398
rect 35530 8336 35586 8392
rect 36520 10906 36576 10908
rect 36600 10906 36656 10908
rect 36680 10906 36736 10908
rect 36760 10906 36816 10908
rect 36520 10854 36566 10906
rect 36566 10854 36576 10906
rect 36600 10854 36630 10906
rect 36630 10854 36642 10906
rect 36642 10854 36656 10906
rect 36680 10854 36694 10906
rect 36694 10854 36706 10906
rect 36706 10854 36736 10906
rect 36760 10854 36770 10906
rect 36770 10854 36816 10906
rect 36520 10852 36576 10854
rect 36600 10852 36656 10854
rect 36680 10852 36736 10854
rect 36760 10852 36816 10854
rect 35860 10362 35916 10364
rect 35940 10362 35996 10364
rect 36020 10362 36076 10364
rect 36100 10362 36156 10364
rect 35860 10310 35906 10362
rect 35906 10310 35916 10362
rect 35940 10310 35970 10362
rect 35970 10310 35982 10362
rect 35982 10310 35996 10362
rect 36020 10310 36034 10362
rect 36034 10310 36046 10362
rect 36046 10310 36076 10362
rect 36100 10310 36110 10362
rect 36110 10310 36156 10362
rect 35860 10308 35916 10310
rect 35940 10308 35996 10310
rect 36020 10308 36076 10310
rect 36100 10308 36156 10310
rect 36634 10004 36636 10024
rect 36636 10004 36688 10024
rect 36688 10004 36690 10024
rect 35898 9868 35900 9888
rect 35900 9868 35952 9888
rect 35952 9868 35954 9888
rect 35898 9832 35954 9868
rect 36634 9968 36690 10004
rect 36520 9818 36576 9820
rect 36600 9818 36656 9820
rect 36680 9818 36736 9820
rect 36760 9818 36816 9820
rect 36520 9766 36566 9818
rect 36566 9766 36576 9818
rect 36600 9766 36630 9818
rect 36630 9766 36642 9818
rect 36642 9766 36656 9818
rect 36680 9766 36694 9818
rect 36694 9766 36706 9818
rect 36706 9766 36736 9818
rect 36760 9766 36770 9818
rect 36770 9766 36816 9818
rect 36520 9764 36576 9766
rect 36600 9764 36656 9766
rect 36680 9764 36736 9766
rect 36760 9764 36816 9766
rect 36358 9424 36414 9480
rect 35860 9274 35916 9276
rect 35940 9274 35996 9276
rect 36020 9274 36076 9276
rect 36100 9274 36156 9276
rect 35860 9222 35906 9274
rect 35906 9222 35916 9274
rect 35940 9222 35970 9274
rect 35970 9222 35982 9274
rect 35982 9222 35996 9274
rect 36020 9222 36034 9274
rect 36034 9222 36046 9274
rect 36046 9222 36076 9274
rect 36100 9222 36110 9274
rect 36110 9222 36156 9274
rect 35860 9220 35916 9222
rect 35940 9220 35996 9222
rect 36020 9220 36076 9222
rect 36100 9220 36156 9222
rect 36266 8744 36322 8800
rect 35860 8186 35916 8188
rect 35940 8186 35996 8188
rect 36020 8186 36076 8188
rect 36100 8186 36156 8188
rect 35860 8134 35906 8186
rect 35906 8134 35916 8186
rect 35940 8134 35970 8186
rect 35970 8134 35982 8186
rect 35982 8134 35996 8186
rect 36020 8134 36034 8186
rect 36034 8134 36046 8186
rect 36046 8134 36076 8186
rect 36100 8134 36110 8186
rect 36110 8134 36156 8186
rect 35860 8132 35916 8134
rect 35940 8132 35996 8134
rect 36020 8132 36076 8134
rect 36100 8132 36156 8134
rect 35530 7540 35586 7576
rect 35530 7520 35532 7540
rect 35532 7520 35584 7540
rect 35584 7520 35586 7540
rect 35860 7098 35916 7100
rect 35940 7098 35996 7100
rect 36020 7098 36076 7100
rect 36100 7098 36156 7100
rect 35860 7046 35906 7098
rect 35906 7046 35916 7098
rect 35940 7046 35970 7098
rect 35970 7046 35982 7098
rect 35982 7046 35996 7098
rect 36020 7046 36034 7098
rect 36034 7046 36046 7098
rect 36046 7046 36076 7098
rect 36100 7046 36110 7098
rect 36110 7046 36156 7098
rect 35860 7044 35916 7046
rect 35940 7044 35996 7046
rect 36020 7044 36076 7046
rect 36100 7044 36156 7046
rect 35438 5480 35494 5536
rect 34978 4528 35034 4584
rect 35714 6024 35770 6080
rect 35860 6010 35916 6012
rect 35940 6010 35996 6012
rect 36020 6010 36076 6012
rect 36100 6010 36156 6012
rect 35860 5958 35906 6010
rect 35906 5958 35916 6010
rect 35940 5958 35970 6010
rect 35970 5958 35982 6010
rect 35982 5958 35996 6010
rect 36020 5958 36034 6010
rect 36034 5958 36046 6010
rect 36046 5958 36076 6010
rect 36100 5958 36110 6010
rect 36110 5958 36156 6010
rect 35860 5956 35916 5958
rect 35940 5956 35996 5958
rect 36020 5956 36076 5958
rect 36100 5956 36156 5958
rect 35714 5752 35770 5808
rect 36520 8730 36576 8732
rect 36600 8730 36656 8732
rect 36680 8730 36736 8732
rect 36760 8730 36816 8732
rect 36520 8678 36566 8730
rect 36566 8678 36576 8730
rect 36600 8678 36630 8730
rect 36630 8678 36642 8730
rect 36642 8678 36656 8730
rect 36680 8678 36694 8730
rect 36694 8678 36706 8730
rect 36706 8678 36736 8730
rect 36760 8678 36770 8730
rect 36770 8678 36816 8730
rect 36520 8676 36576 8678
rect 36600 8676 36656 8678
rect 36680 8676 36736 8678
rect 36760 8676 36816 8678
rect 36520 7642 36576 7644
rect 36600 7642 36656 7644
rect 36680 7642 36736 7644
rect 36760 7642 36816 7644
rect 36520 7590 36566 7642
rect 36566 7590 36576 7642
rect 36600 7590 36630 7642
rect 36630 7590 36642 7642
rect 36642 7590 36656 7642
rect 36680 7590 36694 7642
rect 36694 7590 36706 7642
rect 36706 7590 36736 7642
rect 36760 7590 36770 7642
rect 36770 7590 36816 7642
rect 36520 7588 36576 7590
rect 36600 7588 36656 7590
rect 36680 7588 36736 7590
rect 36760 7588 36816 7590
rect 36910 6840 36966 6896
rect 35898 5480 35954 5536
rect 35860 4922 35916 4924
rect 35940 4922 35996 4924
rect 36020 4922 36076 4924
rect 36100 4922 36156 4924
rect 35860 4870 35906 4922
rect 35906 4870 35916 4922
rect 35940 4870 35970 4922
rect 35970 4870 35982 4922
rect 35982 4870 35996 4922
rect 36020 4870 36034 4922
rect 36034 4870 36046 4922
rect 36046 4870 36076 4922
rect 36100 4870 36110 4922
rect 36110 4870 36156 4922
rect 35860 4868 35916 4870
rect 35940 4868 35996 4870
rect 36020 4868 36076 4870
rect 36100 4868 36156 4870
rect 36520 6554 36576 6556
rect 36600 6554 36656 6556
rect 36680 6554 36736 6556
rect 36760 6554 36816 6556
rect 36520 6502 36566 6554
rect 36566 6502 36576 6554
rect 36600 6502 36630 6554
rect 36630 6502 36642 6554
rect 36642 6502 36656 6554
rect 36680 6502 36694 6554
rect 36694 6502 36706 6554
rect 36706 6502 36736 6554
rect 36760 6502 36770 6554
rect 36770 6502 36816 6554
rect 36520 6500 36576 6502
rect 36600 6500 36656 6502
rect 36680 6500 36736 6502
rect 36760 6500 36816 6502
rect 36910 6160 36966 6216
rect 36450 5636 36506 5672
rect 36450 5616 36452 5636
rect 36452 5616 36504 5636
rect 36504 5616 36506 5636
rect 36520 5466 36576 5468
rect 36600 5466 36656 5468
rect 36680 5466 36736 5468
rect 36760 5466 36816 5468
rect 36520 5414 36566 5466
rect 36566 5414 36576 5466
rect 36600 5414 36630 5466
rect 36630 5414 36642 5466
rect 36642 5414 36656 5466
rect 36680 5414 36694 5466
rect 36694 5414 36706 5466
rect 36706 5414 36736 5466
rect 36760 5414 36770 5466
rect 36770 5414 36816 5466
rect 36520 5412 36576 5414
rect 36600 5412 36656 5414
rect 36680 5412 36736 5414
rect 36760 5412 36816 5414
rect 36450 4800 36506 4856
rect 36266 4120 36322 4176
rect 35860 3834 35916 3836
rect 35940 3834 35996 3836
rect 36020 3834 36076 3836
rect 36100 3834 36156 3836
rect 35860 3782 35906 3834
rect 35906 3782 35916 3834
rect 35940 3782 35970 3834
rect 35970 3782 35982 3834
rect 35982 3782 35996 3834
rect 36020 3782 36034 3834
rect 36034 3782 36046 3834
rect 36046 3782 36076 3834
rect 36100 3782 36110 3834
rect 36110 3782 36156 3834
rect 35860 3780 35916 3782
rect 35940 3780 35996 3782
rect 36020 3780 36076 3782
rect 36100 3780 36156 3782
rect 36520 4378 36576 4380
rect 36600 4378 36656 4380
rect 36680 4378 36736 4380
rect 36760 4378 36816 4380
rect 36520 4326 36566 4378
rect 36566 4326 36576 4378
rect 36600 4326 36630 4378
rect 36630 4326 36642 4378
rect 36642 4326 36656 4378
rect 36680 4326 36694 4378
rect 36694 4326 36706 4378
rect 36706 4326 36736 4378
rect 36760 4326 36770 4378
rect 36770 4326 36816 4378
rect 36520 4324 36576 4326
rect 36600 4324 36656 4326
rect 36680 4324 36736 4326
rect 36760 4324 36816 4326
rect 37370 5208 37426 5264
rect 36520 3290 36576 3292
rect 36600 3290 36656 3292
rect 36680 3290 36736 3292
rect 36760 3290 36816 3292
rect 36520 3238 36566 3290
rect 36566 3238 36576 3290
rect 36600 3238 36630 3290
rect 36630 3238 36642 3290
rect 36642 3238 36656 3290
rect 36680 3238 36694 3290
rect 36694 3238 36706 3290
rect 36706 3238 36736 3290
rect 36760 3238 36770 3290
rect 36770 3238 36816 3290
rect 36520 3236 36576 3238
rect 36600 3236 36656 3238
rect 36680 3236 36736 3238
rect 36760 3236 36816 3238
rect 35860 2746 35916 2748
rect 35940 2746 35996 2748
rect 36020 2746 36076 2748
rect 36100 2746 36156 2748
rect 35860 2694 35906 2746
rect 35906 2694 35916 2746
rect 35940 2694 35970 2746
rect 35970 2694 35982 2746
rect 35982 2694 35996 2746
rect 36020 2694 36034 2746
rect 36034 2694 36046 2746
rect 36046 2694 36076 2746
rect 36100 2694 36110 2746
rect 36110 2694 36156 2746
rect 35860 2692 35916 2694
rect 35940 2692 35996 2694
rect 36020 2692 36076 2694
rect 36100 2692 36156 2694
rect 35438 1264 35494 1320
rect 37554 3984 37610 4040
rect 36520 2202 36576 2204
rect 36600 2202 36656 2204
rect 36680 2202 36736 2204
rect 36760 2202 36816 2204
rect 36520 2150 36566 2202
rect 36566 2150 36576 2202
rect 36600 2150 36630 2202
rect 36630 2150 36642 2202
rect 36642 2150 36656 2202
rect 36680 2150 36694 2202
rect 36694 2150 36706 2202
rect 36706 2150 36736 2202
rect 36760 2150 36770 2202
rect 36770 2150 36816 2202
rect 36520 2148 36576 2150
rect 36600 2148 36656 2150
rect 36680 2148 36736 2150
rect 36760 2148 36816 2150
rect 38198 9016 38254 9072
rect 37738 5108 37740 5128
rect 37740 5108 37792 5128
rect 37792 5108 37794 5128
rect 37738 5072 37794 5108
rect 37738 4800 37794 4856
rect 37738 4020 37740 4040
rect 37740 4020 37792 4040
rect 37792 4020 37794 4040
rect 37738 3984 37794 4020
rect 38198 4800 38254 4856
rect 36726 1400 36782 1456
rect 37646 1400 37702 1456
rect 67240 10906 67296 10908
rect 67320 10906 67376 10908
rect 67400 10906 67456 10908
rect 67480 10906 67536 10908
rect 67240 10854 67286 10906
rect 67286 10854 67296 10906
rect 67320 10854 67350 10906
rect 67350 10854 67362 10906
rect 67362 10854 67376 10906
rect 67400 10854 67414 10906
rect 67414 10854 67426 10906
rect 67426 10854 67456 10906
rect 67480 10854 67490 10906
rect 67490 10854 67536 10906
rect 67240 10852 67296 10854
rect 67320 10852 67376 10854
rect 67400 10852 67456 10854
rect 67480 10852 67536 10854
rect 66580 10362 66636 10364
rect 66660 10362 66716 10364
rect 66740 10362 66796 10364
rect 66820 10362 66876 10364
rect 66580 10310 66626 10362
rect 66626 10310 66636 10362
rect 66660 10310 66690 10362
rect 66690 10310 66702 10362
rect 66702 10310 66716 10362
rect 66740 10310 66754 10362
rect 66754 10310 66766 10362
rect 66766 10310 66796 10362
rect 66820 10310 66830 10362
rect 66830 10310 66876 10362
rect 66580 10308 66636 10310
rect 66660 10308 66716 10310
rect 66740 10308 66796 10310
rect 66820 10308 66876 10310
rect 67240 9818 67296 9820
rect 67320 9818 67376 9820
rect 67400 9818 67456 9820
rect 67480 9818 67536 9820
rect 67240 9766 67286 9818
rect 67286 9766 67296 9818
rect 67320 9766 67350 9818
rect 67350 9766 67362 9818
rect 67362 9766 67376 9818
rect 67400 9766 67414 9818
rect 67414 9766 67426 9818
rect 67426 9766 67456 9818
rect 67480 9766 67490 9818
rect 67490 9766 67536 9818
rect 67240 9764 67296 9766
rect 67320 9764 67376 9766
rect 67400 9764 67456 9766
rect 67480 9764 67536 9766
rect 38474 3712 38530 3768
rect 66580 9274 66636 9276
rect 66660 9274 66716 9276
rect 66740 9274 66796 9276
rect 66820 9274 66876 9276
rect 66580 9222 66626 9274
rect 66626 9222 66636 9274
rect 66660 9222 66690 9274
rect 66690 9222 66702 9274
rect 66702 9222 66716 9274
rect 66740 9222 66754 9274
rect 66754 9222 66766 9274
rect 66766 9222 66796 9274
rect 66820 9222 66830 9274
rect 66830 9222 66876 9274
rect 66580 9220 66636 9222
rect 66660 9220 66716 9222
rect 66740 9220 66796 9222
rect 66820 9220 66876 9222
rect 67240 8730 67296 8732
rect 67320 8730 67376 8732
rect 67400 8730 67456 8732
rect 67480 8730 67536 8732
rect 67240 8678 67286 8730
rect 67286 8678 67296 8730
rect 67320 8678 67350 8730
rect 67350 8678 67362 8730
rect 67362 8678 67376 8730
rect 67400 8678 67414 8730
rect 67414 8678 67426 8730
rect 67426 8678 67456 8730
rect 67480 8678 67490 8730
rect 67490 8678 67536 8730
rect 67240 8676 67296 8678
rect 67320 8676 67376 8678
rect 67400 8676 67456 8678
rect 67480 8676 67536 8678
rect 40222 7928 40278 7984
rect 66580 8186 66636 8188
rect 66660 8186 66716 8188
rect 66740 8186 66796 8188
rect 66820 8186 66876 8188
rect 66580 8134 66626 8186
rect 66626 8134 66636 8186
rect 66660 8134 66690 8186
rect 66690 8134 66702 8186
rect 66702 8134 66716 8186
rect 66740 8134 66754 8186
rect 66754 8134 66766 8186
rect 66766 8134 66796 8186
rect 66820 8134 66830 8186
rect 66830 8134 66876 8186
rect 66580 8132 66636 8134
rect 66660 8132 66716 8134
rect 66740 8132 66796 8134
rect 66820 8132 66876 8134
rect 39946 5072 40002 5128
rect 41602 7812 41658 7848
rect 41602 7792 41604 7812
rect 41604 7792 41656 7812
rect 41656 7792 41658 7812
rect 40130 4664 40186 4720
rect 39946 4392 40002 4448
rect 40498 5072 40554 5128
rect 39946 3576 40002 3632
rect 39854 2896 39910 2952
rect 40498 3576 40554 3632
rect 40774 4256 40830 4312
rect 41326 3712 41382 3768
rect 41786 3848 41842 3904
rect 42522 3304 42578 3360
rect 42706 4528 42762 4584
rect 42706 4392 42762 4448
rect 42890 4256 42946 4312
rect 43258 3576 43314 3632
rect 43902 4120 43958 4176
rect 44178 3304 44234 3360
rect 44730 4020 44732 4040
rect 44732 4020 44784 4040
rect 44784 4020 44786 4040
rect 44730 3984 44786 4020
rect 67240 7642 67296 7644
rect 67320 7642 67376 7644
rect 67400 7642 67456 7644
rect 67480 7642 67536 7644
rect 67240 7590 67286 7642
rect 67286 7590 67296 7642
rect 67320 7590 67350 7642
rect 67350 7590 67362 7642
rect 67362 7590 67376 7642
rect 67400 7590 67414 7642
rect 67414 7590 67426 7642
rect 67426 7590 67456 7642
rect 67480 7590 67490 7642
rect 67490 7590 67536 7642
rect 67240 7588 67296 7590
rect 67320 7588 67376 7590
rect 67400 7588 67456 7590
rect 67480 7588 67536 7590
rect 66580 7098 66636 7100
rect 66660 7098 66716 7100
rect 66740 7098 66796 7100
rect 66820 7098 66876 7100
rect 66580 7046 66626 7098
rect 66626 7046 66636 7098
rect 66660 7046 66690 7098
rect 66690 7046 66702 7098
rect 66702 7046 66716 7098
rect 66740 7046 66754 7098
rect 66754 7046 66766 7098
rect 66766 7046 66796 7098
rect 66820 7046 66830 7098
rect 66830 7046 66876 7098
rect 66580 7044 66636 7046
rect 66660 7044 66716 7046
rect 66740 7044 66796 7046
rect 66820 7044 66876 7046
rect 67240 6554 67296 6556
rect 67320 6554 67376 6556
rect 67400 6554 67456 6556
rect 67480 6554 67536 6556
rect 67240 6502 67286 6554
rect 67286 6502 67296 6554
rect 67320 6502 67350 6554
rect 67350 6502 67362 6554
rect 67362 6502 67376 6554
rect 67400 6502 67414 6554
rect 67414 6502 67426 6554
rect 67426 6502 67456 6554
rect 67480 6502 67490 6554
rect 67490 6502 67536 6554
rect 67240 6500 67296 6502
rect 67320 6500 67376 6502
rect 67400 6500 67456 6502
rect 67480 6500 67536 6502
rect 48318 3848 48374 3904
rect 66580 6010 66636 6012
rect 66660 6010 66716 6012
rect 66740 6010 66796 6012
rect 66820 6010 66876 6012
rect 66580 5958 66626 6010
rect 66626 5958 66636 6010
rect 66660 5958 66690 6010
rect 66690 5958 66702 6010
rect 66702 5958 66716 6010
rect 66740 5958 66754 6010
rect 66754 5958 66766 6010
rect 66766 5958 66796 6010
rect 66820 5958 66830 6010
rect 66830 5958 66876 6010
rect 66580 5956 66636 5958
rect 66660 5956 66716 5958
rect 66740 5956 66796 5958
rect 66820 5956 66876 5958
rect 67240 5466 67296 5468
rect 67320 5466 67376 5468
rect 67400 5466 67456 5468
rect 67480 5466 67536 5468
rect 67240 5414 67286 5466
rect 67286 5414 67296 5466
rect 67320 5414 67350 5466
rect 67350 5414 67362 5466
rect 67362 5414 67376 5466
rect 67400 5414 67414 5466
rect 67414 5414 67426 5466
rect 67426 5414 67456 5466
rect 67480 5414 67490 5466
rect 67490 5414 67536 5466
rect 67240 5412 67296 5414
rect 67320 5412 67376 5414
rect 67400 5412 67456 5414
rect 67480 5412 67536 5414
rect 66580 4922 66636 4924
rect 66660 4922 66716 4924
rect 66740 4922 66796 4924
rect 66820 4922 66876 4924
rect 66580 4870 66626 4922
rect 66626 4870 66636 4922
rect 66660 4870 66690 4922
rect 66690 4870 66702 4922
rect 66702 4870 66716 4922
rect 66740 4870 66754 4922
rect 66754 4870 66766 4922
rect 66766 4870 66796 4922
rect 66820 4870 66830 4922
rect 66830 4870 66876 4922
rect 66580 4868 66636 4870
rect 66660 4868 66716 4870
rect 66740 4868 66796 4870
rect 66820 4868 66876 4870
rect 67240 4378 67296 4380
rect 67320 4378 67376 4380
rect 67400 4378 67456 4380
rect 67480 4378 67536 4380
rect 67240 4326 67286 4378
rect 67286 4326 67296 4378
rect 67320 4326 67350 4378
rect 67350 4326 67362 4378
rect 67362 4326 67376 4378
rect 67400 4326 67414 4378
rect 67414 4326 67426 4378
rect 67426 4326 67456 4378
rect 67480 4326 67490 4378
rect 67490 4326 67536 4378
rect 67240 4324 67296 4326
rect 67320 4324 67376 4326
rect 67400 4324 67456 4326
rect 67480 4324 67536 4326
rect 66580 3834 66636 3836
rect 66660 3834 66716 3836
rect 66740 3834 66796 3836
rect 66820 3834 66876 3836
rect 66580 3782 66626 3834
rect 66626 3782 66636 3834
rect 66660 3782 66690 3834
rect 66690 3782 66702 3834
rect 66702 3782 66716 3834
rect 66740 3782 66754 3834
rect 66754 3782 66766 3834
rect 66766 3782 66796 3834
rect 66820 3782 66830 3834
rect 66830 3782 66876 3834
rect 66580 3780 66636 3782
rect 66660 3780 66716 3782
rect 66740 3780 66796 3782
rect 66820 3780 66876 3782
rect 67240 3290 67296 3292
rect 67320 3290 67376 3292
rect 67400 3290 67456 3292
rect 67480 3290 67536 3292
rect 67240 3238 67286 3290
rect 67286 3238 67296 3290
rect 67320 3238 67350 3290
rect 67350 3238 67362 3290
rect 67362 3238 67376 3290
rect 67400 3238 67414 3290
rect 67414 3238 67426 3290
rect 67426 3238 67456 3290
rect 67480 3238 67490 3290
rect 67490 3238 67536 3290
rect 67240 3236 67296 3238
rect 67320 3236 67376 3238
rect 67400 3236 67456 3238
rect 67480 3236 67536 3238
rect 66580 2746 66636 2748
rect 66660 2746 66716 2748
rect 66740 2746 66796 2748
rect 66820 2746 66876 2748
rect 66580 2694 66626 2746
rect 66626 2694 66636 2746
rect 66660 2694 66690 2746
rect 66690 2694 66702 2746
rect 66702 2694 66716 2746
rect 66740 2694 66754 2746
rect 66754 2694 66766 2746
rect 66766 2694 66796 2746
rect 66820 2694 66830 2746
rect 66830 2694 66876 2746
rect 66580 2692 66636 2694
rect 66660 2692 66716 2694
rect 66740 2692 66796 2694
rect 66820 2692 66876 2694
rect 67240 2202 67296 2204
rect 67320 2202 67376 2204
rect 67400 2202 67456 2204
rect 67480 2202 67536 2204
rect 67240 2150 67286 2202
rect 67286 2150 67296 2202
rect 67320 2150 67350 2202
rect 67350 2150 67362 2202
rect 67362 2150 67376 2202
rect 67400 2150 67414 2202
rect 67414 2150 67426 2202
rect 67426 2150 67456 2202
rect 67480 2150 67490 2202
rect 67490 2150 67536 2202
rect 67240 2148 67296 2150
rect 67320 2148 67376 2150
rect 67400 2148 67456 2150
rect 67480 2148 67536 2150
rect 74262 1808 74318 1864
<< metal3 >>
rect 5130 37568 5446 37569
rect 5130 37504 5136 37568
rect 5200 37504 5216 37568
rect 5280 37504 5296 37568
rect 5360 37504 5376 37568
rect 5440 37504 5446 37568
rect 5130 37503 5446 37504
rect 35850 37568 36166 37569
rect 35850 37504 35856 37568
rect 35920 37504 35936 37568
rect 36000 37504 36016 37568
rect 36080 37504 36096 37568
rect 36160 37504 36166 37568
rect 35850 37503 36166 37504
rect 66570 37568 66886 37569
rect 66570 37504 66576 37568
rect 66640 37504 66656 37568
rect 66720 37504 66736 37568
rect 66800 37504 66816 37568
rect 66880 37504 66886 37568
rect 66570 37503 66886 37504
rect 5790 37024 6106 37025
rect 5790 36960 5796 37024
rect 5860 36960 5876 37024
rect 5940 36960 5956 37024
rect 6020 36960 6036 37024
rect 6100 36960 6106 37024
rect 5790 36959 6106 36960
rect 36510 37024 36826 37025
rect 36510 36960 36516 37024
rect 36580 36960 36596 37024
rect 36660 36960 36676 37024
rect 36740 36960 36756 37024
rect 36820 36960 36826 37024
rect 36510 36959 36826 36960
rect 67230 37024 67546 37025
rect 67230 36960 67236 37024
rect 67300 36960 67316 37024
rect 67380 36960 67396 37024
rect 67460 36960 67476 37024
rect 67540 36960 67546 37024
rect 67230 36959 67546 36960
rect 14549 36548 14615 36549
rect 14549 36544 14596 36548
rect 14660 36546 14666 36548
rect 14549 36488 14554 36544
rect 14549 36484 14596 36488
rect 14660 36486 14706 36546
rect 14660 36484 14666 36486
rect 14549 36483 14615 36484
rect 5130 36480 5446 36481
rect 5130 36416 5136 36480
rect 5200 36416 5216 36480
rect 5280 36416 5296 36480
rect 5360 36416 5376 36480
rect 5440 36416 5446 36480
rect 5130 36415 5446 36416
rect 35850 36480 36166 36481
rect 35850 36416 35856 36480
rect 35920 36416 35936 36480
rect 36000 36416 36016 36480
rect 36080 36416 36096 36480
rect 36160 36416 36166 36480
rect 35850 36415 36166 36416
rect 66570 36480 66886 36481
rect 66570 36416 66576 36480
rect 66640 36416 66656 36480
rect 66720 36416 66736 36480
rect 66800 36416 66816 36480
rect 66880 36416 66886 36480
rect 66570 36415 66886 36416
rect 31518 36348 31524 36412
rect 31588 36410 31594 36412
rect 32673 36410 32739 36413
rect 31588 36408 32739 36410
rect 31588 36352 32678 36408
rect 32734 36352 32739 36408
rect 31588 36350 32739 36352
rect 31588 36348 31594 36350
rect 32673 36347 32739 36350
rect 5790 35936 6106 35937
rect 5790 35872 5796 35936
rect 5860 35872 5876 35936
rect 5940 35872 5956 35936
rect 6020 35872 6036 35936
rect 6100 35872 6106 35936
rect 5790 35871 6106 35872
rect 36510 35936 36826 35937
rect 36510 35872 36516 35936
rect 36580 35872 36596 35936
rect 36660 35872 36676 35936
rect 36740 35872 36756 35936
rect 36820 35872 36826 35936
rect 36510 35871 36826 35872
rect 67230 35936 67546 35937
rect 67230 35872 67236 35936
rect 67300 35872 67316 35936
rect 67380 35872 67396 35936
rect 67460 35872 67476 35936
rect 67540 35872 67546 35936
rect 67230 35871 67546 35872
rect 5130 35392 5446 35393
rect 5130 35328 5136 35392
rect 5200 35328 5216 35392
rect 5280 35328 5296 35392
rect 5360 35328 5376 35392
rect 5440 35328 5446 35392
rect 5130 35327 5446 35328
rect 35850 35392 36166 35393
rect 35850 35328 35856 35392
rect 35920 35328 35936 35392
rect 36000 35328 36016 35392
rect 36080 35328 36096 35392
rect 36160 35328 36166 35392
rect 35850 35327 36166 35328
rect 66570 35392 66886 35393
rect 66570 35328 66576 35392
rect 66640 35328 66656 35392
rect 66720 35328 66736 35392
rect 66800 35328 66816 35392
rect 66880 35328 66886 35392
rect 66570 35327 66886 35328
rect 5790 34848 6106 34849
rect 5790 34784 5796 34848
rect 5860 34784 5876 34848
rect 5940 34784 5956 34848
rect 6020 34784 6036 34848
rect 6100 34784 6106 34848
rect 5790 34783 6106 34784
rect 36510 34848 36826 34849
rect 36510 34784 36516 34848
rect 36580 34784 36596 34848
rect 36660 34784 36676 34848
rect 36740 34784 36756 34848
rect 36820 34784 36826 34848
rect 36510 34783 36826 34784
rect 67230 34848 67546 34849
rect 67230 34784 67236 34848
rect 67300 34784 67316 34848
rect 67380 34784 67396 34848
rect 67460 34784 67476 34848
rect 67540 34784 67546 34848
rect 67230 34783 67546 34784
rect 5130 34304 5446 34305
rect 5130 34240 5136 34304
rect 5200 34240 5216 34304
rect 5280 34240 5296 34304
rect 5360 34240 5376 34304
rect 5440 34240 5446 34304
rect 5130 34239 5446 34240
rect 35850 34304 36166 34305
rect 35850 34240 35856 34304
rect 35920 34240 35936 34304
rect 36000 34240 36016 34304
rect 36080 34240 36096 34304
rect 36160 34240 36166 34304
rect 35850 34239 36166 34240
rect 66570 34304 66886 34305
rect 66570 34240 66576 34304
rect 66640 34240 66656 34304
rect 66720 34240 66736 34304
rect 66800 34240 66816 34304
rect 66880 34240 66886 34304
rect 66570 34239 66886 34240
rect 5790 33760 6106 33761
rect 5790 33696 5796 33760
rect 5860 33696 5876 33760
rect 5940 33696 5956 33760
rect 6020 33696 6036 33760
rect 6100 33696 6106 33760
rect 5790 33695 6106 33696
rect 36510 33760 36826 33761
rect 36510 33696 36516 33760
rect 36580 33696 36596 33760
rect 36660 33696 36676 33760
rect 36740 33696 36756 33760
rect 36820 33696 36826 33760
rect 36510 33695 36826 33696
rect 67230 33760 67546 33761
rect 67230 33696 67236 33760
rect 67300 33696 67316 33760
rect 67380 33696 67396 33760
rect 67460 33696 67476 33760
rect 67540 33696 67546 33760
rect 67230 33695 67546 33696
rect 5130 33216 5446 33217
rect 5130 33152 5136 33216
rect 5200 33152 5216 33216
rect 5280 33152 5296 33216
rect 5360 33152 5376 33216
rect 5440 33152 5446 33216
rect 5130 33151 5446 33152
rect 35850 33216 36166 33217
rect 35850 33152 35856 33216
rect 35920 33152 35936 33216
rect 36000 33152 36016 33216
rect 36080 33152 36096 33216
rect 36160 33152 36166 33216
rect 35850 33151 36166 33152
rect 66570 33216 66886 33217
rect 66570 33152 66576 33216
rect 66640 33152 66656 33216
rect 66720 33152 66736 33216
rect 66800 33152 66816 33216
rect 66880 33152 66886 33216
rect 66570 33151 66886 33152
rect 5790 32672 6106 32673
rect 5790 32608 5796 32672
rect 5860 32608 5876 32672
rect 5940 32608 5956 32672
rect 6020 32608 6036 32672
rect 6100 32608 6106 32672
rect 5790 32607 6106 32608
rect 36510 32672 36826 32673
rect 36510 32608 36516 32672
rect 36580 32608 36596 32672
rect 36660 32608 36676 32672
rect 36740 32608 36756 32672
rect 36820 32608 36826 32672
rect 36510 32607 36826 32608
rect 67230 32672 67546 32673
rect 67230 32608 67236 32672
rect 67300 32608 67316 32672
rect 67380 32608 67396 32672
rect 67460 32608 67476 32672
rect 67540 32608 67546 32672
rect 67230 32607 67546 32608
rect 7097 32466 7163 32469
rect 33174 32466 33180 32468
rect 7097 32464 33180 32466
rect 7097 32408 7102 32464
rect 7158 32408 33180 32464
rect 7097 32406 33180 32408
rect 7097 32403 7163 32406
rect 33174 32404 33180 32406
rect 33244 32404 33250 32468
rect 5130 32128 5446 32129
rect 5130 32064 5136 32128
rect 5200 32064 5216 32128
rect 5280 32064 5296 32128
rect 5360 32064 5376 32128
rect 5440 32064 5446 32128
rect 5130 32063 5446 32064
rect 35850 32128 36166 32129
rect 35850 32064 35856 32128
rect 35920 32064 35936 32128
rect 36000 32064 36016 32128
rect 36080 32064 36096 32128
rect 36160 32064 36166 32128
rect 35850 32063 36166 32064
rect 66570 32128 66886 32129
rect 66570 32064 66576 32128
rect 66640 32064 66656 32128
rect 66720 32064 66736 32128
rect 66800 32064 66816 32128
rect 66880 32064 66886 32128
rect 66570 32063 66886 32064
rect 5790 31584 6106 31585
rect 5790 31520 5796 31584
rect 5860 31520 5876 31584
rect 5940 31520 5956 31584
rect 6020 31520 6036 31584
rect 6100 31520 6106 31584
rect 5790 31519 6106 31520
rect 36510 31584 36826 31585
rect 36510 31520 36516 31584
rect 36580 31520 36596 31584
rect 36660 31520 36676 31584
rect 36740 31520 36756 31584
rect 36820 31520 36826 31584
rect 36510 31519 36826 31520
rect 67230 31584 67546 31585
rect 67230 31520 67236 31584
rect 67300 31520 67316 31584
rect 67380 31520 67396 31584
rect 67460 31520 67476 31584
rect 67540 31520 67546 31584
rect 67230 31519 67546 31520
rect 5130 31040 5446 31041
rect 5130 30976 5136 31040
rect 5200 30976 5216 31040
rect 5280 30976 5296 31040
rect 5360 30976 5376 31040
rect 5440 30976 5446 31040
rect 5130 30975 5446 30976
rect 35850 31040 36166 31041
rect 35850 30976 35856 31040
rect 35920 30976 35936 31040
rect 36000 30976 36016 31040
rect 36080 30976 36096 31040
rect 36160 30976 36166 31040
rect 35850 30975 36166 30976
rect 66570 31040 66886 31041
rect 66570 30976 66576 31040
rect 66640 30976 66656 31040
rect 66720 30976 66736 31040
rect 66800 30976 66816 31040
rect 66880 30976 66886 31040
rect 66570 30975 66886 30976
rect 5790 30496 6106 30497
rect 5790 30432 5796 30496
rect 5860 30432 5876 30496
rect 5940 30432 5956 30496
rect 6020 30432 6036 30496
rect 6100 30432 6106 30496
rect 5790 30431 6106 30432
rect 36510 30496 36826 30497
rect 36510 30432 36516 30496
rect 36580 30432 36596 30496
rect 36660 30432 36676 30496
rect 36740 30432 36756 30496
rect 36820 30432 36826 30496
rect 36510 30431 36826 30432
rect 67230 30496 67546 30497
rect 67230 30432 67236 30496
rect 67300 30432 67316 30496
rect 67380 30432 67396 30496
rect 67460 30432 67476 30496
rect 67540 30432 67546 30496
rect 67230 30431 67546 30432
rect 5130 29952 5446 29953
rect 5130 29888 5136 29952
rect 5200 29888 5216 29952
rect 5280 29888 5296 29952
rect 5360 29888 5376 29952
rect 5440 29888 5446 29952
rect 5130 29887 5446 29888
rect 35850 29952 36166 29953
rect 35850 29888 35856 29952
rect 35920 29888 35936 29952
rect 36000 29888 36016 29952
rect 36080 29888 36096 29952
rect 36160 29888 36166 29952
rect 35850 29887 36166 29888
rect 66570 29952 66886 29953
rect 66570 29888 66576 29952
rect 66640 29888 66656 29952
rect 66720 29888 66736 29952
rect 66800 29888 66816 29952
rect 66880 29888 66886 29952
rect 66570 29887 66886 29888
rect 10961 29610 11027 29613
rect 26734 29610 26740 29612
rect 10961 29608 26740 29610
rect 10961 29552 10966 29608
rect 11022 29552 26740 29608
rect 10961 29550 26740 29552
rect 10961 29547 11027 29550
rect 26734 29548 26740 29550
rect 26804 29548 26810 29612
rect 5790 29408 6106 29409
rect 5790 29344 5796 29408
rect 5860 29344 5876 29408
rect 5940 29344 5956 29408
rect 6020 29344 6036 29408
rect 6100 29344 6106 29408
rect 5790 29343 6106 29344
rect 36510 29408 36826 29409
rect 36510 29344 36516 29408
rect 36580 29344 36596 29408
rect 36660 29344 36676 29408
rect 36740 29344 36756 29408
rect 36820 29344 36826 29408
rect 36510 29343 36826 29344
rect 67230 29408 67546 29409
rect 67230 29344 67236 29408
rect 67300 29344 67316 29408
rect 67380 29344 67396 29408
rect 67460 29344 67476 29408
rect 67540 29344 67546 29408
rect 67230 29343 67546 29344
rect 5130 28864 5446 28865
rect 5130 28800 5136 28864
rect 5200 28800 5216 28864
rect 5280 28800 5296 28864
rect 5360 28800 5376 28864
rect 5440 28800 5446 28864
rect 5130 28799 5446 28800
rect 35850 28864 36166 28865
rect 35850 28800 35856 28864
rect 35920 28800 35936 28864
rect 36000 28800 36016 28864
rect 36080 28800 36096 28864
rect 36160 28800 36166 28864
rect 35850 28799 36166 28800
rect 66570 28864 66886 28865
rect 66570 28800 66576 28864
rect 66640 28800 66656 28864
rect 66720 28800 66736 28864
rect 66800 28800 66816 28864
rect 66880 28800 66886 28864
rect 66570 28799 66886 28800
rect 5790 28320 6106 28321
rect 5790 28256 5796 28320
rect 5860 28256 5876 28320
rect 5940 28256 5956 28320
rect 6020 28256 6036 28320
rect 6100 28256 6106 28320
rect 5790 28255 6106 28256
rect 36510 28320 36826 28321
rect 36510 28256 36516 28320
rect 36580 28256 36596 28320
rect 36660 28256 36676 28320
rect 36740 28256 36756 28320
rect 36820 28256 36826 28320
rect 36510 28255 36826 28256
rect 67230 28320 67546 28321
rect 67230 28256 67236 28320
rect 67300 28256 67316 28320
rect 67380 28256 67396 28320
rect 67460 28256 67476 28320
rect 67540 28256 67546 28320
rect 67230 28255 67546 28256
rect 5130 27776 5446 27777
rect 5130 27712 5136 27776
rect 5200 27712 5216 27776
rect 5280 27712 5296 27776
rect 5360 27712 5376 27776
rect 5440 27712 5446 27776
rect 5130 27711 5446 27712
rect 35850 27776 36166 27777
rect 35850 27712 35856 27776
rect 35920 27712 35936 27776
rect 36000 27712 36016 27776
rect 36080 27712 36096 27776
rect 36160 27712 36166 27776
rect 35850 27711 36166 27712
rect 66570 27776 66886 27777
rect 66570 27712 66576 27776
rect 66640 27712 66656 27776
rect 66720 27712 66736 27776
rect 66800 27712 66816 27776
rect 66880 27712 66886 27776
rect 66570 27711 66886 27712
rect 5790 27232 6106 27233
rect 5790 27168 5796 27232
rect 5860 27168 5876 27232
rect 5940 27168 5956 27232
rect 6020 27168 6036 27232
rect 6100 27168 6106 27232
rect 5790 27167 6106 27168
rect 36510 27232 36826 27233
rect 36510 27168 36516 27232
rect 36580 27168 36596 27232
rect 36660 27168 36676 27232
rect 36740 27168 36756 27232
rect 36820 27168 36826 27232
rect 36510 27167 36826 27168
rect 67230 27232 67546 27233
rect 67230 27168 67236 27232
rect 67300 27168 67316 27232
rect 67380 27168 67396 27232
rect 67460 27168 67476 27232
rect 67540 27168 67546 27232
rect 67230 27167 67546 27168
rect 5130 26688 5446 26689
rect 5130 26624 5136 26688
rect 5200 26624 5216 26688
rect 5280 26624 5296 26688
rect 5360 26624 5376 26688
rect 5440 26624 5446 26688
rect 5130 26623 5446 26624
rect 35850 26688 36166 26689
rect 35850 26624 35856 26688
rect 35920 26624 35936 26688
rect 36000 26624 36016 26688
rect 36080 26624 36096 26688
rect 36160 26624 36166 26688
rect 35850 26623 36166 26624
rect 66570 26688 66886 26689
rect 66570 26624 66576 26688
rect 66640 26624 66656 26688
rect 66720 26624 66736 26688
rect 66800 26624 66816 26688
rect 66880 26624 66886 26688
rect 66570 26623 66886 26624
rect 5790 26144 6106 26145
rect 5790 26080 5796 26144
rect 5860 26080 5876 26144
rect 5940 26080 5956 26144
rect 6020 26080 6036 26144
rect 6100 26080 6106 26144
rect 5790 26079 6106 26080
rect 36510 26144 36826 26145
rect 36510 26080 36516 26144
rect 36580 26080 36596 26144
rect 36660 26080 36676 26144
rect 36740 26080 36756 26144
rect 36820 26080 36826 26144
rect 36510 26079 36826 26080
rect 67230 26144 67546 26145
rect 67230 26080 67236 26144
rect 67300 26080 67316 26144
rect 67380 26080 67396 26144
rect 67460 26080 67476 26144
rect 67540 26080 67546 26144
rect 67230 26079 67546 26080
rect 5130 25600 5446 25601
rect 5130 25536 5136 25600
rect 5200 25536 5216 25600
rect 5280 25536 5296 25600
rect 5360 25536 5376 25600
rect 5440 25536 5446 25600
rect 5130 25535 5446 25536
rect 35850 25600 36166 25601
rect 35850 25536 35856 25600
rect 35920 25536 35936 25600
rect 36000 25536 36016 25600
rect 36080 25536 36096 25600
rect 36160 25536 36166 25600
rect 35850 25535 36166 25536
rect 66570 25600 66886 25601
rect 66570 25536 66576 25600
rect 66640 25536 66656 25600
rect 66720 25536 66736 25600
rect 66800 25536 66816 25600
rect 66880 25536 66886 25600
rect 66570 25535 66886 25536
rect 5790 25056 6106 25057
rect 5790 24992 5796 25056
rect 5860 24992 5876 25056
rect 5940 24992 5956 25056
rect 6020 24992 6036 25056
rect 6100 24992 6106 25056
rect 5790 24991 6106 24992
rect 36510 25056 36826 25057
rect 36510 24992 36516 25056
rect 36580 24992 36596 25056
rect 36660 24992 36676 25056
rect 36740 24992 36756 25056
rect 36820 24992 36826 25056
rect 36510 24991 36826 24992
rect 67230 25056 67546 25057
rect 67230 24992 67236 25056
rect 67300 24992 67316 25056
rect 67380 24992 67396 25056
rect 67460 24992 67476 25056
rect 67540 24992 67546 25056
rect 67230 24991 67546 24992
rect 5130 24512 5446 24513
rect 5130 24448 5136 24512
rect 5200 24448 5216 24512
rect 5280 24448 5296 24512
rect 5360 24448 5376 24512
rect 5440 24448 5446 24512
rect 5130 24447 5446 24448
rect 35850 24512 36166 24513
rect 35850 24448 35856 24512
rect 35920 24448 35936 24512
rect 36000 24448 36016 24512
rect 36080 24448 36096 24512
rect 36160 24448 36166 24512
rect 35850 24447 36166 24448
rect 66570 24512 66886 24513
rect 66570 24448 66576 24512
rect 66640 24448 66656 24512
rect 66720 24448 66736 24512
rect 66800 24448 66816 24512
rect 66880 24448 66886 24512
rect 66570 24447 66886 24448
rect 5790 23968 6106 23969
rect 5790 23904 5796 23968
rect 5860 23904 5876 23968
rect 5940 23904 5956 23968
rect 6020 23904 6036 23968
rect 6100 23904 6106 23968
rect 5790 23903 6106 23904
rect 36510 23968 36826 23969
rect 36510 23904 36516 23968
rect 36580 23904 36596 23968
rect 36660 23904 36676 23968
rect 36740 23904 36756 23968
rect 36820 23904 36826 23968
rect 36510 23903 36826 23904
rect 67230 23968 67546 23969
rect 67230 23904 67236 23968
rect 67300 23904 67316 23968
rect 67380 23904 67396 23968
rect 67460 23904 67476 23968
rect 67540 23904 67546 23968
rect 67230 23903 67546 23904
rect 5130 23424 5446 23425
rect 5130 23360 5136 23424
rect 5200 23360 5216 23424
rect 5280 23360 5296 23424
rect 5360 23360 5376 23424
rect 5440 23360 5446 23424
rect 5130 23359 5446 23360
rect 35850 23424 36166 23425
rect 35850 23360 35856 23424
rect 35920 23360 35936 23424
rect 36000 23360 36016 23424
rect 36080 23360 36096 23424
rect 36160 23360 36166 23424
rect 35850 23359 36166 23360
rect 66570 23424 66886 23425
rect 66570 23360 66576 23424
rect 66640 23360 66656 23424
rect 66720 23360 66736 23424
rect 66800 23360 66816 23424
rect 66880 23360 66886 23424
rect 66570 23359 66886 23360
rect 5790 22880 6106 22881
rect 5790 22816 5796 22880
rect 5860 22816 5876 22880
rect 5940 22816 5956 22880
rect 6020 22816 6036 22880
rect 6100 22816 6106 22880
rect 5790 22815 6106 22816
rect 36510 22880 36826 22881
rect 36510 22816 36516 22880
rect 36580 22816 36596 22880
rect 36660 22816 36676 22880
rect 36740 22816 36756 22880
rect 36820 22816 36826 22880
rect 36510 22815 36826 22816
rect 67230 22880 67546 22881
rect 67230 22816 67236 22880
rect 67300 22816 67316 22880
rect 67380 22816 67396 22880
rect 67460 22816 67476 22880
rect 67540 22816 67546 22880
rect 67230 22815 67546 22816
rect 5130 22336 5446 22337
rect 5130 22272 5136 22336
rect 5200 22272 5216 22336
rect 5280 22272 5296 22336
rect 5360 22272 5376 22336
rect 5440 22272 5446 22336
rect 5130 22271 5446 22272
rect 35850 22336 36166 22337
rect 35850 22272 35856 22336
rect 35920 22272 35936 22336
rect 36000 22272 36016 22336
rect 36080 22272 36096 22336
rect 36160 22272 36166 22336
rect 35850 22271 36166 22272
rect 66570 22336 66886 22337
rect 66570 22272 66576 22336
rect 66640 22272 66656 22336
rect 66720 22272 66736 22336
rect 66800 22272 66816 22336
rect 66880 22272 66886 22336
rect 66570 22271 66886 22272
rect 5790 21792 6106 21793
rect 5790 21728 5796 21792
rect 5860 21728 5876 21792
rect 5940 21728 5956 21792
rect 6020 21728 6036 21792
rect 6100 21728 6106 21792
rect 5790 21727 6106 21728
rect 36510 21792 36826 21793
rect 36510 21728 36516 21792
rect 36580 21728 36596 21792
rect 36660 21728 36676 21792
rect 36740 21728 36756 21792
rect 36820 21728 36826 21792
rect 36510 21727 36826 21728
rect 67230 21792 67546 21793
rect 67230 21728 67236 21792
rect 67300 21728 67316 21792
rect 67380 21728 67396 21792
rect 67460 21728 67476 21792
rect 67540 21728 67546 21792
rect 67230 21727 67546 21728
rect 5130 21248 5446 21249
rect 5130 21184 5136 21248
rect 5200 21184 5216 21248
rect 5280 21184 5296 21248
rect 5360 21184 5376 21248
rect 5440 21184 5446 21248
rect 5130 21183 5446 21184
rect 35850 21248 36166 21249
rect 35850 21184 35856 21248
rect 35920 21184 35936 21248
rect 36000 21184 36016 21248
rect 36080 21184 36096 21248
rect 36160 21184 36166 21248
rect 35850 21183 36166 21184
rect 66570 21248 66886 21249
rect 66570 21184 66576 21248
rect 66640 21184 66656 21248
rect 66720 21184 66736 21248
rect 66800 21184 66816 21248
rect 66880 21184 66886 21248
rect 66570 21183 66886 21184
rect 5790 20704 6106 20705
rect 5790 20640 5796 20704
rect 5860 20640 5876 20704
rect 5940 20640 5956 20704
rect 6020 20640 6036 20704
rect 6100 20640 6106 20704
rect 5790 20639 6106 20640
rect 36510 20704 36826 20705
rect 36510 20640 36516 20704
rect 36580 20640 36596 20704
rect 36660 20640 36676 20704
rect 36740 20640 36756 20704
rect 36820 20640 36826 20704
rect 36510 20639 36826 20640
rect 67230 20704 67546 20705
rect 67230 20640 67236 20704
rect 67300 20640 67316 20704
rect 67380 20640 67396 20704
rect 67460 20640 67476 20704
rect 67540 20640 67546 20704
rect 67230 20639 67546 20640
rect 5130 20160 5446 20161
rect 5130 20096 5136 20160
rect 5200 20096 5216 20160
rect 5280 20096 5296 20160
rect 5360 20096 5376 20160
rect 5440 20096 5446 20160
rect 5130 20095 5446 20096
rect 35850 20160 36166 20161
rect 35850 20096 35856 20160
rect 35920 20096 35936 20160
rect 36000 20096 36016 20160
rect 36080 20096 36096 20160
rect 36160 20096 36166 20160
rect 35850 20095 36166 20096
rect 66570 20160 66886 20161
rect 66570 20096 66576 20160
rect 66640 20096 66656 20160
rect 66720 20096 66736 20160
rect 66800 20096 66816 20160
rect 66880 20096 66886 20160
rect 66570 20095 66886 20096
rect 5790 19616 6106 19617
rect 5790 19552 5796 19616
rect 5860 19552 5876 19616
rect 5940 19552 5956 19616
rect 6020 19552 6036 19616
rect 6100 19552 6106 19616
rect 5790 19551 6106 19552
rect 36510 19616 36826 19617
rect 36510 19552 36516 19616
rect 36580 19552 36596 19616
rect 36660 19552 36676 19616
rect 36740 19552 36756 19616
rect 36820 19552 36826 19616
rect 36510 19551 36826 19552
rect 67230 19616 67546 19617
rect 67230 19552 67236 19616
rect 67300 19552 67316 19616
rect 67380 19552 67396 19616
rect 67460 19552 67476 19616
rect 67540 19552 67546 19616
rect 67230 19551 67546 19552
rect 5130 19072 5446 19073
rect 5130 19008 5136 19072
rect 5200 19008 5216 19072
rect 5280 19008 5296 19072
rect 5360 19008 5376 19072
rect 5440 19008 5446 19072
rect 5130 19007 5446 19008
rect 35850 19072 36166 19073
rect 35850 19008 35856 19072
rect 35920 19008 35936 19072
rect 36000 19008 36016 19072
rect 36080 19008 36096 19072
rect 36160 19008 36166 19072
rect 35850 19007 36166 19008
rect 66570 19072 66886 19073
rect 66570 19008 66576 19072
rect 66640 19008 66656 19072
rect 66720 19008 66736 19072
rect 66800 19008 66816 19072
rect 66880 19008 66886 19072
rect 66570 19007 66886 19008
rect 5790 18528 6106 18529
rect 5790 18464 5796 18528
rect 5860 18464 5876 18528
rect 5940 18464 5956 18528
rect 6020 18464 6036 18528
rect 6100 18464 6106 18528
rect 5790 18463 6106 18464
rect 36510 18528 36826 18529
rect 36510 18464 36516 18528
rect 36580 18464 36596 18528
rect 36660 18464 36676 18528
rect 36740 18464 36756 18528
rect 36820 18464 36826 18528
rect 36510 18463 36826 18464
rect 67230 18528 67546 18529
rect 67230 18464 67236 18528
rect 67300 18464 67316 18528
rect 67380 18464 67396 18528
rect 67460 18464 67476 18528
rect 67540 18464 67546 18528
rect 67230 18463 67546 18464
rect 5130 17984 5446 17985
rect 5130 17920 5136 17984
rect 5200 17920 5216 17984
rect 5280 17920 5296 17984
rect 5360 17920 5376 17984
rect 5440 17920 5446 17984
rect 5130 17919 5446 17920
rect 35850 17984 36166 17985
rect 35850 17920 35856 17984
rect 35920 17920 35936 17984
rect 36000 17920 36016 17984
rect 36080 17920 36096 17984
rect 36160 17920 36166 17984
rect 35850 17919 36166 17920
rect 66570 17984 66886 17985
rect 66570 17920 66576 17984
rect 66640 17920 66656 17984
rect 66720 17920 66736 17984
rect 66800 17920 66816 17984
rect 66880 17920 66886 17984
rect 66570 17919 66886 17920
rect 5790 17440 6106 17441
rect 5790 17376 5796 17440
rect 5860 17376 5876 17440
rect 5940 17376 5956 17440
rect 6020 17376 6036 17440
rect 6100 17376 6106 17440
rect 5790 17375 6106 17376
rect 36510 17440 36826 17441
rect 36510 17376 36516 17440
rect 36580 17376 36596 17440
rect 36660 17376 36676 17440
rect 36740 17376 36756 17440
rect 36820 17376 36826 17440
rect 36510 17375 36826 17376
rect 67230 17440 67546 17441
rect 67230 17376 67236 17440
rect 67300 17376 67316 17440
rect 67380 17376 67396 17440
rect 67460 17376 67476 17440
rect 67540 17376 67546 17440
rect 67230 17375 67546 17376
rect 5130 16896 5446 16897
rect 5130 16832 5136 16896
rect 5200 16832 5216 16896
rect 5280 16832 5296 16896
rect 5360 16832 5376 16896
rect 5440 16832 5446 16896
rect 5130 16831 5446 16832
rect 35850 16896 36166 16897
rect 35850 16832 35856 16896
rect 35920 16832 35936 16896
rect 36000 16832 36016 16896
rect 36080 16832 36096 16896
rect 36160 16832 36166 16896
rect 35850 16831 36166 16832
rect 66570 16896 66886 16897
rect 66570 16832 66576 16896
rect 66640 16832 66656 16896
rect 66720 16832 66736 16896
rect 66800 16832 66816 16896
rect 66880 16832 66886 16896
rect 66570 16831 66886 16832
rect 5790 16352 6106 16353
rect 5790 16288 5796 16352
rect 5860 16288 5876 16352
rect 5940 16288 5956 16352
rect 6020 16288 6036 16352
rect 6100 16288 6106 16352
rect 5790 16287 6106 16288
rect 36510 16352 36826 16353
rect 36510 16288 36516 16352
rect 36580 16288 36596 16352
rect 36660 16288 36676 16352
rect 36740 16288 36756 16352
rect 36820 16288 36826 16352
rect 36510 16287 36826 16288
rect 67230 16352 67546 16353
rect 67230 16288 67236 16352
rect 67300 16288 67316 16352
rect 67380 16288 67396 16352
rect 67460 16288 67476 16352
rect 67540 16288 67546 16352
rect 67230 16287 67546 16288
rect 5130 15808 5446 15809
rect 5130 15744 5136 15808
rect 5200 15744 5216 15808
rect 5280 15744 5296 15808
rect 5360 15744 5376 15808
rect 5440 15744 5446 15808
rect 5130 15743 5446 15744
rect 35850 15808 36166 15809
rect 35850 15744 35856 15808
rect 35920 15744 35936 15808
rect 36000 15744 36016 15808
rect 36080 15744 36096 15808
rect 36160 15744 36166 15808
rect 35850 15743 36166 15744
rect 66570 15808 66886 15809
rect 66570 15744 66576 15808
rect 66640 15744 66656 15808
rect 66720 15744 66736 15808
rect 66800 15744 66816 15808
rect 66880 15744 66886 15808
rect 66570 15743 66886 15744
rect 5790 15264 6106 15265
rect 5790 15200 5796 15264
rect 5860 15200 5876 15264
rect 5940 15200 5956 15264
rect 6020 15200 6036 15264
rect 6100 15200 6106 15264
rect 5790 15199 6106 15200
rect 36510 15264 36826 15265
rect 36510 15200 36516 15264
rect 36580 15200 36596 15264
rect 36660 15200 36676 15264
rect 36740 15200 36756 15264
rect 36820 15200 36826 15264
rect 36510 15199 36826 15200
rect 67230 15264 67546 15265
rect 67230 15200 67236 15264
rect 67300 15200 67316 15264
rect 67380 15200 67396 15264
rect 67460 15200 67476 15264
rect 67540 15200 67546 15264
rect 67230 15199 67546 15200
rect 5130 14720 5446 14721
rect 5130 14656 5136 14720
rect 5200 14656 5216 14720
rect 5280 14656 5296 14720
rect 5360 14656 5376 14720
rect 5440 14656 5446 14720
rect 5130 14655 5446 14656
rect 35850 14720 36166 14721
rect 35850 14656 35856 14720
rect 35920 14656 35936 14720
rect 36000 14656 36016 14720
rect 36080 14656 36096 14720
rect 36160 14656 36166 14720
rect 35850 14655 36166 14656
rect 66570 14720 66886 14721
rect 66570 14656 66576 14720
rect 66640 14656 66656 14720
rect 66720 14656 66736 14720
rect 66800 14656 66816 14720
rect 66880 14656 66886 14720
rect 66570 14655 66886 14656
rect 5790 14176 6106 14177
rect 5790 14112 5796 14176
rect 5860 14112 5876 14176
rect 5940 14112 5956 14176
rect 6020 14112 6036 14176
rect 6100 14112 6106 14176
rect 5790 14111 6106 14112
rect 36510 14176 36826 14177
rect 36510 14112 36516 14176
rect 36580 14112 36596 14176
rect 36660 14112 36676 14176
rect 36740 14112 36756 14176
rect 36820 14112 36826 14176
rect 36510 14111 36826 14112
rect 67230 14176 67546 14177
rect 67230 14112 67236 14176
rect 67300 14112 67316 14176
rect 67380 14112 67396 14176
rect 67460 14112 67476 14176
rect 67540 14112 67546 14176
rect 67230 14111 67546 14112
rect 5130 13632 5446 13633
rect 5130 13568 5136 13632
rect 5200 13568 5216 13632
rect 5280 13568 5296 13632
rect 5360 13568 5376 13632
rect 5440 13568 5446 13632
rect 5130 13567 5446 13568
rect 35850 13632 36166 13633
rect 35850 13568 35856 13632
rect 35920 13568 35936 13632
rect 36000 13568 36016 13632
rect 36080 13568 36096 13632
rect 36160 13568 36166 13632
rect 35850 13567 36166 13568
rect 66570 13632 66886 13633
rect 66570 13568 66576 13632
rect 66640 13568 66656 13632
rect 66720 13568 66736 13632
rect 66800 13568 66816 13632
rect 66880 13568 66886 13632
rect 66570 13567 66886 13568
rect 5790 13088 6106 13089
rect 5790 13024 5796 13088
rect 5860 13024 5876 13088
rect 5940 13024 5956 13088
rect 6020 13024 6036 13088
rect 6100 13024 6106 13088
rect 5790 13023 6106 13024
rect 36510 13088 36826 13089
rect 36510 13024 36516 13088
rect 36580 13024 36596 13088
rect 36660 13024 36676 13088
rect 36740 13024 36756 13088
rect 36820 13024 36826 13088
rect 36510 13023 36826 13024
rect 67230 13088 67546 13089
rect 67230 13024 67236 13088
rect 67300 13024 67316 13088
rect 67380 13024 67396 13088
rect 67460 13024 67476 13088
rect 67540 13024 67546 13088
rect 67230 13023 67546 13024
rect 5130 12544 5446 12545
rect 5130 12480 5136 12544
rect 5200 12480 5216 12544
rect 5280 12480 5296 12544
rect 5360 12480 5376 12544
rect 5440 12480 5446 12544
rect 5130 12479 5446 12480
rect 35850 12544 36166 12545
rect 35850 12480 35856 12544
rect 35920 12480 35936 12544
rect 36000 12480 36016 12544
rect 36080 12480 36096 12544
rect 36160 12480 36166 12544
rect 35850 12479 36166 12480
rect 66570 12544 66886 12545
rect 66570 12480 66576 12544
rect 66640 12480 66656 12544
rect 66720 12480 66736 12544
rect 66800 12480 66816 12544
rect 66880 12480 66886 12544
rect 66570 12479 66886 12480
rect 5790 12000 6106 12001
rect 5790 11936 5796 12000
rect 5860 11936 5876 12000
rect 5940 11936 5956 12000
rect 6020 11936 6036 12000
rect 6100 11936 6106 12000
rect 5790 11935 6106 11936
rect 36510 12000 36826 12001
rect 36510 11936 36516 12000
rect 36580 11936 36596 12000
rect 36660 11936 36676 12000
rect 36740 11936 36756 12000
rect 36820 11936 36826 12000
rect 36510 11935 36826 11936
rect 67230 12000 67546 12001
rect 67230 11936 67236 12000
rect 67300 11936 67316 12000
rect 67380 11936 67396 12000
rect 67460 11936 67476 12000
rect 67540 11936 67546 12000
rect 67230 11935 67546 11936
rect 20662 11868 20668 11932
rect 20732 11930 20738 11932
rect 28809 11930 28875 11933
rect 20732 11928 28875 11930
rect 20732 11872 28814 11928
rect 28870 11872 28875 11928
rect 20732 11870 28875 11872
rect 20732 11868 20738 11870
rect 28809 11867 28875 11870
rect 17534 11596 17540 11660
rect 17604 11658 17610 11660
rect 28441 11658 28507 11661
rect 17604 11656 28507 11658
rect 17604 11600 28446 11656
rect 28502 11600 28507 11656
rect 17604 11598 28507 11600
rect 17604 11596 17610 11598
rect 28441 11595 28507 11598
rect 15694 11460 15700 11524
rect 15764 11522 15770 11524
rect 25221 11522 25287 11525
rect 15764 11520 25287 11522
rect 15764 11464 25226 11520
rect 25282 11464 25287 11520
rect 15764 11462 25287 11464
rect 15764 11460 15770 11462
rect 25221 11459 25287 11462
rect 5130 11456 5446 11457
rect 5130 11392 5136 11456
rect 5200 11392 5216 11456
rect 5280 11392 5296 11456
rect 5360 11392 5376 11456
rect 5440 11392 5446 11456
rect 5130 11391 5446 11392
rect 35850 11456 36166 11457
rect 35850 11392 35856 11456
rect 35920 11392 35936 11456
rect 36000 11392 36016 11456
rect 36080 11392 36096 11456
rect 36160 11392 36166 11456
rect 35850 11391 36166 11392
rect 66570 11456 66886 11457
rect 66570 11392 66576 11456
rect 66640 11392 66656 11456
rect 66720 11392 66736 11456
rect 66800 11392 66816 11456
rect 66880 11392 66886 11456
rect 66570 11391 66886 11392
rect 11462 11324 11468 11388
rect 11532 11386 11538 11388
rect 21725 11386 21791 11389
rect 11532 11384 21791 11386
rect 11532 11328 21730 11384
rect 21786 11328 21791 11384
rect 11532 11326 21791 11328
rect 11532 11324 11538 11326
rect 21725 11323 21791 11326
rect 22461 11386 22527 11389
rect 26049 11386 26115 11389
rect 22461 11384 26115 11386
rect 22461 11328 22466 11384
rect 22522 11328 26054 11384
rect 26110 11328 26115 11384
rect 22461 11326 26115 11328
rect 22461 11323 22527 11326
rect 26049 11323 26115 11326
rect 11646 11188 11652 11252
rect 11716 11250 11722 11252
rect 22737 11250 22803 11253
rect 11716 11248 22803 11250
rect 11716 11192 22742 11248
rect 22798 11192 22803 11248
rect 11716 11190 22803 11192
rect 11716 11188 11722 11190
rect 22737 11187 22803 11190
rect 23197 11250 23263 11253
rect 26233 11252 26299 11253
rect 23422 11250 23428 11252
rect 23197 11248 23428 11250
rect 23197 11192 23202 11248
rect 23258 11192 23428 11248
rect 23197 11190 23428 11192
rect 23197 11187 23263 11190
rect 23422 11188 23428 11190
rect 23492 11188 23498 11252
rect 26182 11250 26188 11252
rect 26142 11190 26188 11250
rect 26252 11248 26299 11252
rect 26294 11192 26299 11248
rect 26182 11188 26188 11190
rect 26252 11188 26299 11192
rect 26233 11187 26299 11188
rect 12198 11052 12204 11116
rect 12268 11114 12274 11116
rect 23381 11114 23447 11117
rect 12268 11112 23447 11114
rect 12268 11056 23386 11112
rect 23442 11056 23447 11112
rect 12268 11054 23447 11056
rect 12268 11052 12274 11054
rect 23381 11051 23447 11054
rect 24526 11052 24532 11116
rect 24596 11114 24602 11116
rect 30465 11114 30531 11117
rect 24596 11112 30531 11114
rect 24596 11056 30470 11112
rect 30526 11056 30531 11112
rect 24596 11054 30531 11056
rect 24596 11052 24602 11054
rect 30465 11051 30531 11054
rect 15878 10916 15884 10980
rect 15948 10978 15954 10980
rect 33317 10978 33383 10981
rect 15948 10976 33383 10978
rect 15948 10920 33322 10976
rect 33378 10920 33383 10976
rect 15948 10918 33383 10920
rect 15948 10916 15954 10918
rect 33317 10915 33383 10918
rect 5790 10912 6106 10913
rect 5790 10848 5796 10912
rect 5860 10848 5876 10912
rect 5940 10848 5956 10912
rect 6020 10848 6036 10912
rect 6100 10848 6106 10912
rect 5790 10847 6106 10848
rect 36510 10912 36826 10913
rect 36510 10848 36516 10912
rect 36580 10848 36596 10912
rect 36660 10848 36676 10912
rect 36740 10848 36756 10912
rect 36820 10848 36826 10912
rect 36510 10847 36826 10848
rect 67230 10912 67546 10913
rect 67230 10848 67236 10912
rect 67300 10848 67316 10912
rect 67380 10848 67396 10912
rect 67460 10848 67476 10912
rect 67540 10848 67546 10912
rect 67230 10847 67546 10848
rect 21817 10842 21883 10845
rect 25313 10842 25379 10845
rect 21817 10840 25379 10842
rect 21817 10784 21822 10840
rect 21878 10784 25318 10840
rect 25374 10784 25379 10840
rect 21817 10782 25379 10784
rect 21817 10779 21883 10782
rect 25313 10779 25379 10782
rect 25814 10780 25820 10844
rect 25884 10842 25890 10844
rect 29545 10842 29611 10845
rect 25884 10840 29611 10842
rect 25884 10784 29550 10840
rect 29606 10784 29611 10840
rect 25884 10782 29611 10784
rect 25884 10780 25890 10782
rect 29545 10779 29611 10782
rect 11605 10706 11671 10709
rect 26049 10706 26115 10709
rect 11605 10704 26115 10706
rect 11605 10648 11610 10704
rect 11666 10648 26054 10704
rect 26110 10648 26115 10704
rect 11605 10646 26115 10648
rect 11605 10643 11671 10646
rect 26049 10643 26115 10646
rect 17953 10570 18019 10573
rect 28809 10570 28875 10573
rect 17953 10568 28875 10570
rect 17953 10512 17958 10568
rect 18014 10512 28814 10568
rect 28870 10512 28875 10568
rect 17953 10510 28875 10512
rect 17953 10507 18019 10510
rect 28809 10507 28875 10510
rect 34973 10570 35039 10573
rect 37406 10570 37412 10572
rect 34973 10568 37412 10570
rect 34973 10512 34978 10568
rect 35034 10512 37412 10568
rect 34973 10510 37412 10512
rect 34973 10507 35039 10510
rect 37406 10508 37412 10510
rect 37476 10508 37482 10572
rect 8150 10372 8156 10436
rect 8220 10434 8226 10436
rect 22185 10434 22251 10437
rect 8220 10432 22251 10434
rect 8220 10376 22190 10432
rect 22246 10376 22251 10432
rect 8220 10374 22251 10376
rect 8220 10372 8226 10374
rect 22185 10371 22251 10374
rect 25998 10372 26004 10436
rect 26068 10434 26074 10436
rect 30465 10434 30531 10437
rect 26068 10432 30531 10434
rect 26068 10376 30470 10432
rect 30526 10376 30531 10432
rect 26068 10374 30531 10376
rect 26068 10372 26074 10374
rect 30465 10371 30531 10374
rect 5130 10368 5446 10369
rect 5130 10304 5136 10368
rect 5200 10304 5216 10368
rect 5280 10304 5296 10368
rect 5360 10304 5376 10368
rect 5440 10304 5446 10368
rect 5130 10303 5446 10304
rect 35850 10368 36166 10369
rect 35850 10304 35856 10368
rect 35920 10304 35936 10368
rect 36000 10304 36016 10368
rect 36080 10304 36096 10368
rect 36160 10304 36166 10368
rect 35850 10303 36166 10304
rect 66570 10368 66886 10369
rect 66570 10304 66576 10368
rect 66640 10304 66656 10368
rect 66720 10304 66736 10368
rect 66800 10304 66816 10368
rect 66880 10304 66886 10368
rect 66570 10303 66886 10304
rect 21173 10300 21239 10301
rect 21173 10298 21220 10300
rect 21128 10296 21220 10298
rect 21128 10240 21178 10296
rect 21128 10238 21220 10240
rect 21173 10236 21220 10238
rect 21284 10236 21290 10300
rect 21173 10235 21239 10236
rect 17217 10162 17283 10165
rect 27613 10162 27679 10165
rect 17217 10160 27679 10162
rect 17217 10104 17222 10160
rect 17278 10104 27618 10160
rect 27674 10104 27679 10160
rect 17217 10102 27679 10104
rect 17217 10099 17283 10102
rect 27613 10099 27679 10102
rect 30373 10162 30439 10165
rect 30782 10162 30788 10164
rect 30373 10160 30788 10162
rect 30373 10104 30378 10160
rect 30434 10104 30788 10160
rect 30373 10102 30788 10104
rect 30373 10099 30439 10102
rect 30782 10100 30788 10102
rect 30852 10100 30858 10164
rect 33593 10162 33659 10165
rect 37222 10162 37228 10164
rect 33593 10160 37228 10162
rect 33593 10104 33598 10160
rect 33654 10104 37228 10160
rect 33593 10102 37228 10104
rect 33593 10099 33659 10102
rect 37222 10100 37228 10102
rect 37292 10100 37298 10164
rect 10174 9964 10180 10028
rect 10244 10026 10250 10028
rect 20437 10026 20503 10029
rect 10244 10024 20503 10026
rect 10244 9968 20442 10024
rect 20498 9968 20503 10024
rect 10244 9966 20503 9968
rect 10244 9964 10250 9966
rect 20437 9963 20503 9966
rect 20846 9964 20852 10028
rect 20916 10026 20922 10028
rect 23473 10026 23539 10029
rect 20916 10024 23539 10026
rect 20916 9968 23478 10024
rect 23534 9968 23539 10024
rect 20916 9966 23539 9968
rect 20916 9964 20922 9966
rect 23473 9963 23539 9966
rect 24853 10026 24919 10029
rect 27705 10026 27771 10029
rect 24853 10024 27771 10026
rect 24853 9968 24858 10024
rect 24914 9968 27710 10024
rect 27766 9968 27771 10024
rect 24853 9966 27771 9968
rect 24853 9963 24919 9966
rect 27705 9963 27771 9966
rect 28022 9964 28028 10028
rect 28092 10026 28098 10028
rect 36629 10026 36695 10029
rect 28092 10024 36695 10026
rect 28092 9968 36634 10024
rect 36690 9968 36695 10024
rect 28092 9966 36695 9968
rect 28092 9964 28098 9966
rect 36629 9963 36695 9966
rect 10726 9828 10732 9892
rect 10796 9890 10802 9892
rect 20805 9890 20871 9893
rect 30557 9890 30623 9893
rect 35893 9890 35959 9893
rect 10796 9888 20871 9890
rect 10796 9832 20810 9888
rect 20866 9832 20871 9888
rect 10796 9830 20871 9832
rect 10796 9828 10802 9830
rect 20805 9827 20871 9830
rect 21038 9888 30623 9890
rect 21038 9832 30562 9888
rect 30618 9832 30623 9888
rect 21038 9830 30623 9832
rect 5790 9824 6106 9825
rect 5790 9760 5796 9824
rect 5860 9760 5876 9824
rect 5940 9760 5956 9824
rect 6020 9760 6036 9824
rect 6100 9760 6106 9824
rect 5790 9759 6106 9760
rect 19609 9754 19675 9757
rect 19742 9754 19748 9756
rect 19609 9752 19748 9754
rect 19609 9696 19614 9752
rect 19670 9696 19748 9752
rect 19609 9694 19748 9696
rect 19609 9691 19675 9694
rect 19742 9692 19748 9694
rect 19812 9692 19818 9756
rect 20478 9692 20484 9756
rect 20548 9754 20554 9756
rect 21038 9754 21098 9830
rect 30557 9827 30623 9830
rect 30790 9888 35959 9890
rect 30790 9832 35898 9888
rect 35954 9832 35959 9888
rect 30790 9830 35959 9832
rect 20548 9694 21098 9754
rect 20548 9692 20554 9694
rect 21398 9692 21404 9756
rect 21468 9754 21474 9756
rect 21817 9754 21883 9757
rect 21468 9752 21883 9754
rect 21468 9696 21822 9752
rect 21878 9696 21883 9752
rect 21468 9694 21883 9696
rect 21468 9692 21474 9694
rect 21817 9691 21883 9694
rect 24158 9692 24164 9756
rect 24228 9754 24234 9756
rect 24669 9754 24735 9757
rect 24228 9752 24735 9754
rect 24228 9696 24674 9752
rect 24730 9696 24735 9752
rect 24228 9694 24735 9696
rect 24228 9692 24234 9694
rect 24669 9691 24735 9694
rect 26182 9692 26188 9756
rect 26252 9754 26258 9756
rect 26325 9754 26391 9757
rect 26252 9752 26391 9754
rect 26252 9696 26330 9752
rect 26386 9696 26391 9752
rect 26252 9694 26391 9696
rect 26252 9692 26258 9694
rect 26325 9691 26391 9694
rect 29126 9692 29132 9756
rect 29196 9754 29202 9756
rect 30790 9754 30850 9830
rect 35893 9827 35959 9830
rect 36510 9824 36826 9825
rect 36510 9760 36516 9824
rect 36580 9760 36596 9824
rect 36660 9760 36676 9824
rect 36740 9760 36756 9824
rect 36820 9760 36826 9824
rect 36510 9759 36826 9760
rect 67230 9824 67546 9825
rect 67230 9760 67236 9824
rect 67300 9760 67316 9824
rect 67380 9760 67396 9824
rect 67460 9760 67476 9824
rect 67540 9760 67546 9824
rect 67230 9759 67546 9760
rect 32765 9754 32831 9757
rect 29196 9694 30850 9754
rect 30974 9752 32831 9754
rect 30974 9696 32770 9752
rect 32826 9696 32831 9752
rect 30974 9694 32831 9696
rect 29196 9692 29202 9694
rect 24209 9618 24275 9621
rect 24342 9618 24348 9620
rect 24209 9616 24348 9618
rect 24209 9560 24214 9616
rect 24270 9560 24348 9616
rect 24209 9558 24348 9560
rect 24209 9555 24275 9558
rect 24342 9556 24348 9558
rect 24412 9556 24418 9620
rect 28993 9618 29059 9621
rect 29310 9618 29316 9620
rect 28993 9616 29316 9618
rect 28993 9560 28998 9616
rect 29054 9560 29316 9616
rect 28993 9558 29316 9560
rect 28993 9555 29059 9558
rect 29310 9556 29316 9558
rect 29380 9556 29386 9620
rect 29678 9556 29684 9620
rect 29748 9618 29754 9620
rect 30974 9618 31034 9694
rect 32765 9691 32831 9694
rect 34237 9756 34303 9757
rect 34237 9752 34284 9756
rect 34348 9754 34354 9756
rect 34237 9696 34242 9752
rect 34237 9692 34284 9696
rect 34348 9694 34394 9754
rect 34348 9692 34354 9694
rect 34237 9691 34303 9692
rect 29748 9558 31034 9618
rect 29748 9556 29754 9558
rect 31150 9556 31156 9620
rect 31220 9618 31226 9620
rect 31569 9618 31635 9621
rect 31220 9616 31635 9618
rect 31220 9560 31574 9616
rect 31630 9560 31635 9616
rect 31220 9558 31635 9560
rect 31220 9556 31226 9558
rect 31569 9555 31635 9558
rect 32622 9556 32628 9620
rect 32692 9618 32698 9620
rect 33225 9618 33291 9621
rect 32692 9616 33291 9618
rect 32692 9560 33230 9616
rect 33286 9560 33291 9616
rect 32692 9558 33291 9560
rect 32692 9556 32698 9558
rect 33225 9555 33291 9558
rect 13670 9420 13676 9484
rect 13740 9482 13746 9484
rect 25957 9482 26023 9485
rect 13740 9480 26023 9482
rect 13740 9424 25962 9480
rect 26018 9424 26023 9480
rect 13740 9422 26023 9424
rect 13740 9420 13746 9422
rect 25957 9419 26023 9422
rect 30966 9420 30972 9484
rect 31036 9482 31042 9484
rect 31109 9482 31175 9485
rect 31036 9480 31175 9482
rect 31036 9424 31114 9480
rect 31170 9424 31175 9480
rect 31036 9422 31175 9424
rect 31036 9420 31042 9422
rect 31109 9419 31175 9422
rect 32438 9420 32444 9484
rect 32508 9482 32514 9484
rect 36353 9482 36419 9485
rect 32508 9480 36419 9482
rect 32508 9424 36358 9480
rect 36414 9424 36419 9480
rect 32508 9422 36419 9424
rect 32508 9420 32514 9422
rect 36353 9419 36419 9422
rect 12985 9346 13051 9349
rect 19425 9346 19491 9349
rect 12985 9344 19491 9346
rect 12985 9288 12990 9344
rect 13046 9288 19430 9344
rect 19486 9288 19491 9344
rect 12985 9286 19491 9288
rect 12985 9283 13051 9286
rect 19425 9283 19491 9286
rect 27102 9284 27108 9348
rect 27172 9346 27178 9348
rect 34973 9346 35039 9349
rect 27172 9344 35039 9346
rect 27172 9288 34978 9344
rect 35034 9288 35039 9344
rect 27172 9286 35039 9288
rect 27172 9284 27178 9286
rect 34973 9283 35039 9286
rect 5130 9280 5446 9281
rect 5130 9216 5136 9280
rect 5200 9216 5216 9280
rect 5280 9216 5296 9280
rect 5360 9216 5376 9280
rect 5440 9216 5446 9280
rect 5130 9215 5446 9216
rect 35850 9280 36166 9281
rect 35850 9216 35856 9280
rect 35920 9216 35936 9280
rect 36000 9216 36016 9280
rect 36080 9216 36096 9280
rect 36160 9216 36166 9280
rect 35850 9215 36166 9216
rect 66570 9280 66886 9281
rect 66570 9216 66576 9280
rect 66640 9216 66656 9280
rect 66720 9216 66736 9280
rect 66800 9216 66816 9280
rect 66880 9216 66886 9280
rect 66570 9215 66886 9216
rect 17166 9148 17172 9212
rect 17236 9210 17242 9212
rect 17953 9210 18019 9213
rect 19241 9212 19307 9213
rect 19190 9210 19196 9212
rect 17236 9208 18019 9210
rect 17236 9152 17958 9208
rect 18014 9152 18019 9208
rect 17236 9150 18019 9152
rect 19150 9150 19196 9210
rect 19260 9208 19307 9212
rect 19302 9152 19307 9208
rect 17236 9148 17242 9150
rect 17953 9147 18019 9150
rect 19190 9148 19196 9150
rect 19260 9148 19307 9152
rect 27286 9148 27292 9212
rect 27356 9210 27362 9212
rect 31293 9210 31359 9213
rect 33685 9210 33751 9213
rect 33961 9212 34027 9213
rect 27356 9208 33751 9210
rect 27356 9152 31298 9208
rect 31354 9152 33690 9208
rect 33746 9152 33751 9208
rect 27356 9150 33751 9152
rect 27356 9148 27362 9150
rect 19241 9147 19307 9148
rect 31293 9147 31359 9150
rect 33685 9147 33751 9150
rect 33910 9148 33916 9212
rect 33980 9210 34027 9212
rect 35157 9210 35223 9213
rect 33980 9208 35223 9210
rect 34022 9152 35162 9208
rect 35218 9152 35223 9208
rect 33980 9150 35223 9152
rect 33980 9148 34027 9150
rect 33961 9147 34027 9148
rect 35157 9147 35223 9150
rect 16798 9012 16804 9076
rect 16868 9074 16874 9076
rect 34605 9074 34671 9077
rect 16868 9072 34671 9074
rect 16868 9016 34610 9072
rect 34666 9016 34671 9072
rect 16868 9014 34671 9016
rect 16868 9012 16874 9014
rect 34605 9011 34671 9014
rect 36302 9012 36308 9076
rect 36372 9074 36378 9076
rect 38193 9074 38259 9077
rect 36372 9072 38259 9074
rect 36372 9016 38198 9072
rect 38254 9016 38259 9072
rect 36372 9014 38259 9016
rect 36372 9012 36378 9014
rect 38193 9011 38259 9014
rect 10409 8938 10475 8941
rect 23013 8938 23079 8941
rect 10409 8936 23079 8938
rect 10409 8880 10414 8936
rect 10470 8880 23018 8936
rect 23074 8880 23079 8936
rect 10409 8878 23079 8880
rect 10409 8875 10475 8878
rect 23013 8875 23079 8878
rect 24894 8876 24900 8940
rect 24964 8938 24970 8940
rect 25865 8938 25931 8941
rect 24964 8936 25931 8938
rect 24964 8880 25870 8936
rect 25926 8880 25931 8936
rect 24964 8878 25931 8880
rect 24964 8876 24970 8878
rect 25865 8875 25931 8878
rect 27470 8876 27476 8940
rect 27540 8938 27546 8940
rect 33133 8938 33199 8941
rect 35249 8940 35315 8941
rect 27540 8936 33199 8938
rect 27540 8880 33138 8936
rect 33194 8880 33199 8936
rect 27540 8878 33199 8880
rect 27540 8876 27546 8878
rect 33133 8875 33199 8878
rect 35198 8876 35204 8940
rect 35268 8938 35315 8940
rect 35268 8936 35360 8938
rect 35310 8880 35360 8936
rect 35268 8878 35360 8880
rect 35268 8876 35315 8878
rect 35249 8875 35315 8876
rect 18086 8740 18092 8804
rect 18156 8802 18162 8804
rect 18597 8802 18663 8805
rect 18156 8800 18663 8802
rect 18156 8744 18602 8800
rect 18658 8744 18663 8800
rect 18156 8742 18663 8744
rect 18156 8740 18162 8742
rect 18597 8739 18663 8742
rect 19425 8802 19491 8805
rect 24301 8802 24367 8805
rect 36261 8802 36327 8805
rect 19425 8800 36327 8802
rect 19425 8744 19430 8800
rect 19486 8744 24306 8800
rect 24362 8744 36266 8800
rect 36322 8744 36327 8800
rect 19425 8742 36327 8744
rect 19425 8739 19491 8742
rect 24301 8739 24367 8742
rect 36261 8739 36327 8742
rect 5790 8736 6106 8737
rect 5790 8672 5796 8736
rect 5860 8672 5876 8736
rect 5940 8672 5956 8736
rect 6020 8672 6036 8736
rect 6100 8672 6106 8736
rect 5790 8671 6106 8672
rect 36510 8736 36826 8737
rect 36510 8672 36516 8736
rect 36580 8672 36596 8736
rect 36660 8672 36676 8736
rect 36740 8672 36756 8736
rect 36820 8672 36826 8736
rect 36510 8671 36826 8672
rect 67230 8736 67546 8737
rect 67230 8672 67236 8736
rect 67300 8672 67316 8736
rect 67380 8672 67396 8736
rect 67460 8672 67476 8736
rect 67540 8672 67546 8736
rect 67230 8671 67546 8672
rect 12249 8666 12315 8669
rect 20345 8666 20411 8669
rect 12249 8664 20411 8666
rect 12249 8608 12254 8664
rect 12310 8608 20350 8664
rect 20406 8608 20411 8664
rect 12249 8606 20411 8608
rect 12249 8603 12315 8606
rect 20345 8603 20411 8606
rect 24393 8666 24459 8669
rect 27429 8666 27495 8669
rect 24393 8664 27495 8666
rect 24393 8608 24398 8664
rect 24454 8608 27434 8664
rect 27490 8608 27495 8664
rect 24393 8606 27495 8608
rect 24393 8603 24459 8606
rect 27429 8603 27495 8606
rect 27654 8604 27660 8668
rect 27724 8666 27730 8668
rect 32213 8666 32279 8669
rect 27724 8664 32279 8666
rect 27724 8608 32218 8664
rect 32274 8608 32279 8664
rect 27724 8606 32279 8608
rect 27724 8604 27730 8606
rect 32213 8603 32279 8606
rect 35065 8666 35131 8669
rect 35566 8666 35572 8668
rect 35065 8664 35572 8666
rect 35065 8608 35070 8664
rect 35126 8608 35572 8664
rect 35065 8606 35572 8608
rect 35065 8603 35131 8606
rect 35566 8604 35572 8606
rect 35636 8604 35642 8668
rect 18137 8530 18203 8533
rect 20110 8530 20116 8532
rect 18137 8528 20116 8530
rect 18137 8472 18142 8528
rect 18198 8472 20116 8528
rect 18137 8470 20116 8472
rect 18137 8467 18203 8470
rect 20110 8468 20116 8470
rect 20180 8468 20186 8532
rect 23054 8468 23060 8532
rect 23124 8530 23130 8532
rect 28441 8530 28507 8533
rect 23124 8528 28507 8530
rect 23124 8472 28446 8528
rect 28502 8472 28507 8528
rect 23124 8470 28507 8472
rect 23124 8468 23130 8470
rect 28441 8467 28507 8470
rect 30598 8468 30604 8532
rect 30668 8530 30674 8532
rect 33041 8530 33107 8533
rect 30668 8528 33107 8530
rect 30668 8472 33046 8528
rect 33102 8472 33107 8528
rect 30668 8470 33107 8472
rect 30668 8468 30674 8470
rect 33041 8467 33107 8470
rect 33225 8530 33291 8533
rect 33358 8530 33364 8532
rect 33225 8528 33364 8530
rect 33225 8472 33230 8528
rect 33286 8472 33364 8528
rect 33225 8470 33364 8472
rect 33225 8467 33291 8470
rect 33358 8468 33364 8470
rect 33428 8468 33434 8532
rect 9990 8332 9996 8396
rect 10060 8394 10066 8396
rect 18137 8394 18203 8397
rect 10060 8392 18203 8394
rect 10060 8336 18142 8392
rect 18198 8336 18203 8392
rect 10060 8334 18203 8336
rect 10060 8332 10066 8334
rect 18137 8331 18203 8334
rect 19558 8332 19564 8396
rect 19628 8394 19634 8396
rect 19885 8394 19951 8397
rect 19628 8392 19951 8394
rect 19628 8336 19890 8392
rect 19946 8336 19951 8392
rect 19628 8334 19951 8336
rect 19628 8332 19634 8334
rect 19885 8331 19951 8334
rect 20529 8394 20595 8397
rect 25313 8394 25379 8397
rect 20529 8392 25379 8394
rect 20529 8336 20534 8392
rect 20590 8336 25318 8392
rect 25374 8336 25379 8392
rect 20529 8334 25379 8336
rect 20529 8331 20595 8334
rect 25313 8331 25379 8334
rect 28206 8332 28212 8396
rect 28276 8394 28282 8396
rect 32489 8394 32555 8397
rect 28276 8392 32555 8394
rect 28276 8336 32494 8392
rect 32550 8336 32555 8392
rect 28276 8334 32555 8336
rect 28276 8332 28282 8334
rect 32489 8331 32555 8334
rect 32990 8332 32996 8396
rect 33060 8394 33066 8396
rect 33409 8394 33475 8397
rect 33060 8392 33475 8394
rect 33060 8336 33414 8392
rect 33470 8336 33475 8392
rect 33060 8334 33475 8336
rect 33060 8332 33066 8334
rect 33409 8331 33475 8334
rect 34830 8332 34836 8396
rect 34900 8394 34906 8396
rect 35525 8394 35591 8397
rect 34900 8392 35591 8394
rect 34900 8336 35530 8392
rect 35586 8336 35591 8392
rect 34900 8334 35591 8336
rect 34900 8332 34906 8334
rect 35525 8331 35591 8334
rect 17769 8258 17835 8261
rect 18270 8258 18276 8260
rect 17769 8256 18276 8258
rect 17769 8200 17774 8256
rect 17830 8200 18276 8256
rect 17769 8198 18276 8200
rect 17769 8195 17835 8198
rect 18270 8196 18276 8198
rect 18340 8196 18346 8260
rect 21173 8258 21239 8261
rect 24761 8258 24827 8261
rect 21173 8256 24827 8258
rect 21173 8200 21178 8256
rect 21234 8200 24766 8256
rect 24822 8200 24827 8256
rect 21173 8198 24827 8200
rect 21173 8195 21239 8198
rect 24761 8195 24827 8198
rect 27429 8258 27495 8261
rect 34789 8258 34855 8261
rect 27429 8256 34855 8258
rect 27429 8200 27434 8256
rect 27490 8200 34794 8256
rect 34850 8200 34855 8256
rect 27429 8198 34855 8200
rect 27429 8195 27495 8198
rect 34789 8195 34855 8198
rect 5130 8192 5446 8193
rect 5130 8128 5136 8192
rect 5200 8128 5216 8192
rect 5280 8128 5296 8192
rect 5360 8128 5376 8192
rect 5440 8128 5446 8192
rect 5130 8127 5446 8128
rect 35850 8192 36166 8193
rect 35850 8128 35856 8192
rect 35920 8128 35936 8192
rect 36000 8128 36016 8192
rect 36080 8128 36096 8192
rect 36160 8128 36166 8192
rect 35850 8127 36166 8128
rect 66570 8192 66886 8193
rect 66570 8128 66576 8192
rect 66640 8128 66656 8192
rect 66720 8128 66736 8192
rect 66800 8128 66816 8192
rect 66880 8128 66886 8192
rect 66570 8127 66886 8128
rect 22502 8060 22508 8124
rect 22572 8122 22578 8124
rect 24342 8122 24348 8124
rect 22572 8062 24348 8122
rect 22572 8060 22578 8062
rect 24342 8060 24348 8062
rect 24412 8122 24418 8124
rect 25865 8122 25931 8125
rect 24412 8120 25931 8122
rect 24412 8064 25870 8120
rect 25926 8064 25931 8120
rect 24412 8062 25931 8064
rect 24412 8060 24418 8062
rect 25865 8059 25931 8062
rect 28441 8122 28507 8125
rect 31937 8122 32003 8125
rect 28441 8120 32003 8122
rect 28441 8064 28446 8120
rect 28502 8064 31942 8120
rect 31998 8064 32003 8120
rect 28441 8062 32003 8064
rect 28441 8059 28507 8062
rect 31937 8059 32003 8062
rect 33174 8060 33180 8124
rect 33244 8122 33250 8124
rect 34237 8122 34303 8125
rect 33244 8120 34303 8122
rect 33244 8064 34242 8120
rect 34298 8064 34303 8120
rect 33244 8062 34303 8064
rect 33244 8060 33250 8062
rect 34237 8059 34303 8062
rect 22737 7986 22803 7989
rect 27061 7986 27127 7989
rect 30557 7986 30623 7989
rect 34329 7986 34395 7989
rect 22737 7984 27354 7986
rect 22737 7928 22742 7984
rect 22798 7928 27066 7984
rect 27122 7928 27354 7984
rect 22737 7926 27354 7928
rect 22737 7923 22803 7926
rect 27061 7923 27127 7926
rect 15009 7852 15075 7853
rect 14958 7850 14964 7852
rect 14918 7790 14964 7850
rect 15028 7848 15075 7852
rect 15070 7792 15075 7848
rect 14958 7788 14964 7790
rect 15028 7788 15075 7792
rect 15009 7787 15075 7788
rect 24761 7850 24827 7853
rect 25078 7850 25084 7852
rect 24761 7848 25084 7850
rect 24761 7792 24766 7848
rect 24822 7792 25084 7848
rect 24761 7790 25084 7792
rect 24761 7787 24827 7790
rect 25078 7788 25084 7790
rect 25148 7788 25154 7852
rect 27294 7850 27354 7926
rect 30557 7984 34395 7986
rect 30557 7928 30562 7984
rect 30618 7928 34334 7984
rect 34390 7928 34395 7984
rect 30557 7926 34395 7928
rect 30557 7923 30623 7926
rect 34329 7923 34395 7926
rect 34973 7986 35039 7989
rect 40217 7986 40283 7989
rect 34973 7984 40283 7986
rect 34973 7928 34978 7984
rect 35034 7928 40222 7984
rect 40278 7928 40283 7984
rect 34973 7926 40283 7928
rect 34973 7923 35039 7926
rect 40217 7923 40283 7926
rect 30465 7850 30531 7853
rect 27294 7848 30531 7850
rect 27294 7792 30470 7848
rect 30526 7792 30531 7848
rect 27294 7790 30531 7792
rect 30465 7787 30531 7790
rect 31937 7850 32003 7853
rect 34789 7850 34855 7853
rect 31937 7848 34855 7850
rect 31937 7792 31942 7848
rect 31998 7792 34794 7848
rect 34850 7792 34855 7848
rect 31937 7790 34855 7792
rect 31937 7787 32003 7790
rect 34789 7787 34855 7790
rect 41454 7788 41460 7852
rect 41524 7850 41530 7852
rect 41597 7850 41663 7853
rect 41524 7848 41663 7850
rect 41524 7792 41602 7848
rect 41658 7792 41663 7848
rect 41524 7790 41663 7792
rect 41524 7788 41530 7790
rect 41597 7787 41663 7790
rect 20989 7714 21055 7717
rect 23749 7714 23815 7717
rect 20989 7712 23815 7714
rect 20989 7656 20994 7712
rect 21050 7656 23754 7712
rect 23810 7656 23815 7712
rect 20989 7654 23815 7656
rect 20989 7651 21055 7654
rect 23749 7651 23815 7654
rect 24301 7714 24367 7717
rect 25037 7714 25103 7717
rect 24301 7712 25103 7714
rect 24301 7656 24306 7712
rect 24362 7656 25042 7712
rect 25098 7656 25103 7712
rect 24301 7654 25103 7656
rect 24301 7651 24367 7654
rect 25037 7651 25103 7654
rect 25681 7714 25747 7717
rect 25681 7712 31586 7714
rect 25681 7656 25686 7712
rect 25742 7656 31586 7712
rect 25681 7654 31586 7656
rect 25681 7651 25747 7654
rect 5790 7648 6106 7649
rect 5790 7584 5796 7648
rect 5860 7584 5876 7648
rect 5940 7584 5956 7648
rect 6020 7584 6036 7648
rect 6100 7584 6106 7648
rect 5790 7583 6106 7584
rect 17902 7516 17908 7580
rect 17972 7578 17978 7580
rect 20161 7578 20227 7581
rect 17972 7576 20227 7578
rect 17972 7520 20166 7576
rect 20222 7520 20227 7576
rect 17972 7518 20227 7520
rect 17972 7516 17978 7518
rect 20161 7515 20227 7518
rect 21449 7578 21515 7581
rect 22502 7578 22508 7580
rect 21449 7576 22508 7578
rect 21449 7520 21454 7576
rect 21510 7520 22508 7576
rect 21449 7518 22508 7520
rect 21449 7515 21515 7518
rect 22502 7516 22508 7518
rect 22572 7516 22578 7580
rect 24945 7578 25011 7581
rect 29269 7578 29335 7581
rect 31526 7580 31586 7654
rect 36510 7648 36826 7649
rect 36510 7584 36516 7648
rect 36580 7584 36596 7648
rect 36660 7584 36676 7648
rect 36740 7584 36756 7648
rect 36820 7584 36826 7648
rect 36510 7583 36826 7584
rect 67230 7648 67546 7649
rect 67230 7584 67236 7648
rect 67300 7584 67316 7648
rect 67380 7584 67396 7648
rect 67460 7584 67476 7648
rect 67540 7584 67546 7648
rect 67230 7583 67546 7584
rect 24945 7576 29335 7578
rect 24945 7520 24950 7576
rect 25006 7520 29274 7576
rect 29330 7520 29335 7576
rect 24945 7518 29335 7520
rect 24945 7515 25011 7518
rect 29269 7515 29335 7518
rect 31518 7516 31524 7580
rect 31588 7578 31594 7580
rect 31753 7578 31819 7581
rect 33869 7578 33935 7581
rect 31588 7576 31819 7578
rect 31588 7520 31758 7576
rect 31814 7520 31819 7576
rect 31588 7518 31819 7520
rect 31588 7516 31594 7518
rect 31753 7515 31819 7518
rect 32216 7576 33935 7578
rect 32216 7520 33874 7576
rect 33930 7520 33935 7576
rect 32216 7518 33935 7520
rect 32216 7445 32276 7518
rect 33869 7515 33935 7518
rect 35382 7516 35388 7580
rect 35452 7578 35458 7580
rect 35525 7578 35591 7581
rect 35452 7576 35591 7578
rect 35452 7520 35530 7576
rect 35586 7520 35591 7576
rect 35452 7518 35591 7520
rect 35452 7516 35458 7518
rect 35525 7515 35591 7518
rect 22461 7442 22527 7445
rect 25814 7442 25820 7444
rect 22461 7440 25820 7442
rect 22461 7384 22466 7440
rect 22522 7384 25820 7440
rect 22461 7382 25820 7384
rect 22461 7379 22527 7382
rect 25814 7380 25820 7382
rect 25884 7380 25890 7444
rect 30097 7442 30163 7445
rect 32213 7442 32279 7445
rect 30097 7440 32279 7442
rect 30097 7384 30102 7440
rect 30158 7384 32218 7440
rect 32274 7384 32279 7440
rect 30097 7382 32279 7384
rect 30097 7379 30163 7382
rect 32213 7379 32279 7382
rect 32806 7380 32812 7444
rect 32876 7442 32882 7444
rect 33409 7442 33475 7445
rect 32876 7440 33475 7442
rect 32876 7384 33414 7440
rect 33470 7384 33475 7440
rect 32876 7382 33475 7384
rect 32876 7380 32882 7382
rect 33409 7379 33475 7382
rect 12065 7306 12131 7309
rect 16757 7306 16823 7309
rect 12065 7304 16823 7306
rect 12065 7248 12070 7304
rect 12126 7248 16762 7304
rect 16818 7248 16823 7304
rect 12065 7246 16823 7248
rect 12065 7243 12131 7246
rect 16757 7243 16823 7246
rect 21173 7306 21239 7309
rect 24025 7306 24091 7309
rect 21173 7304 24091 7306
rect 21173 7248 21178 7304
rect 21234 7248 24030 7304
rect 24086 7248 24091 7304
rect 21173 7246 24091 7248
rect 21173 7243 21239 7246
rect 24025 7243 24091 7246
rect 28257 7306 28323 7309
rect 34881 7306 34947 7309
rect 28257 7304 34947 7306
rect 28257 7248 28262 7304
rect 28318 7248 34886 7304
rect 34942 7248 34947 7304
rect 28257 7246 34947 7248
rect 28257 7243 28323 7246
rect 34881 7243 34947 7246
rect 14273 7170 14339 7173
rect 20253 7170 20319 7173
rect 14273 7168 20319 7170
rect 14273 7112 14278 7168
rect 14334 7112 20258 7168
rect 20314 7112 20319 7168
rect 14273 7110 20319 7112
rect 14273 7107 14339 7110
rect 20253 7107 20319 7110
rect 21909 7170 21975 7173
rect 25998 7170 26004 7172
rect 21909 7168 26004 7170
rect 21909 7112 21914 7168
rect 21970 7112 26004 7168
rect 21909 7110 26004 7112
rect 21909 7107 21975 7110
rect 25998 7108 26004 7110
rect 26068 7108 26074 7172
rect 26141 7170 26207 7173
rect 28206 7170 28212 7172
rect 26141 7168 28212 7170
rect 26141 7112 26146 7168
rect 26202 7112 28212 7168
rect 26141 7110 28212 7112
rect 26141 7107 26207 7110
rect 28206 7108 28212 7110
rect 28276 7108 28282 7172
rect 29913 7170 29979 7173
rect 30373 7170 30439 7173
rect 31937 7170 32003 7173
rect 32213 7170 32279 7173
rect 29913 7168 32279 7170
rect 29913 7112 29918 7168
rect 29974 7112 30378 7168
rect 30434 7112 31942 7168
rect 31998 7112 32218 7168
rect 32274 7112 32279 7168
rect 29913 7110 32279 7112
rect 29913 7107 29979 7110
rect 30373 7107 30439 7110
rect 31937 7107 32003 7110
rect 32213 7107 32279 7110
rect 33041 7170 33107 7173
rect 33317 7170 33383 7173
rect 33041 7168 33383 7170
rect 33041 7112 33046 7168
rect 33102 7112 33322 7168
rect 33378 7112 33383 7168
rect 33041 7110 33383 7112
rect 33041 7107 33107 7110
rect 33317 7107 33383 7110
rect 33869 7172 33935 7173
rect 33869 7168 33916 7172
rect 33980 7170 33986 7172
rect 33869 7112 33874 7168
rect 33869 7108 33916 7112
rect 33980 7110 34026 7170
rect 33980 7108 33986 7110
rect 33869 7107 33935 7108
rect 5130 7104 5446 7105
rect 5130 7040 5136 7104
rect 5200 7040 5216 7104
rect 5280 7040 5296 7104
rect 5360 7040 5376 7104
rect 5440 7040 5446 7104
rect 5130 7039 5446 7040
rect 35850 7104 36166 7105
rect 35850 7040 35856 7104
rect 35920 7040 35936 7104
rect 36000 7040 36016 7104
rect 36080 7040 36096 7104
rect 36160 7040 36166 7104
rect 35850 7039 36166 7040
rect 66570 7104 66886 7105
rect 66570 7040 66576 7104
rect 66640 7040 66656 7104
rect 66720 7040 66736 7104
rect 66800 7040 66816 7104
rect 66880 7040 66886 7104
rect 66570 7039 66886 7040
rect 15142 6972 15148 7036
rect 15212 7034 15218 7036
rect 15377 7034 15443 7037
rect 15212 7032 15443 7034
rect 15212 6976 15382 7032
rect 15438 6976 15443 7032
rect 15212 6974 15443 6976
rect 15212 6972 15218 6974
rect 15377 6971 15443 6974
rect 22277 7034 22343 7037
rect 23841 7034 23907 7037
rect 29729 7034 29795 7037
rect 22277 7032 22800 7034
rect 22277 6976 22282 7032
rect 22338 6976 22800 7032
rect 22277 6974 22800 6976
rect 22277 6971 22343 6974
rect 22553 6900 22619 6901
rect 22502 6836 22508 6900
rect 22572 6898 22619 6900
rect 22740 6898 22800 6974
rect 23841 7032 29795 7034
rect 23841 6976 23846 7032
rect 23902 6976 29734 7032
rect 29790 6976 29795 7032
rect 23841 6974 29795 6976
rect 23841 6971 23907 6974
rect 29729 6971 29795 6974
rect 31293 7034 31359 7037
rect 31569 7034 31635 7037
rect 31293 7032 31635 7034
rect 31293 6976 31298 7032
rect 31354 6976 31574 7032
rect 31630 6976 31635 7032
rect 31293 6974 31635 6976
rect 31293 6971 31359 6974
rect 31569 6971 31635 6974
rect 32397 7034 32463 7037
rect 34329 7034 34395 7037
rect 32397 7032 34395 7034
rect 32397 6976 32402 7032
rect 32458 6976 34334 7032
rect 34390 6976 34395 7032
rect 32397 6974 34395 6976
rect 32397 6971 32463 6974
rect 34329 6971 34395 6974
rect 25773 6898 25839 6901
rect 22572 6896 22664 6898
rect 22614 6840 22664 6896
rect 22572 6838 22664 6840
rect 22740 6896 25839 6898
rect 22740 6840 25778 6896
rect 25834 6840 25839 6896
rect 22740 6838 25839 6840
rect 22572 6836 22619 6838
rect 22553 6835 22619 6836
rect 25773 6835 25839 6838
rect 26601 6898 26667 6901
rect 27286 6898 27292 6900
rect 26601 6896 27292 6898
rect 26601 6840 26606 6896
rect 26662 6840 27292 6896
rect 26601 6838 27292 6840
rect 26601 6835 26667 6838
rect 27286 6836 27292 6838
rect 27356 6836 27362 6900
rect 30741 6898 30807 6901
rect 36905 6898 36971 6901
rect 30741 6896 36971 6898
rect 30741 6840 30746 6896
rect 30802 6840 36910 6896
rect 36966 6840 36971 6896
rect 30741 6838 36971 6840
rect 30741 6835 30807 6838
rect 36905 6835 36971 6838
rect 22185 6762 22251 6765
rect 25497 6762 25563 6765
rect 25630 6762 25636 6764
rect 22185 6760 25636 6762
rect 22185 6704 22190 6760
rect 22246 6704 25502 6760
rect 25558 6704 25636 6760
rect 22185 6702 25636 6704
rect 22185 6699 22251 6702
rect 25497 6699 25563 6702
rect 25630 6700 25636 6702
rect 25700 6762 25706 6764
rect 28533 6762 28599 6765
rect 25700 6760 28599 6762
rect 25700 6704 28538 6760
rect 28594 6704 28599 6760
rect 25700 6702 28599 6704
rect 25700 6700 25706 6702
rect 28533 6699 28599 6702
rect 29729 6762 29795 6765
rect 32622 6762 32628 6764
rect 29729 6760 32628 6762
rect 29729 6704 29734 6760
rect 29790 6704 32628 6760
rect 29729 6702 32628 6704
rect 29729 6699 29795 6702
rect 32622 6700 32628 6702
rect 32692 6700 32698 6764
rect 18505 6626 18571 6629
rect 21449 6626 21515 6629
rect 29310 6626 29316 6628
rect 18505 6624 19258 6626
rect 18505 6568 18510 6624
rect 18566 6568 19258 6624
rect 18505 6566 19258 6568
rect 18505 6563 18571 6566
rect 5790 6560 6106 6561
rect 5790 6496 5796 6560
rect 5860 6496 5876 6560
rect 5940 6496 5956 6560
rect 6020 6496 6036 6560
rect 6100 6496 6106 6560
rect 5790 6495 6106 6496
rect 19198 6493 19258 6566
rect 21449 6624 29316 6626
rect 21449 6568 21454 6624
rect 21510 6568 29316 6624
rect 21449 6566 29316 6568
rect 21449 6563 21515 6566
rect 29310 6564 29316 6566
rect 29380 6564 29386 6628
rect 30925 6626 30991 6629
rect 34145 6626 34211 6629
rect 30925 6624 34211 6626
rect 30925 6568 30930 6624
rect 30986 6568 34150 6624
rect 34206 6568 34211 6624
rect 30925 6566 34211 6568
rect 30925 6563 30991 6566
rect 34145 6563 34211 6566
rect 36510 6560 36826 6561
rect 36510 6496 36516 6560
rect 36580 6496 36596 6560
rect 36660 6496 36676 6560
rect 36740 6496 36756 6560
rect 36820 6496 36826 6560
rect 36510 6495 36826 6496
rect 67230 6560 67546 6561
rect 67230 6496 67236 6560
rect 67300 6496 67316 6560
rect 67380 6496 67396 6560
rect 67460 6496 67476 6560
rect 67540 6496 67546 6560
rect 67230 6495 67546 6496
rect 19198 6488 19307 6493
rect 19198 6432 19246 6488
rect 19302 6432 19307 6488
rect 19198 6430 19307 6432
rect 19241 6427 19307 6430
rect 21357 6490 21423 6493
rect 23289 6490 23355 6493
rect 21357 6488 23355 6490
rect 21357 6432 21362 6488
rect 21418 6432 23294 6488
rect 23350 6432 23355 6488
rect 21357 6430 23355 6432
rect 21357 6427 21423 6430
rect 23289 6427 23355 6430
rect 23749 6490 23815 6493
rect 24393 6490 24459 6493
rect 24526 6490 24532 6492
rect 23749 6488 24226 6490
rect 23749 6432 23754 6488
rect 23810 6432 24226 6488
rect 23749 6430 24226 6432
rect 23749 6427 23815 6430
rect 14590 6292 14596 6356
rect 14660 6354 14666 6356
rect 24025 6354 24091 6357
rect 14660 6352 24091 6354
rect 14660 6296 24030 6352
rect 24086 6296 24091 6352
rect 14660 6294 24091 6296
rect 24166 6354 24226 6430
rect 24393 6488 24532 6490
rect 24393 6432 24398 6488
rect 24454 6432 24532 6488
rect 24393 6430 24532 6432
rect 24393 6427 24459 6430
rect 24526 6428 24532 6430
rect 24596 6428 24602 6492
rect 24669 6490 24735 6493
rect 31150 6490 31156 6492
rect 24669 6488 31156 6490
rect 24669 6432 24674 6488
rect 24730 6432 31156 6488
rect 24669 6430 31156 6432
rect 24669 6427 24735 6430
rect 31150 6428 31156 6430
rect 31220 6428 31226 6492
rect 31661 6490 31727 6493
rect 31526 6488 31727 6490
rect 31526 6432 31666 6488
rect 31722 6432 31727 6488
rect 31526 6430 31727 6432
rect 28441 6354 28507 6357
rect 24166 6352 28507 6354
rect 24166 6296 28446 6352
rect 28502 6296 28507 6352
rect 24166 6294 28507 6296
rect 14660 6292 14666 6294
rect 24025 6291 24091 6294
rect 28441 6291 28507 6294
rect 28625 6354 28691 6357
rect 31526 6354 31586 6430
rect 31661 6427 31727 6430
rect 34513 6354 34579 6357
rect 28625 6352 31586 6354
rect 28625 6296 28630 6352
rect 28686 6296 31586 6352
rect 28625 6294 31586 6296
rect 31710 6352 34579 6354
rect 31710 6296 34518 6352
rect 34574 6296 34579 6352
rect 31710 6294 34579 6296
rect 28625 6291 28691 6294
rect 18045 6218 18111 6221
rect 21214 6218 21220 6220
rect 18045 6216 21220 6218
rect 18045 6160 18050 6216
rect 18106 6160 21220 6216
rect 18045 6158 21220 6160
rect 18045 6155 18111 6158
rect 21214 6156 21220 6158
rect 21284 6218 21290 6220
rect 31710 6218 31770 6294
rect 34513 6291 34579 6294
rect 21284 6158 31770 6218
rect 31937 6218 32003 6221
rect 36905 6218 36971 6221
rect 31937 6216 36971 6218
rect 31937 6160 31942 6216
rect 31998 6160 36910 6216
rect 36966 6160 36971 6216
rect 31937 6158 36971 6160
rect 21284 6156 21290 6158
rect 31937 6155 32003 6158
rect 36905 6155 36971 6158
rect 18505 6082 18571 6085
rect 19149 6082 19215 6085
rect 18505 6080 19215 6082
rect 18505 6024 18510 6080
rect 18566 6024 19154 6080
rect 19210 6024 19215 6080
rect 18505 6022 19215 6024
rect 18505 6019 18571 6022
rect 19149 6019 19215 6022
rect 19333 6082 19399 6085
rect 19885 6082 19951 6085
rect 19333 6080 19951 6082
rect 19333 6024 19338 6080
rect 19394 6024 19890 6080
rect 19946 6024 19951 6080
rect 19333 6022 19951 6024
rect 19333 6019 19399 6022
rect 19885 6019 19951 6022
rect 25681 6082 25747 6085
rect 29913 6082 29979 6085
rect 25681 6080 29979 6082
rect 25681 6024 25686 6080
rect 25742 6024 29918 6080
rect 29974 6024 29979 6080
rect 25681 6022 29979 6024
rect 25681 6019 25747 6022
rect 29913 6019 29979 6022
rect 31753 6082 31819 6085
rect 35709 6082 35775 6085
rect 31753 6080 35775 6082
rect 31753 6024 31758 6080
rect 31814 6024 35714 6080
rect 35770 6024 35775 6080
rect 31753 6022 35775 6024
rect 31753 6019 31819 6022
rect 35709 6019 35775 6022
rect 5130 6016 5446 6017
rect 5130 5952 5136 6016
rect 5200 5952 5216 6016
rect 5280 5952 5296 6016
rect 5360 5952 5376 6016
rect 5440 5952 5446 6016
rect 5130 5951 5446 5952
rect 35850 6016 36166 6017
rect 35850 5952 35856 6016
rect 35920 5952 35936 6016
rect 36000 5952 36016 6016
rect 36080 5952 36096 6016
rect 36160 5952 36166 6016
rect 35850 5951 36166 5952
rect 66570 6016 66886 6017
rect 66570 5952 66576 6016
rect 66640 5952 66656 6016
rect 66720 5952 66736 6016
rect 66800 5952 66816 6016
rect 66880 5952 66886 6016
rect 66570 5951 66886 5952
rect 11881 5946 11947 5949
rect 16297 5946 16363 5949
rect 11881 5944 16363 5946
rect 11881 5888 11886 5944
rect 11942 5888 16302 5944
rect 16358 5888 16363 5944
rect 11881 5886 16363 5888
rect 11881 5883 11947 5886
rect 16297 5883 16363 5886
rect 17125 5946 17191 5949
rect 20437 5946 20503 5949
rect 17125 5944 20503 5946
rect 17125 5888 17130 5944
rect 17186 5888 20442 5944
rect 20498 5888 20503 5944
rect 17125 5886 20503 5888
rect 17125 5883 17191 5886
rect 20437 5883 20503 5886
rect 24025 5946 24091 5949
rect 26918 5946 26924 5948
rect 24025 5944 26924 5946
rect 24025 5888 24030 5944
rect 24086 5888 26924 5944
rect 24025 5886 26924 5888
rect 24025 5883 24091 5886
rect 26918 5884 26924 5886
rect 26988 5884 26994 5948
rect 29545 5946 29611 5949
rect 29545 5944 35634 5946
rect 29545 5888 29550 5944
rect 29606 5888 35634 5944
rect 29545 5886 35634 5888
rect 29545 5883 29611 5886
rect 14825 5810 14891 5813
rect 17769 5810 17835 5813
rect 14825 5808 17835 5810
rect 14825 5752 14830 5808
rect 14886 5752 17774 5808
rect 17830 5752 17835 5808
rect 14825 5750 17835 5752
rect 14825 5747 14891 5750
rect 17769 5747 17835 5750
rect 20805 5810 20871 5813
rect 27337 5810 27403 5813
rect 27470 5810 27476 5812
rect 20805 5808 25146 5810
rect 20805 5752 20810 5808
rect 20866 5752 25146 5808
rect 20805 5750 25146 5752
rect 20805 5747 20871 5750
rect 25086 5677 25146 5750
rect 27337 5808 27476 5810
rect 27337 5752 27342 5808
rect 27398 5752 27476 5808
rect 27337 5750 27476 5752
rect 27337 5747 27403 5750
rect 27470 5748 27476 5750
rect 27540 5748 27546 5812
rect 29085 5810 29151 5813
rect 29453 5810 29519 5813
rect 31518 5810 31524 5812
rect 29085 5808 29332 5810
rect 29085 5752 29090 5808
rect 29146 5752 29332 5808
rect 29085 5750 29332 5752
rect 29085 5747 29151 5750
rect 10961 5674 11027 5677
rect 16573 5674 16639 5677
rect 19241 5676 19307 5677
rect 19190 5674 19196 5676
rect 10961 5672 16639 5674
rect 10961 5616 10966 5672
rect 11022 5616 16578 5672
rect 16634 5616 16639 5672
rect 10961 5614 16639 5616
rect 19150 5614 19196 5674
rect 19260 5672 19307 5676
rect 20805 5676 20871 5677
rect 23013 5676 23079 5677
rect 24117 5676 24183 5677
rect 25086 5676 25195 5677
rect 20805 5674 20852 5676
rect 19302 5616 19307 5672
rect 10961 5611 11027 5614
rect 16573 5611 16639 5614
rect 19190 5612 19196 5614
rect 19260 5612 19307 5616
rect 20760 5672 20852 5674
rect 20760 5616 20810 5672
rect 20760 5614 20852 5616
rect 19241 5611 19307 5612
rect 20805 5612 20852 5614
rect 20916 5612 20922 5676
rect 23013 5674 23060 5676
rect 22968 5672 23060 5674
rect 22968 5616 23018 5672
rect 22968 5614 23060 5616
rect 23013 5612 23060 5614
rect 23124 5612 23130 5676
rect 24117 5674 24164 5676
rect 24072 5672 24164 5674
rect 24072 5616 24122 5672
rect 24072 5614 24164 5616
rect 24117 5612 24164 5614
rect 24228 5612 24234 5676
rect 25078 5674 25084 5676
rect 25038 5614 25084 5674
rect 25148 5672 25195 5676
rect 25190 5616 25195 5672
rect 25078 5612 25084 5614
rect 25148 5612 25195 5616
rect 20805 5611 20871 5612
rect 23013 5611 23079 5612
rect 24117 5611 24183 5612
rect 25129 5611 25195 5612
rect 25497 5674 25563 5677
rect 27429 5674 27495 5677
rect 25497 5672 27495 5674
rect 25497 5616 25502 5672
rect 25558 5616 27434 5672
rect 27490 5616 27495 5672
rect 25497 5614 27495 5616
rect 25497 5611 25563 5614
rect 27429 5611 27495 5614
rect 29126 5612 29132 5676
rect 29196 5612 29202 5676
rect 15561 5538 15627 5541
rect 15694 5538 15700 5540
rect 15561 5536 15700 5538
rect 15561 5480 15566 5536
rect 15622 5480 15700 5536
rect 15561 5478 15700 5480
rect 15561 5475 15627 5478
rect 15694 5476 15700 5478
rect 15764 5476 15770 5540
rect 15837 5538 15903 5541
rect 17493 5538 17559 5541
rect 15837 5536 17559 5538
rect 15837 5480 15842 5536
rect 15898 5480 17498 5536
rect 17554 5480 17559 5536
rect 15837 5478 17559 5480
rect 15837 5475 15903 5478
rect 17493 5475 17559 5478
rect 18505 5538 18571 5541
rect 22461 5538 22527 5541
rect 18505 5536 22527 5538
rect 18505 5480 18510 5536
rect 18566 5480 22466 5536
rect 22522 5480 22527 5536
rect 18505 5478 22527 5480
rect 18505 5475 18571 5478
rect 22461 5475 22527 5478
rect 23381 5538 23447 5541
rect 27613 5538 27679 5541
rect 23381 5536 27679 5538
rect 23381 5480 23386 5536
rect 23442 5480 27618 5536
rect 27674 5480 27679 5536
rect 23381 5478 27679 5480
rect 23381 5475 23447 5478
rect 27613 5475 27679 5478
rect 27889 5538 27955 5541
rect 29134 5538 29194 5612
rect 27889 5536 29194 5538
rect 27889 5480 27894 5536
rect 27950 5480 29194 5536
rect 27889 5478 29194 5480
rect 29272 5538 29332 5750
rect 29453 5808 31524 5810
rect 29453 5752 29458 5808
rect 29514 5752 31524 5808
rect 29453 5750 31524 5752
rect 29453 5747 29519 5750
rect 31518 5748 31524 5750
rect 31588 5748 31594 5812
rect 31661 5810 31727 5813
rect 34421 5810 34487 5813
rect 31661 5808 34487 5810
rect 31661 5752 31666 5808
rect 31722 5752 34426 5808
rect 34482 5752 34487 5808
rect 31661 5750 34487 5752
rect 35574 5810 35634 5886
rect 35709 5810 35775 5813
rect 35574 5808 35775 5810
rect 35574 5752 35714 5808
rect 35770 5752 35775 5808
rect 35574 5750 35775 5752
rect 31661 5747 31727 5750
rect 34421 5747 34487 5750
rect 35709 5747 35775 5750
rect 29637 5674 29703 5677
rect 32581 5674 32647 5677
rect 36445 5674 36511 5677
rect 29637 5672 36511 5674
rect 29637 5616 29642 5672
rect 29698 5616 32586 5672
rect 32642 5616 36450 5672
rect 36506 5616 36511 5672
rect 29637 5614 36511 5616
rect 29637 5611 29703 5614
rect 32581 5611 32647 5614
rect 36445 5611 36511 5614
rect 31661 5538 31727 5541
rect 29272 5536 31727 5538
rect 29272 5480 31666 5536
rect 31722 5480 31727 5536
rect 29272 5478 31727 5480
rect 27889 5475 27955 5478
rect 31661 5475 31727 5478
rect 32029 5538 32095 5541
rect 32949 5538 33015 5541
rect 35433 5540 35499 5541
rect 32029 5536 33015 5538
rect 32029 5480 32034 5536
rect 32090 5480 32954 5536
rect 33010 5480 33015 5536
rect 32029 5478 33015 5480
rect 32029 5475 32095 5478
rect 32949 5475 33015 5478
rect 35382 5476 35388 5540
rect 35452 5538 35499 5540
rect 35893 5538 35959 5541
rect 35452 5536 35959 5538
rect 35494 5480 35898 5536
rect 35954 5480 35959 5536
rect 35452 5478 35959 5480
rect 35452 5476 35499 5478
rect 35433 5475 35499 5476
rect 35893 5475 35959 5478
rect 5790 5472 6106 5473
rect 5790 5408 5796 5472
rect 5860 5408 5876 5472
rect 5940 5408 5956 5472
rect 6020 5408 6036 5472
rect 6100 5408 6106 5472
rect 5790 5407 6106 5408
rect 36510 5472 36826 5473
rect 36510 5408 36516 5472
rect 36580 5408 36596 5472
rect 36660 5408 36676 5472
rect 36740 5408 36756 5472
rect 36820 5408 36826 5472
rect 36510 5407 36826 5408
rect 67230 5472 67546 5473
rect 67230 5408 67236 5472
rect 67300 5408 67316 5472
rect 67380 5408 67396 5472
rect 67460 5408 67476 5472
rect 67540 5408 67546 5472
rect 67230 5407 67546 5408
rect 9305 5402 9371 5405
rect 17902 5402 17908 5404
rect 9305 5400 17908 5402
rect 9305 5344 9310 5400
rect 9366 5344 17908 5400
rect 9305 5342 17908 5344
rect 9305 5339 9371 5342
rect 17902 5340 17908 5342
rect 17972 5340 17978 5404
rect 18321 5402 18387 5405
rect 19057 5402 19123 5405
rect 18321 5400 19123 5402
rect 18321 5344 18326 5400
rect 18382 5344 19062 5400
rect 19118 5344 19123 5400
rect 18321 5342 19123 5344
rect 18321 5339 18387 5342
rect 19057 5339 19123 5342
rect 20897 5402 20963 5405
rect 24669 5402 24735 5405
rect 20897 5400 24735 5402
rect 20897 5344 20902 5400
rect 20958 5344 24674 5400
rect 24730 5344 24735 5400
rect 20897 5342 24735 5344
rect 20897 5339 20963 5342
rect 24669 5339 24735 5342
rect 25497 5402 25563 5405
rect 32438 5402 32444 5404
rect 25497 5400 32444 5402
rect 25497 5344 25502 5400
rect 25558 5344 32444 5400
rect 25497 5342 32444 5344
rect 25497 5339 25563 5342
rect 32438 5340 32444 5342
rect 32508 5340 32514 5404
rect 10133 5266 10199 5269
rect 14273 5266 14339 5269
rect 10133 5264 14339 5266
rect 10133 5208 10138 5264
rect 10194 5208 14278 5264
rect 14334 5208 14339 5264
rect 10133 5206 14339 5208
rect 10133 5203 10199 5206
rect 14273 5203 14339 5206
rect 15009 5266 15075 5269
rect 21357 5266 21423 5269
rect 15009 5264 21423 5266
rect 15009 5208 15014 5264
rect 15070 5208 21362 5264
rect 21418 5208 21423 5264
rect 15009 5206 21423 5208
rect 15009 5203 15075 5206
rect 21357 5203 21423 5206
rect 24853 5266 24919 5269
rect 27654 5266 27660 5268
rect 24853 5264 27660 5266
rect 24853 5208 24858 5264
rect 24914 5208 27660 5264
rect 24853 5206 27660 5208
rect 24853 5203 24919 5206
rect 27654 5204 27660 5206
rect 27724 5204 27730 5268
rect 28349 5266 28415 5269
rect 30598 5266 30604 5268
rect 28349 5264 30604 5266
rect 28349 5208 28354 5264
rect 28410 5208 30604 5264
rect 28349 5206 30604 5208
rect 28349 5203 28415 5206
rect 30598 5204 30604 5206
rect 30668 5204 30674 5268
rect 30833 5266 30899 5269
rect 37365 5266 37431 5269
rect 30833 5264 37431 5266
rect 30833 5208 30838 5264
rect 30894 5208 37370 5264
rect 37426 5208 37431 5264
rect 30833 5206 37431 5208
rect 30833 5203 30899 5206
rect 37365 5203 37431 5206
rect 14641 5130 14707 5133
rect 14774 5130 14780 5132
rect 14641 5128 14780 5130
rect 14641 5072 14646 5128
rect 14702 5072 14780 5128
rect 14641 5070 14780 5072
rect 14641 5067 14707 5070
rect 14774 5068 14780 5070
rect 14844 5068 14850 5132
rect 15837 5130 15903 5133
rect 19149 5130 19215 5133
rect 15837 5128 19215 5130
rect 15837 5072 15842 5128
rect 15898 5072 19154 5128
rect 19210 5072 19215 5128
rect 15837 5070 19215 5072
rect 15837 5067 15903 5070
rect 19149 5067 19215 5070
rect 21817 5130 21883 5133
rect 27521 5130 27587 5133
rect 21817 5128 27587 5130
rect 21817 5072 21822 5128
rect 21878 5072 27526 5128
rect 27582 5072 27587 5128
rect 21817 5070 27587 5072
rect 21817 5067 21883 5070
rect 27521 5067 27587 5070
rect 29269 5130 29335 5133
rect 30097 5130 30163 5133
rect 34789 5132 34855 5133
rect 34789 5130 34836 5132
rect 29269 5128 30163 5130
rect 29269 5072 29274 5128
rect 29330 5072 30102 5128
rect 30158 5072 30163 5128
rect 29269 5070 30163 5072
rect 34744 5128 34836 5130
rect 34744 5072 34794 5128
rect 34744 5070 34836 5072
rect 29269 5067 29335 5070
rect 30097 5067 30163 5070
rect 34789 5068 34836 5070
rect 34900 5068 34906 5132
rect 35566 5068 35572 5132
rect 35636 5130 35642 5132
rect 37733 5130 37799 5133
rect 39941 5130 40007 5133
rect 35636 5128 40007 5130
rect 35636 5072 37738 5128
rect 37794 5072 39946 5128
rect 40002 5072 40007 5128
rect 35636 5070 40007 5072
rect 35636 5068 35642 5070
rect 34789 5067 34855 5068
rect 37733 5067 37799 5070
rect 39941 5067 40007 5070
rect 40350 5068 40356 5132
rect 40420 5130 40426 5132
rect 40493 5130 40559 5133
rect 40420 5128 40559 5130
rect 40420 5072 40498 5128
rect 40554 5072 40559 5128
rect 40420 5070 40559 5072
rect 40420 5068 40426 5070
rect 40493 5067 40559 5070
rect 7833 4994 7899 4997
rect 18137 4994 18203 4997
rect 7833 4992 18203 4994
rect 7833 4936 7838 4992
rect 7894 4936 18142 4992
rect 18198 4936 18203 4992
rect 7833 4934 18203 4936
rect 7833 4931 7899 4934
rect 18137 4931 18203 4934
rect 24301 4994 24367 4997
rect 27613 4994 27679 4997
rect 24301 4992 27679 4994
rect 24301 4936 24306 4992
rect 24362 4936 27618 4992
rect 27674 4936 27679 4992
rect 24301 4934 27679 4936
rect 24301 4931 24367 4934
rect 27613 4931 27679 4934
rect 28901 4994 28967 4997
rect 34697 4994 34763 4997
rect 28901 4992 34763 4994
rect 28901 4936 28906 4992
rect 28962 4936 34702 4992
rect 34758 4936 34763 4992
rect 28901 4934 34763 4936
rect 28901 4931 28967 4934
rect 34697 4931 34763 4934
rect 5130 4928 5446 4929
rect 5130 4864 5136 4928
rect 5200 4864 5216 4928
rect 5280 4864 5296 4928
rect 5360 4864 5376 4928
rect 5440 4864 5446 4928
rect 5130 4863 5446 4864
rect 35850 4928 36166 4929
rect 35850 4864 35856 4928
rect 35920 4864 35936 4928
rect 36000 4864 36016 4928
rect 36080 4864 36096 4928
rect 36160 4864 36166 4928
rect 35850 4863 36166 4864
rect 66570 4928 66886 4929
rect 66570 4864 66576 4928
rect 66640 4864 66656 4928
rect 66720 4864 66736 4928
rect 66800 4864 66816 4928
rect 66880 4864 66886 4928
rect 66570 4863 66886 4864
rect 17861 4858 17927 4861
rect 21265 4858 21331 4861
rect 17861 4856 21331 4858
rect 17861 4800 17866 4856
rect 17922 4800 21270 4856
rect 21326 4800 21331 4856
rect 17861 4798 21331 4800
rect 17861 4795 17927 4798
rect 21265 4795 21331 4798
rect 23565 4858 23631 4861
rect 30966 4858 30972 4860
rect 23565 4856 30972 4858
rect 23565 4800 23570 4856
rect 23626 4800 30972 4856
rect 23565 4798 30972 4800
rect 23565 4795 23631 4798
rect 30966 4796 30972 4798
rect 31036 4796 31042 4860
rect 36445 4858 36511 4861
rect 37733 4858 37799 4861
rect 38193 4858 38259 4861
rect 36445 4856 38259 4858
rect 36445 4800 36450 4856
rect 36506 4800 37738 4856
rect 37794 4800 38198 4856
rect 38254 4800 38259 4856
rect 36445 4798 38259 4800
rect 36445 4795 36511 4798
rect 37733 4795 37799 4798
rect 38193 4795 38259 4798
rect 10593 4722 10659 4725
rect 10726 4722 10732 4724
rect 10593 4720 10732 4722
rect 10593 4664 10598 4720
rect 10654 4664 10732 4720
rect 10593 4662 10732 4664
rect 10593 4659 10659 4662
rect 10726 4660 10732 4662
rect 10796 4660 10802 4724
rect 11329 4722 11395 4725
rect 11462 4722 11468 4724
rect 11329 4720 11468 4722
rect 11329 4664 11334 4720
rect 11390 4664 11468 4720
rect 11329 4662 11468 4664
rect 11329 4659 11395 4662
rect 11462 4660 11468 4662
rect 11532 4660 11538 4724
rect 11973 4722 12039 4725
rect 12198 4722 12204 4724
rect 11973 4720 12204 4722
rect 11973 4664 11978 4720
rect 12034 4664 12204 4720
rect 11973 4662 12204 4664
rect 11973 4659 12039 4662
rect 12198 4660 12204 4662
rect 12268 4660 12274 4724
rect 13537 4722 13603 4725
rect 13670 4722 13676 4724
rect 13537 4720 13676 4722
rect 13537 4664 13542 4720
rect 13598 4664 13676 4720
rect 13537 4662 13676 4664
rect 13537 4659 13603 4662
rect 13670 4660 13676 4662
rect 13740 4660 13746 4724
rect 16481 4722 16547 4725
rect 17585 4722 17651 4725
rect 16481 4720 17651 4722
rect 16481 4664 16486 4720
rect 16542 4664 17590 4720
rect 17646 4664 17651 4720
rect 16481 4662 17651 4664
rect 16481 4659 16547 4662
rect 17585 4659 17651 4662
rect 17769 4722 17835 4725
rect 18137 4722 18203 4725
rect 23422 4722 23428 4724
rect 17769 4720 17970 4722
rect 17769 4664 17774 4720
rect 17830 4664 17970 4720
rect 17769 4662 17970 4664
rect 17769 4659 17835 4662
rect 15009 4450 15075 4453
rect 17677 4450 17743 4453
rect 15009 4448 17743 4450
rect 15009 4392 15014 4448
rect 15070 4392 17682 4448
rect 17738 4392 17743 4448
rect 15009 4390 17743 4392
rect 15009 4387 15075 4390
rect 17677 4387 17743 4390
rect 5790 4384 6106 4385
rect 5790 4320 5796 4384
rect 5860 4320 5876 4384
rect 5940 4320 5956 4384
rect 6020 4320 6036 4384
rect 6100 4320 6106 4384
rect 5790 4319 6106 4320
rect 12249 4314 12315 4317
rect 16389 4314 16455 4317
rect 12249 4312 16455 4314
rect 12249 4256 12254 4312
rect 12310 4256 16394 4312
rect 16450 4256 16455 4312
rect 12249 4254 16455 4256
rect 12249 4251 12315 4254
rect 16389 4251 16455 4254
rect 17534 4252 17540 4316
rect 17604 4314 17610 4316
rect 17604 4254 17786 4314
rect 17604 4252 17610 4254
rect 17726 4181 17786 4254
rect 11973 4178 12039 4181
rect 14733 4178 14799 4181
rect 11973 4176 14799 4178
rect 11973 4120 11978 4176
rect 12034 4120 14738 4176
rect 14794 4120 14799 4176
rect 11973 4118 14799 4120
rect 11973 4115 12039 4118
rect 14733 4115 14799 4118
rect 17309 4178 17375 4181
rect 17309 4176 17602 4178
rect 17309 4120 17314 4176
rect 17370 4120 17602 4176
rect 17309 4118 17602 4120
rect 17726 4176 17835 4181
rect 17726 4120 17774 4176
rect 17830 4120 17835 4176
rect 17726 4118 17835 4120
rect 17910 4178 17970 4662
rect 18137 4720 23428 4722
rect 18137 4664 18142 4720
rect 18198 4664 23428 4720
rect 18137 4662 23428 4664
rect 18137 4659 18203 4662
rect 23422 4660 23428 4662
rect 23492 4660 23498 4724
rect 26417 4722 26483 4725
rect 40125 4722 40191 4725
rect 26417 4720 40191 4722
rect 26417 4664 26422 4720
rect 26478 4664 40130 4720
rect 40186 4664 40191 4720
rect 26417 4662 40191 4664
rect 26417 4659 26483 4662
rect 40125 4659 40191 4662
rect 21725 4586 21791 4589
rect 24301 4586 24367 4589
rect 27981 4588 28047 4589
rect 28993 4588 29059 4589
rect 27981 4586 28028 4588
rect 21725 4584 24367 4586
rect 21725 4528 21730 4584
rect 21786 4528 24306 4584
rect 24362 4528 24367 4584
rect 21725 4526 24367 4528
rect 27936 4584 28028 4586
rect 27936 4528 27986 4584
rect 27936 4526 28028 4528
rect 21725 4523 21791 4526
rect 24301 4523 24367 4526
rect 27981 4524 28028 4526
rect 28092 4524 28098 4588
rect 28942 4586 28948 4588
rect 28902 4526 28948 4586
rect 29012 4584 29059 4588
rect 29054 4528 29059 4584
rect 28942 4524 28948 4526
rect 29012 4524 29059 4528
rect 27981 4523 28047 4524
rect 28993 4523 29059 4524
rect 29637 4586 29703 4589
rect 33133 4586 33199 4589
rect 29637 4584 33199 4586
rect 29637 4528 29642 4584
rect 29698 4528 33138 4584
rect 33194 4528 33199 4584
rect 29637 4526 33199 4528
rect 29637 4523 29703 4526
rect 33133 4523 33199 4526
rect 34973 4586 35039 4589
rect 42701 4586 42767 4589
rect 34973 4584 42767 4586
rect 34973 4528 34978 4584
rect 35034 4528 42706 4584
rect 42762 4528 42767 4584
rect 34973 4526 42767 4528
rect 34973 4523 35039 4526
rect 42701 4523 42767 4526
rect 20897 4450 20963 4453
rect 25865 4450 25931 4453
rect 20897 4448 25931 4450
rect 20897 4392 20902 4448
rect 20958 4392 25870 4448
rect 25926 4392 25931 4448
rect 20897 4390 25931 4392
rect 20897 4387 20963 4390
rect 25865 4387 25931 4390
rect 26918 4388 26924 4452
rect 26988 4450 26994 4452
rect 35566 4450 35572 4452
rect 26988 4390 35572 4450
rect 26988 4388 26994 4390
rect 35566 4388 35572 4390
rect 35636 4388 35642 4452
rect 39941 4450 40007 4453
rect 42701 4450 42767 4453
rect 39941 4448 42767 4450
rect 39941 4392 39946 4448
rect 40002 4392 42706 4448
rect 42762 4392 42767 4448
rect 39941 4390 42767 4392
rect 39941 4387 40007 4390
rect 42701 4387 42767 4390
rect 36510 4384 36826 4385
rect 36510 4320 36516 4384
rect 36580 4320 36596 4384
rect 36660 4320 36676 4384
rect 36740 4320 36756 4384
rect 36820 4320 36826 4384
rect 36510 4319 36826 4320
rect 67230 4384 67546 4385
rect 67230 4320 67236 4384
rect 67300 4320 67316 4384
rect 67380 4320 67396 4384
rect 67460 4320 67476 4384
rect 67540 4320 67546 4384
rect 67230 4319 67546 4320
rect 19977 4314 20043 4317
rect 22185 4314 22251 4317
rect 23197 4314 23263 4317
rect 25589 4314 25655 4317
rect 19977 4312 25655 4314
rect 19977 4256 19982 4312
rect 20038 4256 22190 4312
rect 22246 4256 23202 4312
rect 23258 4256 25594 4312
rect 25650 4256 25655 4312
rect 19977 4254 25655 4256
rect 19977 4251 20043 4254
rect 22185 4251 22251 4254
rect 23197 4251 23263 4254
rect 25589 4251 25655 4254
rect 27337 4314 27403 4317
rect 34697 4314 34763 4317
rect 27337 4312 34763 4314
rect 27337 4256 27342 4312
rect 27398 4256 34702 4312
rect 34758 4256 34763 4312
rect 27337 4254 34763 4256
rect 27337 4251 27403 4254
rect 34697 4251 34763 4254
rect 40769 4314 40835 4317
rect 42885 4314 42951 4317
rect 40769 4312 42951 4314
rect 40769 4256 40774 4312
rect 40830 4256 42890 4312
rect 42946 4256 42951 4312
rect 40769 4254 42951 4256
rect 40769 4251 40835 4254
rect 42885 4251 42951 4254
rect 24577 4178 24643 4181
rect 17910 4176 24643 4178
rect 17910 4120 24582 4176
rect 24638 4120 24643 4176
rect 17910 4118 24643 4120
rect 17309 4115 17375 4118
rect 17542 4045 17602 4118
rect 17769 4115 17835 4118
rect 24577 4115 24643 4118
rect 24894 4116 24900 4180
rect 24964 4178 24970 4180
rect 29637 4178 29703 4181
rect 24964 4176 29703 4178
rect 24964 4120 29642 4176
rect 29698 4120 29703 4176
rect 24964 4118 29703 4120
rect 24964 4116 24970 4118
rect 29637 4115 29703 4118
rect 36261 4178 36327 4181
rect 43897 4178 43963 4181
rect 36261 4176 43963 4178
rect 36261 4120 36266 4176
rect 36322 4120 43902 4176
rect 43958 4120 43963 4176
rect 36261 4118 43963 4120
rect 36261 4115 36327 4118
rect 43897 4115 43963 4118
rect 10041 4042 10107 4045
rect 16757 4044 16823 4045
rect 10174 4042 10180 4044
rect 10041 4040 10180 4042
rect 10041 3984 10046 4040
rect 10102 3984 10180 4040
rect 10041 3982 10180 3984
rect 10041 3979 10107 3982
rect 10174 3980 10180 3982
rect 10244 3980 10250 4044
rect 16757 4042 16804 4044
rect 16712 4040 16804 4042
rect 16712 3984 16762 4040
rect 16712 3982 16804 3984
rect 16757 3980 16804 3982
rect 16868 3980 16874 4044
rect 17542 4040 17651 4045
rect 17542 3984 17590 4040
rect 17646 3984 17651 4040
rect 17542 3982 17651 3984
rect 16757 3979 16823 3980
rect 17585 3979 17651 3982
rect 19885 4042 19951 4045
rect 21357 4044 21423 4045
rect 20662 4042 20668 4044
rect 19885 4040 20668 4042
rect 19885 3984 19890 4040
rect 19946 3984 20668 4040
rect 19885 3982 20668 3984
rect 19885 3979 19951 3982
rect 20662 3980 20668 3982
rect 20732 3980 20738 4044
rect 21357 4042 21404 4044
rect 21312 4040 21404 4042
rect 21312 3984 21362 4040
rect 21312 3982 21404 3984
rect 21357 3980 21404 3982
rect 21468 3980 21474 4044
rect 37549 4042 37615 4045
rect 37733 4042 37799 4045
rect 44725 4042 44791 4045
rect 22050 4040 37658 4042
rect 22050 3984 37554 4040
rect 37610 3984 37658 4040
rect 22050 3982 37658 3984
rect 21357 3979 21423 3980
rect 9489 3906 9555 3909
rect 15377 3906 15443 3909
rect 9489 3904 15443 3906
rect 9489 3848 9494 3904
rect 9550 3848 15382 3904
rect 15438 3848 15443 3904
rect 9489 3846 15443 3848
rect 9489 3843 9555 3846
rect 15377 3843 15443 3846
rect 15745 3906 15811 3909
rect 15878 3906 15884 3908
rect 15745 3904 15884 3906
rect 15745 3848 15750 3904
rect 15806 3848 15884 3904
rect 15745 3846 15884 3848
rect 15745 3843 15811 3846
rect 15878 3844 15884 3846
rect 15948 3844 15954 3908
rect 17309 3906 17375 3909
rect 18137 3906 18203 3909
rect 17309 3904 18203 3906
rect 17309 3848 17314 3904
rect 17370 3848 18142 3904
rect 18198 3848 18203 3904
rect 17309 3846 18203 3848
rect 17309 3843 17375 3846
rect 18137 3843 18203 3846
rect 19517 3906 19583 3909
rect 21633 3906 21699 3909
rect 19517 3904 21699 3906
rect 19517 3848 19522 3904
rect 19578 3848 21638 3904
rect 21694 3848 21699 3904
rect 19517 3846 21699 3848
rect 19517 3843 19583 3846
rect 21633 3843 21699 3846
rect 5130 3840 5446 3841
rect 5130 3776 5136 3840
rect 5200 3776 5216 3840
rect 5280 3776 5296 3840
rect 5360 3776 5376 3840
rect 5440 3776 5446 3840
rect 5130 3775 5446 3776
rect 11513 3770 11579 3773
rect 11646 3770 11652 3772
rect 11513 3768 11652 3770
rect 11513 3712 11518 3768
rect 11574 3712 11652 3768
rect 11513 3710 11652 3712
rect 11513 3707 11579 3710
rect 11646 3708 11652 3710
rect 11716 3708 11722 3772
rect 12801 3770 12867 3773
rect 18270 3770 18276 3772
rect 12801 3768 18276 3770
rect 12801 3712 12806 3768
rect 12862 3712 18276 3768
rect 12801 3710 18276 3712
rect 12801 3707 12867 3710
rect 18270 3708 18276 3710
rect 18340 3708 18346 3772
rect 20253 3770 20319 3773
rect 20478 3770 20484 3772
rect 20253 3768 20484 3770
rect 20253 3712 20258 3768
rect 20314 3712 20484 3768
rect 20253 3710 20484 3712
rect 20253 3707 20319 3710
rect 20478 3708 20484 3710
rect 20548 3708 20554 3772
rect 14222 3572 14228 3636
rect 14292 3634 14298 3636
rect 14641 3634 14707 3637
rect 14292 3632 14707 3634
rect 14292 3576 14646 3632
rect 14702 3576 14707 3632
rect 14292 3574 14707 3576
rect 14292 3572 14298 3574
rect 14641 3571 14707 3574
rect 14958 3572 14964 3636
rect 15028 3634 15034 3636
rect 15101 3634 15167 3637
rect 15028 3632 15167 3634
rect 15028 3576 15106 3632
rect 15162 3576 15167 3632
rect 15028 3574 15167 3576
rect 15028 3572 15034 3574
rect 15101 3571 15167 3574
rect 16297 3634 16363 3637
rect 22050 3634 22110 3982
rect 37549 3979 37658 3982
rect 37733 4040 44791 4042
rect 37733 3984 37738 4040
rect 37794 3984 44730 4040
rect 44786 3984 44791 4040
rect 37733 3982 44791 3984
rect 37733 3979 37799 3982
rect 44725 3979 44791 3982
rect 24945 3906 25011 3909
rect 26141 3908 26207 3909
rect 26141 3906 26188 3908
rect 24945 3904 25882 3906
rect 24945 3848 24950 3904
rect 25006 3848 25882 3904
rect 24945 3846 25882 3848
rect 26096 3904 26188 3906
rect 26096 3848 26146 3904
rect 26096 3846 26188 3848
rect 24945 3843 25011 3846
rect 25589 3772 25655 3773
rect 25589 3770 25636 3772
rect 25544 3768 25636 3770
rect 25544 3712 25594 3768
rect 25544 3710 25636 3712
rect 25589 3708 25636 3710
rect 25700 3708 25706 3772
rect 25822 3770 25882 3846
rect 26141 3844 26188 3846
rect 26252 3844 26258 3908
rect 26325 3906 26391 3909
rect 30925 3906 30991 3909
rect 26325 3904 30991 3906
rect 26325 3848 26330 3904
rect 26386 3848 30930 3904
rect 30986 3848 30991 3904
rect 26325 3846 30991 3848
rect 37598 3906 37658 3979
rect 41781 3906 41847 3909
rect 48313 3906 48379 3909
rect 37598 3904 48379 3906
rect 37598 3848 41786 3904
rect 41842 3848 48318 3904
rect 48374 3848 48379 3904
rect 37598 3846 48379 3848
rect 26141 3843 26207 3844
rect 26325 3843 26391 3846
rect 30925 3843 30991 3846
rect 41781 3843 41847 3846
rect 48313 3843 48379 3846
rect 35850 3840 36166 3841
rect 35850 3776 35856 3840
rect 35920 3776 35936 3840
rect 36000 3776 36016 3840
rect 36080 3776 36096 3840
rect 36160 3776 36166 3840
rect 35850 3775 36166 3776
rect 66570 3840 66886 3841
rect 66570 3776 66576 3840
rect 66640 3776 66656 3840
rect 66720 3776 66736 3840
rect 66800 3776 66816 3840
rect 66880 3776 66886 3840
rect 66570 3775 66886 3776
rect 30925 3770 30991 3773
rect 31201 3770 31267 3773
rect 25822 3768 31267 3770
rect 25822 3712 30930 3768
rect 30986 3712 31206 3768
rect 31262 3712 31267 3768
rect 25822 3710 31267 3712
rect 25589 3707 25655 3708
rect 30925 3707 30991 3710
rect 31201 3707 31267 3710
rect 38469 3770 38535 3773
rect 41321 3770 41387 3773
rect 38469 3768 41387 3770
rect 38469 3712 38474 3768
rect 38530 3712 41326 3768
rect 41382 3712 41387 3768
rect 38469 3710 41387 3712
rect 38469 3707 38535 3710
rect 41321 3707 41387 3710
rect 16297 3632 22110 3634
rect 16297 3576 16302 3632
rect 16358 3576 22110 3632
rect 16297 3574 22110 3576
rect 24761 3634 24827 3637
rect 29453 3634 29519 3637
rect 24761 3632 29519 3634
rect 24761 3576 24766 3632
rect 24822 3576 29458 3632
rect 29514 3576 29519 3632
rect 24761 3574 29519 3576
rect 16297 3571 16363 3574
rect 24761 3571 24827 3574
rect 29453 3571 29519 3574
rect 34605 3634 34671 3637
rect 39941 3634 40007 3637
rect 34605 3632 40007 3634
rect 34605 3576 34610 3632
rect 34666 3576 39946 3632
rect 40002 3576 40007 3632
rect 34605 3574 40007 3576
rect 34605 3571 34671 3574
rect 39941 3571 40007 3574
rect 40493 3634 40559 3637
rect 43253 3634 43319 3637
rect 40493 3632 43319 3634
rect 40493 3576 40498 3632
rect 40554 3576 43258 3632
rect 43314 3576 43319 3632
rect 40493 3574 43319 3576
rect 40493 3571 40559 3574
rect 43253 3571 43319 3574
rect 10961 3498 11027 3501
rect 26141 3498 26207 3501
rect 10961 3496 26207 3498
rect 10961 3440 10966 3496
rect 11022 3440 26146 3496
rect 26202 3440 26207 3496
rect 10961 3438 26207 3440
rect 10961 3435 11027 3438
rect 26141 3435 26207 3438
rect 28717 3498 28783 3501
rect 28717 3496 41430 3498
rect 28717 3440 28722 3496
rect 28778 3440 41430 3496
rect 28717 3438 41430 3440
rect 28717 3435 28783 3438
rect 11237 3362 11303 3365
rect 12341 3362 12407 3365
rect 11237 3360 12407 3362
rect 11237 3304 11242 3360
rect 11298 3304 12346 3360
rect 12402 3304 12407 3360
rect 11237 3302 12407 3304
rect 11237 3299 11303 3302
rect 12341 3299 12407 3302
rect 17166 3300 17172 3364
rect 17236 3362 17242 3364
rect 17309 3362 17375 3365
rect 17236 3360 17375 3362
rect 17236 3304 17314 3360
rect 17370 3304 17375 3360
rect 17236 3302 17375 3304
rect 17236 3300 17242 3302
rect 17309 3299 17375 3302
rect 17677 3362 17743 3365
rect 25681 3362 25747 3365
rect 26969 3364 27035 3365
rect 17677 3360 25747 3362
rect 17677 3304 17682 3360
rect 17738 3304 25686 3360
rect 25742 3304 25747 3360
rect 17677 3302 25747 3304
rect 17677 3299 17743 3302
rect 25681 3299 25747 3302
rect 26918 3300 26924 3364
rect 26988 3362 27035 3364
rect 29913 3362 29979 3365
rect 32806 3362 32812 3364
rect 26988 3360 27080 3362
rect 27030 3304 27080 3360
rect 26988 3302 27080 3304
rect 29913 3360 32812 3362
rect 29913 3304 29918 3360
rect 29974 3304 32812 3360
rect 29913 3302 32812 3304
rect 26988 3300 27035 3302
rect 26969 3299 27035 3300
rect 29913 3299 29979 3302
rect 32806 3300 32812 3302
rect 32876 3300 32882 3364
rect 33869 3362 33935 3365
rect 35198 3362 35204 3364
rect 33869 3360 35204 3362
rect 33869 3304 33874 3360
rect 33930 3304 35204 3360
rect 33869 3302 35204 3304
rect 33869 3299 33935 3302
rect 35198 3300 35204 3302
rect 35268 3300 35274 3364
rect 41370 3362 41430 3438
rect 42517 3362 42583 3365
rect 44173 3362 44239 3365
rect 41370 3360 44239 3362
rect 41370 3304 42522 3360
rect 42578 3304 44178 3360
rect 44234 3304 44239 3360
rect 41370 3302 44239 3304
rect 42517 3299 42583 3302
rect 44173 3299 44239 3302
rect 5790 3296 6106 3297
rect 5790 3232 5796 3296
rect 5860 3232 5876 3296
rect 5940 3232 5956 3296
rect 6020 3232 6036 3296
rect 6100 3232 6106 3296
rect 5790 3231 6106 3232
rect 36510 3296 36826 3297
rect 36510 3232 36516 3296
rect 36580 3232 36596 3296
rect 36660 3232 36676 3296
rect 36740 3232 36756 3296
rect 36820 3232 36826 3296
rect 36510 3231 36826 3232
rect 67230 3296 67546 3297
rect 67230 3232 67236 3296
rect 67300 3232 67316 3296
rect 67380 3232 67396 3296
rect 67460 3232 67476 3296
rect 67540 3232 67546 3296
rect 67230 3231 67546 3232
rect 8201 3228 8267 3229
rect 8150 3164 8156 3228
rect 8220 3226 8267 3228
rect 12617 3226 12683 3229
rect 20161 3226 20227 3229
rect 28717 3226 28783 3229
rect 8220 3224 8312 3226
rect 8262 3168 8312 3224
rect 8220 3166 8312 3168
rect 12617 3224 28783 3226
rect 12617 3168 12622 3224
rect 12678 3168 20166 3224
rect 20222 3168 28722 3224
rect 28778 3168 28783 3224
rect 12617 3166 28783 3168
rect 8220 3164 8267 3166
rect 8201 3163 8267 3164
rect 12617 3163 12683 3166
rect 20161 3163 20227 3166
rect 28717 3163 28783 3166
rect 28901 3226 28967 3229
rect 33358 3226 33364 3228
rect 28901 3224 33364 3226
rect 28901 3168 28906 3224
rect 28962 3168 33364 3224
rect 28901 3166 33364 3168
rect 28901 3163 28967 3166
rect 33358 3164 33364 3166
rect 33428 3164 33434 3228
rect 9949 3092 10015 3093
rect 9949 3090 9996 3092
rect 9904 3088 9996 3090
rect 9904 3032 9954 3088
rect 9904 3030 9996 3032
rect 9949 3028 9996 3030
rect 10060 3028 10066 3092
rect 13813 3090 13879 3093
rect 15101 3090 15167 3093
rect 17309 3090 17375 3093
rect 37406 3090 37412 3092
rect 13813 3088 17375 3090
rect 13813 3032 13818 3088
rect 13874 3032 15106 3088
rect 15162 3032 17314 3088
rect 17370 3032 17375 3088
rect 13813 3030 17375 3032
rect 9949 3027 10015 3028
rect 13813 3027 13879 3030
rect 15101 3027 15167 3030
rect 17309 3027 17375 3030
rect 22050 3030 37412 3090
rect 17493 2818 17559 2821
rect 22050 2818 22110 3030
rect 37406 3028 37412 3030
rect 37476 3028 37482 3092
rect 27102 2892 27108 2956
rect 27172 2954 27178 2956
rect 27337 2954 27403 2957
rect 27172 2952 27403 2954
rect 27172 2896 27342 2952
rect 27398 2896 27403 2952
rect 27172 2894 27403 2896
rect 27172 2892 27178 2894
rect 27337 2891 27403 2894
rect 28533 2952 28599 2957
rect 28533 2896 28538 2952
rect 28594 2896 28599 2952
rect 28533 2891 28599 2896
rect 30741 2954 30807 2957
rect 32765 2954 32831 2957
rect 33041 2956 33107 2957
rect 30741 2952 32831 2954
rect 30741 2896 30746 2952
rect 30802 2896 32770 2952
rect 32826 2896 32831 2952
rect 30741 2894 32831 2896
rect 30741 2891 30807 2894
rect 32765 2891 32831 2894
rect 32990 2892 32996 2956
rect 33060 2954 33107 2956
rect 39849 2954 39915 2957
rect 33060 2952 33152 2954
rect 33102 2896 33152 2952
rect 33060 2894 33152 2896
rect 35574 2952 39915 2954
rect 35574 2896 39854 2952
rect 39910 2896 39915 2952
rect 35574 2894 39915 2896
rect 33060 2892 33107 2894
rect 33041 2891 33107 2892
rect 28536 2818 28596 2891
rect 17493 2816 22110 2818
rect 17493 2760 17498 2816
rect 17554 2760 22110 2816
rect 17493 2758 22110 2760
rect 22372 2758 28596 2818
rect 31385 2818 31451 2821
rect 35574 2818 35634 2894
rect 39849 2891 39915 2894
rect 31385 2816 35634 2818
rect 31385 2760 31390 2816
rect 31446 2760 35634 2816
rect 31385 2758 35634 2760
rect 17493 2755 17559 2758
rect 5130 2752 5446 2753
rect 5130 2688 5136 2752
rect 5200 2688 5216 2752
rect 5280 2688 5296 2752
rect 5360 2688 5376 2752
rect 5440 2688 5446 2752
rect 5130 2687 5446 2688
rect 6545 2682 6611 2685
rect 15142 2682 15148 2684
rect 6545 2680 15148 2682
rect 6545 2624 6550 2680
rect 6606 2624 15148 2680
rect 6545 2622 15148 2624
rect 6545 2619 6611 2622
rect 15142 2620 15148 2622
rect 15212 2620 15218 2684
rect 20713 2682 20779 2685
rect 22372 2682 22432 2758
rect 31385 2755 31451 2758
rect 35850 2752 36166 2753
rect 35850 2688 35856 2752
rect 35920 2688 35936 2752
rect 36000 2688 36016 2752
rect 36080 2688 36096 2752
rect 36160 2688 36166 2752
rect 35850 2687 36166 2688
rect 66570 2752 66886 2753
rect 66570 2688 66576 2752
rect 66640 2688 66656 2752
rect 66720 2688 66736 2752
rect 66800 2688 66816 2752
rect 66880 2688 66886 2752
rect 66570 2687 66886 2688
rect 20713 2680 22432 2682
rect 20713 2624 20718 2680
rect 20774 2624 22432 2680
rect 20713 2622 22432 2624
rect 20713 2619 20779 2622
rect 22502 2620 22508 2684
rect 22572 2682 22578 2684
rect 22921 2682 22987 2685
rect 22572 2680 22987 2682
rect 22572 2624 22926 2680
rect 22982 2624 22987 2680
rect 22572 2622 22987 2624
rect 22572 2620 22578 2622
rect 22921 2619 22987 2622
rect 5625 2546 5691 2549
rect 19742 2546 19748 2548
rect 5625 2544 19748 2546
rect 5625 2488 5630 2544
rect 5686 2488 19748 2544
rect 5625 2486 19748 2488
rect 5625 2483 5691 2486
rect 19742 2484 19748 2486
rect 19812 2484 19818 2548
rect 22001 2546 22067 2549
rect 37222 2546 37228 2548
rect 22001 2544 37228 2546
rect 22001 2488 22006 2544
rect 22062 2488 37228 2544
rect 22001 2486 37228 2488
rect 22001 2483 22067 2486
rect 37222 2484 37228 2486
rect 37292 2484 37298 2548
rect 4889 2410 4955 2413
rect 19558 2410 19564 2412
rect 4889 2408 19564 2410
rect 4889 2352 4894 2408
rect 4950 2352 19564 2408
rect 4889 2350 19564 2352
rect 4889 2347 4955 2350
rect 19558 2348 19564 2350
rect 19628 2348 19634 2412
rect 28257 2410 28323 2413
rect 36302 2410 36308 2412
rect 28257 2408 36308 2410
rect 28257 2352 28262 2408
rect 28318 2352 36308 2408
rect 28257 2350 36308 2352
rect 28257 2347 28323 2350
rect 36302 2348 36308 2350
rect 36372 2348 36378 2412
rect 10593 2274 10659 2277
rect 18086 2274 18092 2276
rect 10593 2272 18092 2274
rect 10593 2216 10598 2272
rect 10654 2216 18092 2272
rect 10593 2214 18092 2216
rect 10593 2211 10659 2214
rect 18086 2212 18092 2214
rect 18156 2212 18162 2276
rect 21081 2274 21147 2277
rect 29678 2274 29684 2276
rect 21081 2272 29684 2274
rect 21081 2216 21086 2272
rect 21142 2216 29684 2272
rect 21081 2214 29684 2216
rect 21081 2211 21147 2214
rect 29678 2212 29684 2214
rect 29748 2212 29754 2276
rect 5790 2208 6106 2209
rect 5790 2144 5796 2208
rect 5860 2144 5876 2208
rect 5940 2144 5956 2208
rect 6020 2144 6036 2208
rect 6100 2144 6106 2208
rect 5790 2143 6106 2144
rect 36510 2208 36826 2209
rect 36510 2144 36516 2208
rect 36580 2144 36596 2208
rect 36660 2144 36676 2208
rect 36740 2144 36756 2208
rect 36820 2144 36826 2208
rect 36510 2143 36826 2144
rect 67230 2208 67546 2209
rect 67230 2144 67236 2208
rect 67300 2144 67316 2208
rect 67380 2144 67396 2208
rect 67460 2144 67476 2208
rect 67540 2144 67546 2208
rect 67230 2143 67546 2144
rect 17309 2138 17375 2141
rect 24894 2138 24900 2140
rect 17309 2136 24900 2138
rect 17309 2080 17314 2136
rect 17370 2080 24900 2136
rect 17309 2078 24900 2080
rect 17309 2075 17375 2078
rect 24894 2076 24900 2078
rect 24964 2076 24970 2140
rect 34278 2138 34284 2140
rect 31710 2078 34284 2138
rect 9029 2002 9095 2005
rect 18689 2002 18755 2005
rect 9029 2000 18755 2002
rect 9029 1944 9034 2000
rect 9090 1944 18694 2000
rect 18750 1944 18755 2000
rect 9029 1942 18755 1944
rect 9029 1939 9095 1942
rect 18689 1939 18755 1942
rect 22829 2002 22895 2005
rect 31710 2002 31770 2078
rect 34278 2076 34284 2078
rect 34348 2076 34354 2140
rect 22829 2000 31770 2002
rect 22829 1944 22834 2000
rect 22890 1944 31770 2000
rect 22829 1942 31770 1944
rect 22829 1939 22895 1942
rect 18270 1804 18276 1868
rect 18340 1866 18346 1868
rect 74257 1866 74323 1869
rect 18340 1864 74323 1866
rect 18340 1808 74262 1864
rect 74318 1808 74323 1864
rect 18340 1806 74323 1808
rect 18340 1804 18346 1806
rect 74257 1803 74323 1806
rect 27705 1594 27771 1597
rect 30782 1594 30788 1596
rect 27705 1592 30788 1594
rect 27705 1536 27710 1592
rect 27766 1536 30788 1592
rect 27705 1534 30788 1536
rect 27705 1531 27771 1534
rect 30782 1532 30788 1534
rect 30852 1532 30858 1596
rect 28349 1458 28415 1461
rect 29361 1458 29427 1461
rect 28349 1456 29427 1458
rect 28349 1400 28354 1456
rect 28410 1400 29366 1456
rect 29422 1400 29427 1456
rect 28349 1398 29427 1400
rect 28349 1395 28415 1398
rect 29361 1395 29427 1398
rect 36721 1458 36787 1461
rect 37641 1458 37707 1461
rect 36721 1456 37707 1458
rect 36721 1400 36726 1456
rect 36782 1400 37646 1456
rect 37702 1400 37707 1456
rect 36721 1398 37707 1400
rect 36721 1395 36787 1398
rect 37641 1395 37707 1398
rect 6729 1322 6795 1325
rect 10961 1322 11027 1325
rect 6729 1320 11027 1322
rect 6729 1264 6734 1320
rect 6790 1264 10966 1320
rect 11022 1264 11027 1320
rect 6729 1262 11027 1264
rect 6729 1259 6795 1262
rect 10961 1259 11027 1262
rect 31518 1260 31524 1324
rect 31588 1322 31594 1324
rect 35433 1322 35499 1325
rect 31588 1320 35499 1322
rect 31588 1264 35438 1320
rect 35494 1264 35499 1320
rect 31588 1262 35499 1264
rect 31588 1260 31594 1262
rect 35433 1259 35499 1262
rect 14774 172 14780 236
rect 14844 234 14850 236
rect 25037 234 25103 237
rect 14844 232 25103 234
rect 14844 176 25042 232
rect 25098 176 25103 232
rect 14844 174 25103 176
rect 14844 172 14850 174
rect 25037 171 25103 174
rect 9121 98 9187 101
rect 28942 98 28948 100
rect 9121 96 28948 98
rect 9121 40 9126 96
rect 9182 40 28948 96
rect 9121 38 28948 40
rect 9121 35 9187 38
rect 28942 36 28948 38
rect 29012 36 29018 100
<< via3 >>
rect 5136 37564 5200 37568
rect 5136 37508 5140 37564
rect 5140 37508 5196 37564
rect 5196 37508 5200 37564
rect 5136 37504 5200 37508
rect 5216 37564 5280 37568
rect 5216 37508 5220 37564
rect 5220 37508 5276 37564
rect 5276 37508 5280 37564
rect 5216 37504 5280 37508
rect 5296 37564 5360 37568
rect 5296 37508 5300 37564
rect 5300 37508 5356 37564
rect 5356 37508 5360 37564
rect 5296 37504 5360 37508
rect 5376 37564 5440 37568
rect 5376 37508 5380 37564
rect 5380 37508 5436 37564
rect 5436 37508 5440 37564
rect 5376 37504 5440 37508
rect 35856 37564 35920 37568
rect 35856 37508 35860 37564
rect 35860 37508 35916 37564
rect 35916 37508 35920 37564
rect 35856 37504 35920 37508
rect 35936 37564 36000 37568
rect 35936 37508 35940 37564
rect 35940 37508 35996 37564
rect 35996 37508 36000 37564
rect 35936 37504 36000 37508
rect 36016 37564 36080 37568
rect 36016 37508 36020 37564
rect 36020 37508 36076 37564
rect 36076 37508 36080 37564
rect 36016 37504 36080 37508
rect 36096 37564 36160 37568
rect 36096 37508 36100 37564
rect 36100 37508 36156 37564
rect 36156 37508 36160 37564
rect 36096 37504 36160 37508
rect 66576 37564 66640 37568
rect 66576 37508 66580 37564
rect 66580 37508 66636 37564
rect 66636 37508 66640 37564
rect 66576 37504 66640 37508
rect 66656 37564 66720 37568
rect 66656 37508 66660 37564
rect 66660 37508 66716 37564
rect 66716 37508 66720 37564
rect 66656 37504 66720 37508
rect 66736 37564 66800 37568
rect 66736 37508 66740 37564
rect 66740 37508 66796 37564
rect 66796 37508 66800 37564
rect 66736 37504 66800 37508
rect 66816 37564 66880 37568
rect 66816 37508 66820 37564
rect 66820 37508 66876 37564
rect 66876 37508 66880 37564
rect 66816 37504 66880 37508
rect 5796 37020 5860 37024
rect 5796 36964 5800 37020
rect 5800 36964 5856 37020
rect 5856 36964 5860 37020
rect 5796 36960 5860 36964
rect 5876 37020 5940 37024
rect 5876 36964 5880 37020
rect 5880 36964 5936 37020
rect 5936 36964 5940 37020
rect 5876 36960 5940 36964
rect 5956 37020 6020 37024
rect 5956 36964 5960 37020
rect 5960 36964 6016 37020
rect 6016 36964 6020 37020
rect 5956 36960 6020 36964
rect 6036 37020 6100 37024
rect 6036 36964 6040 37020
rect 6040 36964 6096 37020
rect 6096 36964 6100 37020
rect 6036 36960 6100 36964
rect 36516 37020 36580 37024
rect 36516 36964 36520 37020
rect 36520 36964 36576 37020
rect 36576 36964 36580 37020
rect 36516 36960 36580 36964
rect 36596 37020 36660 37024
rect 36596 36964 36600 37020
rect 36600 36964 36656 37020
rect 36656 36964 36660 37020
rect 36596 36960 36660 36964
rect 36676 37020 36740 37024
rect 36676 36964 36680 37020
rect 36680 36964 36736 37020
rect 36736 36964 36740 37020
rect 36676 36960 36740 36964
rect 36756 37020 36820 37024
rect 36756 36964 36760 37020
rect 36760 36964 36816 37020
rect 36816 36964 36820 37020
rect 36756 36960 36820 36964
rect 67236 37020 67300 37024
rect 67236 36964 67240 37020
rect 67240 36964 67296 37020
rect 67296 36964 67300 37020
rect 67236 36960 67300 36964
rect 67316 37020 67380 37024
rect 67316 36964 67320 37020
rect 67320 36964 67376 37020
rect 67376 36964 67380 37020
rect 67316 36960 67380 36964
rect 67396 37020 67460 37024
rect 67396 36964 67400 37020
rect 67400 36964 67456 37020
rect 67456 36964 67460 37020
rect 67396 36960 67460 36964
rect 67476 37020 67540 37024
rect 67476 36964 67480 37020
rect 67480 36964 67536 37020
rect 67536 36964 67540 37020
rect 67476 36960 67540 36964
rect 14596 36544 14660 36548
rect 14596 36488 14610 36544
rect 14610 36488 14660 36544
rect 14596 36484 14660 36488
rect 5136 36476 5200 36480
rect 5136 36420 5140 36476
rect 5140 36420 5196 36476
rect 5196 36420 5200 36476
rect 5136 36416 5200 36420
rect 5216 36476 5280 36480
rect 5216 36420 5220 36476
rect 5220 36420 5276 36476
rect 5276 36420 5280 36476
rect 5216 36416 5280 36420
rect 5296 36476 5360 36480
rect 5296 36420 5300 36476
rect 5300 36420 5356 36476
rect 5356 36420 5360 36476
rect 5296 36416 5360 36420
rect 5376 36476 5440 36480
rect 5376 36420 5380 36476
rect 5380 36420 5436 36476
rect 5436 36420 5440 36476
rect 5376 36416 5440 36420
rect 35856 36476 35920 36480
rect 35856 36420 35860 36476
rect 35860 36420 35916 36476
rect 35916 36420 35920 36476
rect 35856 36416 35920 36420
rect 35936 36476 36000 36480
rect 35936 36420 35940 36476
rect 35940 36420 35996 36476
rect 35996 36420 36000 36476
rect 35936 36416 36000 36420
rect 36016 36476 36080 36480
rect 36016 36420 36020 36476
rect 36020 36420 36076 36476
rect 36076 36420 36080 36476
rect 36016 36416 36080 36420
rect 36096 36476 36160 36480
rect 36096 36420 36100 36476
rect 36100 36420 36156 36476
rect 36156 36420 36160 36476
rect 36096 36416 36160 36420
rect 66576 36476 66640 36480
rect 66576 36420 66580 36476
rect 66580 36420 66636 36476
rect 66636 36420 66640 36476
rect 66576 36416 66640 36420
rect 66656 36476 66720 36480
rect 66656 36420 66660 36476
rect 66660 36420 66716 36476
rect 66716 36420 66720 36476
rect 66656 36416 66720 36420
rect 66736 36476 66800 36480
rect 66736 36420 66740 36476
rect 66740 36420 66796 36476
rect 66796 36420 66800 36476
rect 66736 36416 66800 36420
rect 66816 36476 66880 36480
rect 66816 36420 66820 36476
rect 66820 36420 66876 36476
rect 66876 36420 66880 36476
rect 66816 36416 66880 36420
rect 31524 36348 31588 36412
rect 5796 35932 5860 35936
rect 5796 35876 5800 35932
rect 5800 35876 5856 35932
rect 5856 35876 5860 35932
rect 5796 35872 5860 35876
rect 5876 35932 5940 35936
rect 5876 35876 5880 35932
rect 5880 35876 5936 35932
rect 5936 35876 5940 35932
rect 5876 35872 5940 35876
rect 5956 35932 6020 35936
rect 5956 35876 5960 35932
rect 5960 35876 6016 35932
rect 6016 35876 6020 35932
rect 5956 35872 6020 35876
rect 6036 35932 6100 35936
rect 6036 35876 6040 35932
rect 6040 35876 6096 35932
rect 6096 35876 6100 35932
rect 6036 35872 6100 35876
rect 36516 35932 36580 35936
rect 36516 35876 36520 35932
rect 36520 35876 36576 35932
rect 36576 35876 36580 35932
rect 36516 35872 36580 35876
rect 36596 35932 36660 35936
rect 36596 35876 36600 35932
rect 36600 35876 36656 35932
rect 36656 35876 36660 35932
rect 36596 35872 36660 35876
rect 36676 35932 36740 35936
rect 36676 35876 36680 35932
rect 36680 35876 36736 35932
rect 36736 35876 36740 35932
rect 36676 35872 36740 35876
rect 36756 35932 36820 35936
rect 36756 35876 36760 35932
rect 36760 35876 36816 35932
rect 36816 35876 36820 35932
rect 36756 35872 36820 35876
rect 67236 35932 67300 35936
rect 67236 35876 67240 35932
rect 67240 35876 67296 35932
rect 67296 35876 67300 35932
rect 67236 35872 67300 35876
rect 67316 35932 67380 35936
rect 67316 35876 67320 35932
rect 67320 35876 67376 35932
rect 67376 35876 67380 35932
rect 67316 35872 67380 35876
rect 67396 35932 67460 35936
rect 67396 35876 67400 35932
rect 67400 35876 67456 35932
rect 67456 35876 67460 35932
rect 67396 35872 67460 35876
rect 67476 35932 67540 35936
rect 67476 35876 67480 35932
rect 67480 35876 67536 35932
rect 67536 35876 67540 35932
rect 67476 35872 67540 35876
rect 5136 35388 5200 35392
rect 5136 35332 5140 35388
rect 5140 35332 5196 35388
rect 5196 35332 5200 35388
rect 5136 35328 5200 35332
rect 5216 35388 5280 35392
rect 5216 35332 5220 35388
rect 5220 35332 5276 35388
rect 5276 35332 5280 35388
rect 5216 35328 5280 35332
rect 5296 35388 5360 35392
rect 5296 35332 5300 35388
rect 5300 35332 5356 35388
rect 5356 35332 5360 35388
rect 5296 35328 5360 35332
rect 5376 35388 5440 35392
rect 5376 35332 5380 35388
rect 5380 35332 5436 35388
rect 5436 35332 5440 35388
rect 5376 35328 5440 35332
rect 35856 35388 35920 35392
rect 35856 35332 35860 35388
rect 35860 35332 35916 35388
rect 35916 35332 35920 35388
rect 35856 35328 35920 35332
rect 35936 35388 36000 35392
rect 35936 35332 35940 35388
rect 35940 35332 35996 35388
rect 35996 35332 36000 35388
rect 35936 35328 36000 35332
rect 36016 35388 36080 35392
rect 36016 35332 36020 35388
rect 36020 35332 36076 35388
rect 36076 35332 36080 35388
rect 36016 35328 36080 35332
rect 36096 35388 36160 35392
rect 36096 35332 36100 35388
rect 36100 35332 36156 35388
rect 36156 35332 36160 35388
rect 36096 35328 36160 35332
rect 66576 35388 66640 35392
rect 66576 35332 66580 35388
rect 66580 35332 66636 35388
rect 66636 35332 66640 35388
rect 66576 35328 66640 35332
rect 66656 35388 66720 35392
rect 66656 35332 66660 35388
rect 66660 35332 66716 35388
rect 66716 35332 66720 35388
rect 66656 35328 66720 35332
rect 66736 35388 66800 35392
rect 66736 35332 66740 35388
rect 66740 35332 66796 35388
rect 66796 35332 66800 35388
rect 66736 35328 66800 35332
rect 66816 35388 66880 35392
rect 66816 35332 66820 35388
rect 66820 35332 66876 35388
rect 66876 35332 66880 35388
rect 66816 35328 66880 35332
rect 5796 34844 5860 34848
rect 5796 34788 5800 34844
rect 5800 34788 5856 34844
rect 5856 34788 5860 34844
rect 5796 34784 5860 34788
rect 5876 34844 5940 34848
rect 5876 34788 5880 34844
rect 5880 34788 5936 34844
rect 5936 34788 5940 34844
rect 5876 34784 5940 34788
rect 5956 34844 6020 34848
rect 5956 34788 5960 34844
rect 5960 34788 6016 34844
rect 6016 34788 6020 34844
rect 5956 34784 6020 34788
rect 6036 34844 6100 34848
rect 6036 34788 6040 34844
rect 6040 34788 6096 34844
rect 6096 34788 6100 34844
rect 6036 34784 6100 34788
rect 36516 34844 36580 34848
rect 36516 34788 36520 34844
rect 36520 34788 36576 34844
rect 36576 34788 36580 34844
rect 36516 34784 36580 34788
rect 36596 34844 36660 34848
rect 36596 34788 36600 34844
rect 36600 34788 36656 34844
rect 36656 34788 36660 34844
rect 36596 34784 36660 34788
rect 36676 34844 36740 34848
rect 36676 34788 36680 34844
rect 36680 34788 36736 34844
rect 36736 34788 36740 34844
rect 36676 34784 36740 34788
rect 36756 34844 36820 34848
rect 36756 34788 36760 34844
rect 36760 34788 36816 34844
rect 36816 34788 36820 34844
rect 36756 34784 36820 34788
rect 67236 34844 67300 34848
rect 67236 34788 67240 34844
rect 67240 34788 67296 34844
rect 67296 34788 67300 34844
rect 67236 34784 67300 34788
rect 67316 34844 67380 34848
rect 67316 34788 67320 34844
rect 67320 34788 67376 34844
rect 67376 34788 67380 34844
rect 67316 34784 67380 34788
rect 67396 34844 67460 34848
rect 67396 34788 67400 34844
rect 67400 34788 67456 34844
rect 67456 34788 67460 34844
rect 67396 34784 67460 34788
rect 67476 34844 67540 34848
rect 67476 34788 67480 34844
rect 67480 34788 67536 34844
rect 67536 34788 67540 34844
rect 67476 34784 67540 34788
rect 5136 34300 5200 34304
rect 5136 34244 5140 34300
rect 5140 34244 5196 34300
rect 5196 34244 5200 34300
rect 5136 34240 5200 34244
rect 5216 34300 5280 34304
rect 5216 34244 5220 34300
rect 5220 34244 5276 34300
rect 5276 34244 5280 34300
rect 5216 34240 5280 34244
rect 5296 34300 5360 34304
rect 5296 34244 5300 34300
rect 5300 34244 5356 34300
rect 5356 34244 5360 34300
rect 5296 34240 5360 34244
rect 5376 34300 5440 34304
rect 5376 34244 5380 34300
rect 5380 34244 5436 34300
rect 5436 34244 5440 34300
rect 5376 34240 5440 34244
rect 35856 34300 35920 34304
rect 35856 34244 35860 34300
rect 35860 34244 35916 34300
rect 35916 34244 35920 34300
rect 35856 34240 35920 34244
rect 35936 34300 36000 34304
rect 35936 34244 35940 34300
rect 35940 34244 35996 34300
rect 35996 34244 36000 34300
rect 35936 34240 36000 34244
rect 36016 34300 36080 34304
rect 36016 34244 36020 34300
rect 36020 34244 36076 34300
rect 36076 34244 36080 34300
rect 36016 34240 36080 34244
rect 36096 34300 36160 34304
rect 36096 34244 36100 34300
rect 36100 34244 36156 34300
rect 36156 34244 36160 34300
rect 36096 34240 36160 34244
rect 66576 34300 66640 34304
rect 66576 34244 66580 34300
rect 66580 34244 66636 34300
rect 66636 34244 66640 34300
rect 66576 34240 66640 34244
rect 66656 34300 66720 34304
rect 66656 34244 66660 34300
rect 66660 34244 66716 34300
rect 66716 34244 66720 34300
rect 66656 34240 66720 34244
rect 66736 34300 66800 34304
rect 66736 34244 66740 34300
rect 66740 34244 66796 34300
rect 66796 34244 66800 34300
rect 66736 34240 66800 34244
rect 66816 34300 66880 34304
rect 66816 34244 66820 34300
rect 66820 34244 66876 34300
rect 66876 34244 66880 34300
rect 66816 34240 66880 34244
rect 5796 33756 5860 33760
rect 5796 33700 5800 33756
rect 5800 33700 5856 33756
rect 5856 33700 5860 33756
rect 5796 33696 5860 33700
rect 5876 33756 5940 33760
rect 5876 33700 5880 33756
rect 5880 33700 5936 33756
rect 5936 33700 5940 33756
rect 5876 33696 5940 33700
rect 5956 33756 6020 33760
rect 5956 33700 5960 33756
rect 5960 33700 6016 33756
rect 6016 33700 6020 33756
rect 5956 33696 6020 33700
rect 6036 33756 6100 33760
rect 6036 33700 6040 33756
rect 6040 33700 6096 33756
rect 6096 33700 6100 33756
rect 6036 33696 6100 33700
rect 36516 33756 36580 33760
rect 36516 33700 36520 33756
rect 36520 33700 36576 33756
rect 36576 33700 36580 33756
rect 36516 33696 36580 33700
rect 36596 33756 36660 33760
rect 36596 33700 36600 33756
rect 36600 33700 36656 33756
rect 36656 33700 36660 33756
rect 36596 33696 36660 33700
rect 36676 33756 36740 33760
rect 36676 33700 36680 33756
rect 36680 33700 36736 33756
rect 36736 33700 36740 33756
rect 36676 33696 36740 33700
rect 36756 33756 36820 33760
rect 36756 33700 36760 33756
rect 36760 33700 36816 33756
rect 36816 33700 36820 33756
rect 36756 33696 36820 33700
rect 67236 33756 67300 33760
rect 67236 33700 67240 33756
rect 67240 33700 67296 33756
rect 67296 33700 67300 33756
rect 67236 33696 67300 33700
rect 67316 33756 67380 33760
rect 67316 33700 67320 33756
rect 67320 33700 67376 33756
rect 67376 33700 67380 33756
rect 67316 33696 67380 33700
rect 67396 33756 67460 33760
rect 67396 33700 67400 33756
rect 67400 33700 67456 33756
rect 67456 33700 67460 33756
rect 67396 33696 67460 33700
rect 67476 33756 67540 33760
rect 67476 33700 67480 33756
rect 67480 33700 67536 33756
rect 67536 33700 67540 33756
rect 67476 33696 67540 33700
rect 5136 33212 5200 33216
rect 5136 33156 5140 33212
rect 5140 33156 5196 33212
rect 5196 33156 5200 33212
rect 5136 33152 5200 33156
rect 5216 33212 5280 33216
rect 5216 33156 5220 33212
rect 5220 33156 5276 33212
rect 5276 33156 5280 33212
rect 5216 33152 5280 33156
rect 5296 33212 5360 33216
rect 5296 33156 5300 33212
rect 5300 33156 5356 33212
rect 5356 33156 5360 33212
rect 5296 33152 5360 33156
rect 5376 33212 5440 33216
rect 5376 33156 5380 33212
rect 5380 33156 5436 33212
rect 5436 33156 5440 33212
rect 5376 33152 5440 33156
rect 35856 33212 35920 33216
rect 35856 33156 35860 33212
rect 35860 33156 35916 33212
rect 35916 33156 35920 33212
rect 35856 33152 35920 33156
rect 35936 33212 36000 33216
rect 35936 33156 35940 33212
rect 35940 33156 35996 33212
rect 35996 33156 36000 33212
rect 35936 33152 36000 33156
rect 36016 33212 36080 33216
rect 36016 33156 36020 33212
rect 36020 33156 36076 33212
rect 36076 33156 36080 33212
rect 36016 33152 36080 33156
rect 36096 33212 36160 33216
rect 36096 33156 36100 33212
rect 36100 33156 36156 33212
rect 36156 33156 36160 33212
rect 36096 33152 36160 33156
rect 66576 33212 66640 33216
rect 66576 33156 66580 33212
rect 66580 33156 66636 33212
rect 66636 33156 66640 33212
rect 66576 33152 66640 33156
rect 66656 33212 66720 33216
rect 66656 33156 66660 33212
rect 66660 33156 66716 33212
rect 66716 33156 66720 33212
rect 66656 33152 66720 33156
rect 66736 33212 66800 33216
rect 66736 33156 66740 33212
rect 66740 33156 66796 33212
rect 66796 33156 66800 33212
rect 66736 33152 66800 33156
rect 66816 33212 66880 33216
rect 66816 33156 66820 33212
rect 66820 33156 66876 33212
rect 66876 33156 66880 33212
rect 66816 33152 66880 33156
rect 5796 32668 5860 32672
rect 5796 32612 5800 32668
rect 5800 32612 5856 32668
rect 5856 32612 5860 32668
rect 5796 32608 5860 32612
rect 5876 32668 5940 32672
rect 5876 32612 5880 32668
rect 5880 32612 5936 32668
rect 5936 32612 5940 32668
rect 5876 32608 5940 32612
rect 5956 32668 6020 32672
rect 5956 32612 5960 32668
rect 5960 32612 6016 32668
rect 6016 32612 6020 32668
rect 5956 32608 6020 32612
rect 6036 32668 6100 32672
rect 6036 32612 6040 32668
rect 6040 32612 6096 32668
rect 6096 32612 6100 32668
rect 6036 32608 6100 32612
rect 36516 32668 36580 32672
rect 36516 32612 36520 32668
rect 36520 32612 36576 32668
rect 36576 32612 36580 32668
rect 36516 32608 36580 32612
rect 36596 32668 36660 32672
rect 36596 32612 36600 32668
rect 36600 32612 36656 32668
rect 36656 32612 36660 32668
rect 36596 32608 36660 32612
rect 36676 32668 36740 32672
rect 36676 32612 36680 32668
rect 36680 32612 36736 32668
rect 36736 32612 36740 32668
rect 36676 32608 36740 32612
rect 36756 32668 36820 32672
rect 36756 32612 36760 32668
rect 36760 32612 36816 32668
rect 36816 32612 36820 32668
rect 36756 32608 36820 32612
rect 67236 32668 67300 32672
rect 67236 32612 67240 32668
rect 67240 32612 67296 32668
rect 67296 32612 67300 32668
rect 67236 32608 67300 32612
rect 67316 32668 67380 32672
rect 67316 32612 67320 32668
rect 67320 32612 67376 32668
rect 67376 32612 67380 32668
rect 67316 32608 67380 32612
rect 67396 32668 67460 32672
rect 67396 32612 67400 32668
rect 67400 32612 67456 32668
rect 67456 32612 67460 32668
rect 67396 32608 67460 32612
rect 67476 32668 67540 32672
rect 67476 32612 67480 32668
rect 67480 32612 67536 32668
rect 67536 32612 67540 32668
rect 67476 32608 67540 32612
rect 33180 32404 33244 32468
rect 5136 32124 5200 32128
rect 5136 32068 5140 32124
rect 5140 32068 5196 32124
rect 5196 32068 5200 32124
rect 5136 32064 5200 32068
rect 5216 32124 5280 32128
rect 5216 32068 5220 32124
rect 5220 32068 5276 32124
rect 5276 32068 5280 32124
rect 5216 32064 5280 32068
rect 5296 32124 5360 32128
rect 5296 32068 5300 32124
rect 5300 32068 5356 32124
rect 5356 32068 5360 32124
rect 5296 32064 5360 32068
rect 5376 32124 5440 32128
rect 5376 32068 5380 32124
rect 5380 32068 5436 32124
rect 5436 32068 5440 32124
rect 5376 32064 5440 32068
rect 35856 32124 35920 32128
rect 35856 32068 35860 32124
rect 35860 32068 35916 32124
rect 35916 32068 35920 32124
rect 35856 32064 35920 32068
rect 35936 32124 36000 32128
rect 35936 32068 35940 32124
rect 35940 32068 35996 32124
rect 35996 32068 36000 32124
rect 35936 32064 36000 32068
rect 36016 32124 36080 32128
rect 36016 32068 36020 32124
rect 36020 32068 36076 32124
rect 36076 32068 36080 32124
rect 36016 32064 36080 32068
rect 36096 32124 36160 32128
rect 36096 32068 36100 32124
rect 36100 32068 36156 32124
rect 36156 32068 36160 32124
rect 36096 32064 36160 32068
rect 66576 32124 66640 32128
rect 66576 32068 66580 32124
rect 66580 32068 66636 32124
rect 66636 32068 66640 32124
rect 66576 32064 66640 32068
rect 66656 32124 66720 32128
rect 66656 32068 66660 32124
rect 66660 32068 66716 32124
rect 66716 32068 66720 32124
rect 66656 32064 66720 32068
rect 66736 32124 66800 32128
rect 66736 32068 66740 32124
rect 66740 32068 66796 32124
rect 66796 32068 66800 32124
rect 66736 32064 66800 32068
rect 66816 32124 66880 32128
rect 66816 32068 66820 32124
rect 66820 32068 66876 32124
rect 66876 32068 66880 32124
rect 66816 32064 66880 32068
rect 5796 31580 5860 31584
rect 5796 31524 5800 31580
rect 5800 31524 5856 31580
rect 5856 31524 5860 31580
rect 5796 31520 5860 31524
rect 5876 31580 5940 31584
rect 5876 31524 5880 31580
rect 5880 31524 5936 31580
rect 5936 31524 5940 31580
rect 5876 31520 5940 31524
rect 5956 31580 6020 31584
rect 5956 31524 5960 31580
rect 5960 31524 6016 31580
rect 6016 31524 6020 31580
rect 5956 31520 6020 31524
rect 6036 31580 6100 31584
rect 6036 31524 6040 31580
rect 6040 31524 6096 31580
rect 6096 31524 6100 31580
rect 6036 31520 6100 31524
rect 36516 31580 36580 31584
rect 36516 31524 36520 31580
rect 36520 31524 36576 31580
rect 36576 31524 36580 31580
rect 36516 31520 36580 31524
rect 36596 31580 36660 31584
rect 36596 31524 36600 31580
rect 36600 31524 36656 31580
rect 36656 31524 36660 31580
rect 36596 31520 36660 31524
rect 36676 31580 36740 31584
rect 36676 31524 36680 31580
rect 36680 31524 36736 31580
rect 36736 31524 36740 31580
rect 36676 31520 36740 31524
rect 36756 31580 36820 31584
rect 36756 31524 36760 31580
rect 36760 31524 36816 31580
rect 36816 31524 36820 31580
rect 36756 31520 36820 31524
rect 67236 31580 67300 31584
rect 67236 31524 67240 31580
rect 67240 31524 67296 31580
rect 67296 31524 67300 31580
rect 67236 31520 67300 31524
rect 67316 31580 67380 31584
rect 67316 31524 67320 31580
rect 67320 31524 67376 31580
rect 67376 31524 67380 31580
rect 67316 31520 67380 31524
rect 67396 31580 67460 31584
rect 67396 31524 67400 31580
rect 67400 31524 67456 31580
rect 67456 31524 67460 31580
rect 67396 31520 67460 31524
rect 67476 31580 67540 31584
rect 67476 31524 67480 31580
rect 67480 31524 67536 31580
rect 67536 31524 67540 31580
rect 67476 31520 67540 31524
rect 5136 31036 5200 31040
rect 5136 30980 5140 31036
rect 5140 30980 5196 31036
rect 5196 30980 5200 31036
rect 5136 30976 5200 30980
rect 5216 31036 5280 31040
rect 5216 30980 5220 31036
rect 5220 30980 5276 31036
rect 5276 30980 5280 31036
rect 5216 30976 5280 30980
rect 5296 31036 5360 31040
rect 5296 30980 5300 31036
rect 5300 30980 5356 31036
rect 5356 30980 5360 31036
rect 5296 30976 5360 30980
rect 5376 31036 5440 31040
rect 5376 30980 5380 31036
rect 5380 30980 5436 31036
rect 5436 30980 5440 31036
rect 5376 30976 5440 30980
rect 35856 31036 35920 31040
rect 35856 30980 35860 31036
rect 35860 30980 35916 31036
rect 35916 30980 35920 31036
rect 35856 30976 35920 30980
rect 35936 31036 36000 31040
rect 35936 30980 35940 31036
rect 35940 30980 35996 31036
rect 35996 30980 36000 31036
rect 35936 30976 36000 30980
rect 36016 31036 36080 31040
rect 36016 30980 36020 31036
rect 36020 30980 36076 31036
rect 36076 30980 36080 31036
rect 36016 30976 36080 30980
rect 36096 31036 36160 31040
rect 36096 30980 36100 31036
rect 36100 30980 36156 31036
rect 36156 30980 36160 31036
rect 36096 30976 36160 30980
rect 66576 31036 66640 31040
rect 66576 30980 66580 31036
rect 66580 30980 66636 31036
rect 66636 30980 66640 31036
rect 66576 30976 66640 30980
rect 66656 31036 66720 31040
rect 66656 30980 66660 31036
rect 66660 30980 66716 31036
rect 66716 30980 66720 31036
rect 66656 30976 66720 30980
rect 66736 31036 66800 31040
rect 66736 30980 66740 31036
rect 66740 30980 66796 31036
rect 66796 30980 66800 31036
rect 66736 30976 66800 30980
rect 66816 31036 66880 31040
rect 66816 30980 66820 31036
rect 66820 30980 66876 31036
rect 66876 30980 66880 31036
rect 66816 30976 66880 30980
rect 5796 30492 5860 30496
rect 5796 30436 5800 30492
rect 5800 30436 5856 30492
rect 5856 30436 5860 30492
rect 5796 30432 5860 30436
rect 5876 30492 5940 30496
rect 5876 30436 5880 30492
rect 5880 30436 5936 30492
rect 5936 30436 5940 30492
rect 5876 30432 5940 30436
rect 5956 30492 6020 30496
rect 5956 30436 5960 30492
rect 5960 30436 6016 30492
rect 6016 30436 6020 30492
rect 5956 30432 6020 30436
rect 6036 30492 6100 30496
rect 6036 30436 6040 30492
rect 6040 30436 6096 30492
rect 6096 30436 6100 30492
rect 6036 30432 6100 30436
rect 36516 30492 36580 30496
rect 36516 30436 36520 30492
rect 36520 30436 36576 30492
rect 36576 30436 36580 30492
rect 36516 30432 36580 30436
rect 36596 30492 36660 30496
rect 36596 30436 36600 30492
rect 36600 30436 36656 30492
rect 36656 30436 36660 30492
rect 36596 30432 36660 30436
rect 36676 30492 36740 30496
rect 36676 30436 36680 30492
rect 36680 30436 36736 30492
rect 36736 30436 36740 30492
rect 36676 30432 36740 30436
rect 36756 30492 36820 30496
rect 36756 30436 36760 30492
rect 36760 30436 36816 30492
rect 36816 30436 36820 30492
rect 36756 30432 36820 30436
rect 67236 30492 67300 30496
rect 67236 30436 67240 30492
rect 67240 30436 67296 30492
rect 67296 30436 67300 30492
rect 67236 30432 67300 30436
rect 67316 30492 67380 30496
rect 67316 30436 67320 30492
rect 67320 30436 67376 30492
rect 67376 30436 67380 30492
rect 67316 30432 67380 30436
rect 67396 30492 67460 30496
rect 67396 30436 67400 30492
rect 67400 30436 67456 30492
rect 67456 30436 67460 30492
rect 67396 30432 67460 30436
rect 67476 30492 67540 30496
rect 67476 30436 67480 30492
rect 67480 30436 67536 30492
rect 67536 30436 67540 30492
rect 67476 30432 67540 30436
rect 5136 29948 5200 29952
rect 5136 29892 5140 29948
rect 5140 29892 5196 29948
rect 5196 29892 5200 29948
rect 5136 29888 5200 29892
rect 5216 29948 5280 29952
rect 5216 29892 5220 29948
rect 5220 29892 5276 29948
rect 5276 29892 5280 29948
rect 5216 29888 5280 29892
rect 5296 29948 5360 29952
rect 5296 29892 5300 29948
rect 5300 29892 5356 29948
rect 5356 29892 5360 29948
rect 5296 29888 5360 29892
rect 5376 29948 5440 29952
rect 5376 29892 5380 29948
rect 5380 29892 5436 29948
rect 5436 29892 5440 29948
rect 5376 29888 5440 29892
rect 35856 29948 35920 29952
rect 35856 29892 35860 29948
rect 35860 29892 35916 29948
rect 35916 29892 35920 29948
rect 35856 29888 35920 29892
rect 35936 29948 36000 29952
rect 35936 29892 35940 29948
rect 35940 29892 35996 29948
rect 35996 29892 36000 29948
rect 35936 29888 36000 29892
rect 36016 29948 36080 29952
rect 36016 29892 36020 29948
rect 36020 29892 36076 29948
rect 36076 29892 36080 29948
rect 36016 29888 36080 29892
rect 36096 29948 36160 29952
rect 36096 29892 36100 29948
rect 36100 29892 36156 29948
rect 36156 29892 36160 29948
rect 36096 29888 36160 29892
rect 66576 29948 66640 29952
rect 66576 29892 66580 29948
rect 66580 29892 66636 29948
rect 66636 29892 66640 29948
rect 66576 29888 66640 29892
rect 66656 29948 66720 29952
rect 66656 29892 66660 29948
rect 66660 29892 66716 29948
rect 66716 29892 66720 29948
rect 66656 29888 66720 29892
rect 66736 29948 66800 29952
rect 66736 29892 66740 29948
rect 66740 29892 66796 29948
rect 66796 29892 66800 29948
rect 66736 29888 66800 29892
rect 66816 29948 66880 29952
rect 66816 29892 66820 29948
rect 66820 29892 66876 29948
rect 66876 29892 66880 29948
rect 66816 29888 66880 29892
rect 26740 29548 26804 29612
rect 5796 29404 5860 29408
rect 5796 29348 5800 29404
rect 5800 29348 5856 29404
rect 5856 29348 5860 29404
rect 5796 29344 5860 29348
rect 5876 29404 5940 29408
rect 5876 29348 5880 29404
rect 5880 29348 5936 29404
rect 5936 29348 5940 29404
rect 5876 29344 5940 29348
rect 5956 29404 6020 29408
rect 5956 29348 5960 29404
rect 5960 29348 6016 29404
rect 6016 29348 6020 29404
rect 5956 29344 6020 29348
rect 6036 29404 6100 29408
rect 6036 29348 6040 29404
rect 6040 29348 6096 29404
rect 6096 29348 6100 29404
rect 6036 29344 6100 29348
rect 36516 29404 36580 29408
rect 36516 29348 36520 29404
rect 36520 29348 36576 29404
rect 36576 29348 36580 29404
rect 36516 29344 36580 29348
rect 36596 29404 36660 29408
rect 36596 29348 36600 29404
rect 36600 29348 36656 29404
rect 36656 29348 36660 29404
rect 36596 29344 36660 29348
rect 36676 29404 36740 29408
rect 36676 29348 36680 29404
rect 36680 29348 36736 29404
rect 36736 29348 36740 29404
rect 36676 29344 36740 29348
rect 36756 29404 36820 29408
rect 36756 29348 36760 29404
rect 36760 29348 36816 29404
rect 36816 29348 36820 29404
rect 36756 29344 36820 29348
rect 67236 29404 67300 29408
rect 67236 29348 67240 29404
rect 67240 29348 67296 29404
rect 67296 29348 67300 29404
rect 67236 29344 67300 29348
rect 67316 29404 67380 29408
rect 67316 29348 67320 29404
rect 67320 29348 67376 29404
rect 67376 29348 67380 29404
rect 67316 29344 67380 29348
rect 67396 29404 67460 29408
rect 67396 29348 67400 29404
rect 67400 29348 67456 29404
rect 67456 29348 67460 29404
rect 67396 29344 67460 29348
rect 67476 29404 67540 29408
rect 67476 29348 67480 29404
rect 67480 29348 67536 29404
rect 67536 29348 67540 29404
rect 67476 29344 67540 29348
rect 5136 28860 5200 28864
rect 5136 28804 5140 28860
rect 5140 28804 5196 28860
rect 5196 28804 5200 28860
rect 5136 28800 5200 28804
rect 5216 28860 5280 28864
rect 5216 28804 5220 28860
rect 5220 28804 5276 28860
rect 5276 28804 5280 28860
rect 5216 28800 5280 28804
rect 5296 28860 5360 28864
rect 5296 28804 5300 28860
rect 5300 28804 5356 28860
rect 5356 28804 5360 28860
rect 5296 28800 5360 28804
rect 5376 28860 5440 28864
rect 5376 28804 5380 28860
rect 5380 28804 5436 28860
rect 5436 28804 5440 28860
rect 5376 28800 5440 28804
rect 35856 28860 35920 28864
rect 35856 28804 35860 28860
rect 35860 28804 35916 28860
rect 35916 28804 35920 28860
rect 35856 28800 35920 28804
rect 35936 28860 36000 28864
rect 35936 28804 35940 28860
rect 35940 28804 35996 28860
rect 35996 28804 36000 28860
rect 35936 28800 36000 28804
rect 36016 28860 36080 28864
rect 36016 28804 36020 28860
rect 36020 28804 36076 28860
rect 36076 28804 36080 28860
rect 36016 28800 36080 28804
rect 36096 28860 36160 28864
rect 36096 28804 36100 28860
rect 36100 28804 36156 28860
rect 36156 28804 36160 28860
rect 36096 28800 36160 28804
rect 66576 28860 66640 28864
rect 66576 28804 66580 28860
rect 66580 28804 66636 28860
rect 66636 28804 66640 28860
rect 66576 28800 66640 28804
rect 66656 28860 66720 28864
rect 66656 28804 66660 28860
rect 66660 28804 66716 28860
rect 66716 28804 66720 28860
rect 66656 28800 66720 28804
rect 66736 28860 66800 28864
rect 66736 28804 66740 28860
rect 66740 28804 66796 28860
rect 66796 28804 66800 28860
rect 66736 28800 66800 28804
rect 66816 28860 66880 28864
rect 66816 28804 66820 28860
rect 66820 28804 66876 28860
rect 66876 28804 66880 28860
rect 66816 28800 66880 28804
rect 5796 28316 5860 28320
rect 5796 28260 5800 28316
rect 5800 28260 5856 28316
rect 5856 28260 5860 28316
rect 5796 28256 5860 28260
rect 5876 28316 5940 28320
rect 5876 28260 5880 28316
rect 5880 28260 5936 28316
rect 5936 28260 5940 28316
rect 5876 28256 5940 28260
rect 5956 28316 6020 28320
rect 5956 28260 5960 28316
rect 5960 28260 6016 28316
rect 6016 28260 6020 28316
rect 5956 28256 6020 28260
rect 6036 28316 6100 28320
rect 6036 28260 6040 28316
rect 6040 28260 6096 28316
rect 6096 28260 6100 28316
rect 6036 28256 6100 28260
rect 36516 28316 36580 28320
rect 36516 28260 36520 28316
rect 36520 28260 36576 28316
rect 36576 28260 36580 28316
rect 36516 28256 36580 28260
rect 36596 28316 36660 28320
rect 36596 28260 36600 28316
rect 36600 28260 36656 28316
rect 36656 28260 36660 28316
rect 36596 28256 36660 28260
rect 36676 28316 36740 28320
rect 36676 28260 36680 28316
rect 36680 28260 36736 28316
rect 36736 28260 36740 28316
rect 36676 28256 36740 28260
rect 36756 28316 36820 28320
rect 36756 28260 36760 28316
rect 36760 28260 36816 28316
rect 36816 28260 36820 28316
rect 36756 28256 36820 28260
rect 67236 28316 67300 28320
rect 67236 28260 67240 28316
rect 67240 28260 67296 28316
rect 67296 28260 67300 28316
rect 67236 28256 67300 28260
rect 67316 28316 67380 28320
rect 67316 28260 67320 28316
rect 67320 28260 67376 28316
rect 67376 28260 67380 28316
rect 67316 28256 67380 28260
rect 67396 28316 67460 28320
rect 67396 28260 67400 28316
rect 67400 28260 67456 28316
rect 67456 28260 67460 28316
rect 67396 28256 67460 28260
rect 67476 28316 67540 28320
rect 67476 28260 67480 28316
rect 67480 28260 67536 28316
rect 67536 28260 67540 28316
rect 67476 28256 67540 28260
rect 5136 27772 5200 27776
rect 5136 27716 5140 27772
rect 5140 27716 5196 27772
rect 5196 27716 5200 27772
rect 5136 27712 5200 27716
rect 5216 27772 5280 27776
rect 5216 27716 5220 27772
rect 5220 27716 5276 27772
rect 5276 27716 5280 27772
rect 5216 27712 5280 27716
rect 5296 27772 5360 27776
rect 5296 27716 5300 27772
rect 5300 27716 5356 27772
rect 5356 27716 5360 27772
rect 5296 27712 5360 27716
rect 5376 27772 5440 27776
rect 5376 27716 5380 27772
rect 5380 27716 5436 27772
rect 5436 27716 5440 27772
rect 5376 27712 5440 27716
rect 35856 27772 35920 27776
rect 35856 27716 35860 27772
rect 35860 27716 35916 27772
rect 35916 27716 35920 27772
rect 35856 27712 35920 27716
rect 35936 27772 36000 27776
rect 35936 27716 35940 27772
rect 35940 27716 35996 27772
rect 35996 27716 36000 27772
rect 35936 27712 36000 27716
rect 36016 27772 36080 27776
rect 36016 27716 36020 27772
rect 36020 27716 36076 27772
rect 36076 27716 36080 27772
rect 36016 27712 36080 27716
rect 36096 27772 36160 27776
rect 36096 27716 36100 27772
rect 36100 27716 36156 27772
rect 36156 27716 36160 27772
rect 36096 27712 36160 27716
rect 66576 27772 66640 27776
rect 66576 27716 66580 27772
rect 66580 27716 66636 27772
rect 66636 27716 66640 27772
rect 66576 27712 66640 27716
rect 66656 27772 66720 27776
rect 66656 27716 66660 27772
rect 66660 27716 66716 27772
rect 66716 27716 66720 27772
rect 66656 27712 66720 27716
rect 66736 27772 66800 27776
rect 66736 27716 66740 27772
rect 66740 27716 66796 27772
rect 66796 27716 66800 27772
rect 66736 27712 66800 27716
rect 66816 27772 66880 27776
rect 66816 27716 66820 27772
rect 66820 27716 66876 27772
rect 66876 27716 66880 27772
rect 66816 27712 66880 27716
rect 5796 27228 5860 27232
rect 5796 27172 5800 27228
rect 5800 27172 5856 27228
rect 5856 27172 5860 27228
rect 5796 27168 5860 27172
rect 5876 27228 5940 27232
rect 5876 27172 5880 27228
rect 5880 27172 5936 27228
rect 5936 27172 5940 27228
rect 5876 27168 5940 27172
rect 5956 27228 6020 27232
rect 5956 27172 5960 27228
rect 5960 27172 6016 27228
rect 6016 27172 6020 27228
rect 5956 27168 6020 27172
rect 6036 27228 6100 27232
rect 6036 27172 6040 27228
rect 6040 27172 6096 27228
rect 6096 27172 6100 27228
rect 6036 27168 6100 27172
rect 36516 27228 36580 27232
rect 36516 27172 36520 27228
rect 36520 27172 36576 27228
rect 36576 27172 36580 27228
rect 36516 27168 36580 27172
rect 36596 27228 36660 27232
rect 36596 27172 36600 27228
rect 36600 27172 36656 27228
rect 36656 27172 36660 27228
rect 36596 27168 36660 27172
rect 36676 27228 36740 27232
rect 36676 27172 36680 27228
rect 36680 27172 36736 27228
rect 36736 27172 36740 27228
rect 36676 27168 36740 27172
rect 36756 27228 36820 27232
rect 36756 27172 36760 27228
rect 36760 27172 36816 27228
rect 36816 27172 36820 27228
rect 36756 27168 36820 27172
rect 67236 27228 67300 27232
rect 67236 27172 67240 27228
rect 67240 27172 67296 27228
rect 67296 27172 67300 27228
rect 67236 27168 67300 27172
rect 67316 27228 67380 27232
rect 67316 27172 67320 27228
rect 67320 27172 67376 27228
rect 67376 27172 67380 27228
rect 67316 27168 67380 27172
rect 67396 27228 67460 27232
rect 67396 27172 67400 27228
rect 67400 27172 67456 27228
rect 67456 27172 67460 27228
rect 67396 27168 67460 27172
rect 67476 27228 67540 27232
rect 67476 27172 67480 27228
rect 67480 27172 67536 27228
rect 67536 27172 67540 27228
rect 67476 27168 67540 27172
rect 5136 26684 5200 26688
rect 5136 26628 5140 26684
rect 5140 26628 5196 26684
rect 5196 26628 5200 26684
rect 5136 26624 5200 26628
rect 5216 26684 5280 26688
rect 5216 26628 5220 26684
rect 5220 26628 5276 26684
rect 5276 26628 5280 26684
rect 5216 26624 5280 26628
rect 5296 26684 5360 26688
rect 5296 26628 5300 26684
rect 5300 26628 5356 26684
rect 5356 26628 5360 26684
rect 5296 26624 5360 26628
rect 5376 26684 5440 26688
rect 5376 26628 5380 26684
rect 5380 26628 5436 26684
rect 5436 26628 5440 26684
rect 5376 26624 5440 26628
rect 35856 26684 35920 26688
rect 35856 26628 35860 26684
rect 35860 26628 35916 26684
rect 35916 26628 35920 26684
rect 35856 26624 35920 26628
rect 35936 26684 36000 26688
rect 35936 26628 35940 26684
rect 35940 26628 35996 26684
rect 35996 26628 36000 26684
rect 35936 26624 36000 26628
rect 36016 26684 36080 26688
rect 36016 26628 36020 26684
rect 36020 26628 36076 26684
rect 36076 26628 36080 26684
rect 36016 26624 36080 26628
rect 36096 26684 36160 26688
rect 36096 26628 36100 26684
rect 36100 26628 36156 26684
rect 36156 26628 36160 26684
rect 36096 26624 36160 26628
rect 66576 26684 66640 26688
rect 66576 26628 66580 26684
rect 66580 26628 66636 26684
rect 66636 26628 66640 26684
rect 66576 26624 66640 26628
rect 66656 26684 66720 26688
rect 66656 26628 66660 26684
rect 66660 26628 66716 26684
rect 66716 26628 66720 26684
rect 66656 26624 66720 26628
rect 66736 26684 66800 26688
rect 66736 26628 66740 26684
rect 66740 26628 66796 26684
rect 66796 26628 66800 26684
rect 66736 26624 66800 26628
rect 66816 26684 66880 26688
rect 66816 26628 66820 26684
rect 66820 26628 66876 26684
rect 66876 26628 66880 26684
rect 66816 26624 66880 26628
rect 5796 26140 5860 26144
rect 5796 26084 5800 26140
rect 5800 26084 5856 26140
rect 5856 26084 5860 26140
rect 5796 26080 5860 26084
rect 5876 26140 5940 26144
rect 5876 26084 5880 26140
rect 5880 26084 5936 26140
rect 5936 26084 5940 26140
rect 5876 26080 5940 26084
rect 5956 26140 6020 26144
rect 5956 26084 5960 26140
rect 5960 26084 6016 26140
rect 6016 26084 6020 26140
rect 5956 26080 6020 26084
rect 6036 26140 6100 26144
rect 6036 26084 6040 26140
rect 6040 26084 6096 26140
rect 6096 26084 6100 26140
rect 6036 26080 6100 26084
rect 36516 26140 36580 26144
rect 36516 26084 36520 26140
rect 36520 26084 36576 26140
rect 36576 26084 36580 26140
rect 36516 26080 36580 26084
rect 36596 26140 36660 26144
rect 36596 26084 36600 26140
rect 36600 26084 36656 26140
rect 36656 26084 36660 26140
rect 36596 26080 36660 26084
rect 36676 26140 36740 26144
rect 36676 26084 36680 26140
rect 36680 26084 36736 26140
rect 36736 26084 36740 26140
rect 36676 26080 36740 26084
rect 36756 26140 36820 26144
rect 36756 26084 36760 26140
rect 36760 26084 36816 26140
rect 36816 26084 36820 26140
rect 36756 26080 36820 26084
rect 67236 26140 67300 26144
rect 67236 26084 67240 26140
rect 67240 26084 67296 26140
rect 67296 26084 67300 26140
rect 67236 26080 67300 26084
rect 67316 26140 67380 26144
rect 67316 26084 67320 26140
rect 67320 26084 67376 26140
rect 67376 26084 67380 26140
rect 67316 26080 67380 26084
rect 67396 26140 67460 26144
rect 67396 26084 67400 26140
rect 67400 26084 67456 26140
rect 67456 26084 67460 26140
rect 67396 26080 67460 26084
rect 67476 26140 67540 26144
rect 67476 26084 67480 26140
rect 67480 26084 67536 26140
rect 67536 26084 67540 26140
rect 67476 26080 67540 26084
rect 5136 25596 5200 25600
rect 5136 25540 5140 25596
rect 5140 25540 5196 25596
rect 5196 25540 5200 25596
rect 5136 25536 5200 25540
rect 5216 25596 5280 25600
rect 5216 25540 5220 25596
rect 5220 25540 5276 25596
rect 5276 25540 5280 25596
rect 5216 25536 5280 25540
rect 5296 25596 5360 25600
rect 5296 25540 5300 25596
rect 5300 25540 5356 25596
rect 5356 25540 5360 25596
rect 5296 25536 5360 25540
rect 5376 25596 5440 25600
rect 5376 25540 5380 25596
rect 5380 25540 5436 25596
rect 5436 25540 5440 25596
rect 5376 25536 5440 25540
rect 35856 25596 35920 25600
rect 35856 25540 35860 25596
rect 35860 25540 35916 25596
rect 35916 25540 35920 25596
rect 35856 25536 35920 25540
rect 35936 25596 36000 25600
rect 35936 25540 35940 25596
rect 35940 25540 35996 25596
rect 35996 25540 36000 25596
rect 35936 25536 36000 25540
rect 36016 25596 36080 25600
rect 36016 25540 36020 25596
rect 36020 25540 36076 25596
rect 36076 25540 36080 25596
rect 36016 25536 36080 25540
rect 36096 25596 36160 25600
rect 36096 25540 36100 25596
rect 36100 25540 36156 25596
rect 36156 25540 36160 25596
rect 36096 25536 36160 25540
rect 66576 25596 66640 25600
rect 66576 25540 66580 25596
rect 66580 25540 66636 25596
rect 66636 25540 66640 25596
rect 66576 25536 66640 25540
rect 66656 25596 66720 25600
rect 66656 25540 66660 25596
rect 66660 25540 66716 25596
rect 66716 25540 66720 25596
rect 66656 25536 66720 25540
rect 66736 25596 66800 25600
rect 66736 25540 66740 25596
rect 66740 25540 66796 25596
rect 66796 25540 66800 25596
rect 66736 25536 66800 25540
rect 66816 25596 66880 25600
rect 66816 25540 66820 25596
rect 66820 25540 66876 25596
rect 66876 25540 66880 25596
rect 66816 25536 66880 25540
rect 5796 25052 5860 25056
rect 5796 24996 5800 25052
rect 5800 24996 5856 25052
rect 5856 24996 5860 25052
rect 5796 24992 5860 24996
rect 5876 25052 5940 25056
rect 5876 24996 5880 25052
rect 5880 24996 5936 25052
rect 5936 24996 5940 25052
rect 5876 24992 5940 24996
rect 5956 25052 6020 25056
rect 5956 24996 5960 25052
rect 5960 24996 6016 25052
rect 6016 24996 6020 25052
rect 5956 24992 6020 24996
rect 6036 25052 6100 25056
rect 6036 24996 6040 25052
rect 6040 24996 6096 25052
rect 6096 24996 6100 25052
rect 6036 24992 6100 24996
rect 36516 25052 36580 25056
rect 36516 24996 36520 25052
rect 36520 24996 36576 25052
rect 36576 24996 36580 25052
rect 36516 24992 36580 24996
rect 36596 25052 36660 25056
rect 36596 24996 36600 25052
rect 36600 24996 36656 25052
rect 36656 24996 36660 25052
rect 36596 24992 36660 24996
rect 36676 25052 36740 25056
rect 36676 24996 36680 25052
rect 36680 24996 36736 25052
rect 36736 24996 36740 25052
rect 36676 24992 36740 24996
rect 36756 25052 36820 25056
rect 36756 24996 36760 25052
rect 36760 24996 36816 25052
rect 36816 24996 36820 25052
rect 36756 24992 36820 24996
rect 67236 25052 67300 25056
rect 67236 24996 67240 25052
rect 67240 24996 67296 25052
rect 67296 24996 67300 25052
rect 67236 24992 67300 24996
rect 67316 25052 67380 25056
rect 67316 24996 67320 25052
rect 67320 24996 67376 25052
rect 67376 24996 67380 25052
rect 67316 24992 67380 24996
rect 67396 25052 67460 25056
rect 67396 24996 67400 25052
rect 67400 24996 67456 25052
rect 67456 24996 67460 25052
rect 67396 24992 67460 24996
rect 67476 25052 67540 25056
rect 67476 24996 67480 25052
rect 67480 24996 67536 25052
rect 67536 24996 67540 25052
rect 67476 24992 67540 24996
rect 5136 24508 5200 24512
rect 5136 24452 5140 24508
rect 5140 24452 5196 24508
rect 5196 24452 5200 24508
rect 5136 24448 5200 24452
rect 5216 24508 5280 24512
rect 5216 24452 5220 24508
rect 5220 24452 5276 24508
rect 5276 24452 5280 24508
rect 5216 24448 5280 24452
rect 5296 24508 5360 24512
rect 5296 24452 5300 24508
rect 5300 24452 5356 24508
rect 5356 24452 5360 24508
rect 5296 24448 5360 24452
rect 5376 24508 5440 24512
rect 5376 24452 5380 24508
rect 5380 24452 5436 24508
rect 5436 24452 5440 24508
rect 5376 24448 5440 24452
rect 35856 24508 35920 24512
rect 35856 24452 35860 24508
rect 35860 24452 35916 24508
rect 35916 24452 35920 24508
rect 35856 24448 35920 24452
rect 35936 24508 36000 24512
rect 35936 24452 35940 24508
rect 35940 24452 35996 24508
rect 35996 24452 36000 24508
rect 35936 24448 36000 24452
rect 36016 24508 36080 24512
rect 36016 24452 36020 24508
rect 36020 24452 36076 24508
rect 36076 24452 36080 24508
rect 36016 24448 36080 24452
rect 36096 24508 36160 24512
rect 36096 24452 36100 24508
rect 36100 24452 36156 24508
rect 36156 24452 36160 24508
rect 36096 24448 36160 24452
rect 66576 24508 66640 24512
rect 66576 24452 66580 24508
rect 66580 24452 66636 24508
rect 66636 24452 66640 24508
rect 66576 24448 66640 24452
rect 66656 24508 66720 24512
rect 66656 24452 66660 24508
rect 66660 24452 66716 24508
rect 66716 24452 66720 24508
rect 66656 24448 66720 24452
rect 66736 24508 66800 24512
rect 66736 24452 66740 24508
rect 66740 24452 66796 24508
rect 66796 24452 66800 24508
rect 66736 24448 66800 24452
rect 66816 24508 66880 24512
rect 66816 24452 66820 24508
rect 66820 24452 66876 24508
rect 66876 24452 66880 24508
rect 66816 24448 66880 24452
rect 5796 23964 5860 23968
rect 5796 23908 5800 23964
rect 5800 23908 5856 23964
rect 5856 23908 5860 23964
rect 5796 23904 5860 23908
rect 5876 23964 5940 23968
rect 5876 23908 5880 23964
rect 5880 23908 5936 23964
rect 5936 23908 5940 23964
rect 5876 23904 5940 23908
rect 5956 23964 6020 23968
rect 5956 23908 5960 23964
rect 5960 23908 6016 23964
rect 6016 23908 6020 23964
rect 5956 23904 6020 23908
rect 6036 23964 6100 23968
rect 6036 23908 6040 23964
rect 6040 23908 6096 23964
rect 6096 23908 6100 23964
rect 6036 23904 6100 23908
rect 36516 23964 36580 23968
rect 36516 23908 36520 23964
rect 36520 23908 36576 23964
rect 36576 23908 36580 23964
rect 36516 23904 36580 23908
rect 36596 23964 36660 23968
rect 36596 23908 36600 23964
rect 36600 23908 36656 23964
rect 36656 23908 36660 23964
rect 36596 23904 36660 23908
rect 36676 23964 36740 23968
rect 36676 23908 36680 23964
rect 36680 23908 36736 23964
rect 36736 23908 36740 23964
rect 36676 23904 36740 23908
rect 36756 23964 36820 23968
rect 36756 23908 36760 23964
rect 36760 23908 36816 23964
rect 36816 23908 36820 23964
rect 36756 23904 36820 23908
rect 67236 23964 67300 23968
rect 67236 23908 67240 23964
rect 67240 23908 67296 23964
rect 67296 23908 67300 23964
rect 67236 23904 67300 23908
rect 67316 23964 67380 23968
rect 67316 23908 67320 23964
rect 67320 23908 67376 23964
rect 67376 23908 67380 23964
rect 67316 23904 67380 23908
rect 67396 23964 67460 23968
rect 67396 23908 67400 23964
rect 67400 23908 67456 23964
rect 67456 23908 67460 23964
rect 67396 23904 67460 23908
rect 67476 23964 67540 23968
rect 67476 23908 67480 23964
rect 67480 23908 67536 23964
rect 67536 23908 67540 23964
rect 67476 23904 67540 23908
rect 5136 23420 5200 23424
rect 5136 23364 5140 23420
rect 5140 23364 5196 23420
rect 5196 23364 5200 23420
rect 5136 23360 5200 23364
rect 5216 23420 5280 23424
rect 5216 23364 5220 23420
rect 5220 23364 5276 23420
rect 5276 23364 5280 23420
rect 5216 23360 5280 23364
rect 5296 23420 5360 23424
rect 5296 23364 5300 23420
rect 5300 23364 5356 23420
rect 5356 23364 5360 23420
rect 5296 23360 5360 23364
rect 5376 23420 5440 23424
rect 5376 23364 5380 23420
rect 5380 23364 5436 23420
rect 5436 23364 5440 23420
rect 5376 23360 5440 23364
rect 35856 23420 35920 23424
rect 35856 23364 35860 23420
rect 35860 23364 35916 23420
rect 35916 23364 35920 23420
rect 35856 23360 35920 23364
rect 35936 23420 36000 23424
rect 35936 23364 35940 23420
rect 35940 23364 35996 23420
rect 35996 23364 36000 23420
rect 35936 23360 36000 23364
rect 36016 23420 36080 23424
rect 36016 23364 36020 23420
rect 36020 23364 36076 23420
rect 36076 23364 36080 23420
rect 36016 23360 36080 23364
rect 36096 23420 36160 23424
rect 36096 23364 36100 23420
rect 36100 23364 36156 23420
rect 36156 23364 36160 23420
rect 36096 23360 36160 23364
rect 66576 23420 66640 23424
rect 66576 23364 66580 23420
rect 66580 23364 66636 23420
rect 66636 23364 66640 23420
rect 66576 23360 66640 23364
rect 66656 23420 66720 23424
rect 66656 23364 66660 23420
rect 66660 23364 66716 23420
rect 66716 23364 66720 23420
rect 66656 23360 66720 23364
rect 66736 23420 66800 23424
rect 66736 23364 66740 23420
rect 66740 23364 66796 23420
rect 66796 23364 66800 23420
rect 66736 23360 66800 23364
rect 66816 23420 66880 23424
rect 66816 23364 66820 23420
rect 66820 23364 66876 23420
rect 66876 23364 66880 23420
rect 66816 23360 66880 23364
rect 5796 22876 5860 22880
rect 5796 22820 5800 22876
rect 5800 22820 5856 22876
rect 5856 22820 5860 22876
rect 5796 22816 5860 22820
rect 5876 22876 5940 22880
rect 5876 22820 5880 22876
rect 5880 22820 5936 22876
rect 5936 22820 5940 22876
rect 5876 22816 5940 22820
rect 5956 22876 6020 22880
rect 5956 22820 5960 22876
rect 5960 22820 6016 22876
rect 6016 22820 6020 22876
rect 5956 22816 6020 22820
rect 6036 22876 6100 22880
rect 6036 22820 6040 22876
rect 6040 22820 6096 22876
rect 6096 22820 6100 22876
rect 6036 22816 6100 22820
rect 36516 22876 36580 22880
rect 36516 22820 36520 22876
rect 36520 22820 36576 22876
rect 36576 22820 36580 22876
rect 36516 22816 36580 22820
rect 36596 22876 36660 22880
rect 36596 22820 36600 22876
rect 36600 22820 36656 22876
rect 36656 22820 36660 22876
rect 36596 22816 36660 22820
rect 36676 22876 36740 22880
rect 36676 22820 36680 22876
rect 36680 22820 36736 22876
rect 36736 22820 36740 22876
rect 36676 22816 36740 22820
rect 36756 22876 36820 22880
rect 36756 22820 36760 22876
rect 36760 22820 36816 22876
rect 36816 22820 36820 22876
rect 36756 22816 36820 22820
rect 67236 22876 67300 22880
rect 67236 22820 67240 22876
rect 67240 22820 67296 22876
rect 67296 22820 67300 22876
rect 67236 22816 67300 22820
rect 67316 22876 67380 22880
rect 67316 22820 67320 22876
rect 67320 22820 67376 22876
rect 67376 22820 67380 22876
rect 67316 22816 67380 22820
rect 67396 22876 67460 22880
rect 67396 22820 67400 22876
rect 67400 22820 67456 22876
rect 67456 22820 67460 22876
rect 67396 22816 67460 22820
rect 67476 22876 67540 22880
rect 67476 22820 67480 22876
rect 67480 22820 67536 22876
rect 67536 22820 67540 22876
rect 67476 22816 67540 22820
rect 5136 22332 5200 22336
rect 5136 22276 5140 22332
rect 5140 22276 5196 22332
rect 5196 22276 5200 22332
rect 5136 22272 5200 22276
rect 5216 22332 5280 22336
rect 5216 22276 5220 22332
rect 5220 22276 5276 22332
rect 5276 22276 5280 22332
rect 5216 22272 5280 22276
rect 5296 22332 5360 22336
rect 5296 22276 5300 22332
rect 5300 22276 5356 22332
rect 5356 22276 5360 22332
rect 5296 22272 5360 22276
rect 5376 22332 5440 22336
rect 5376 22276 5380 22332
rect 5380 22276 5436 22332
rect 5436 22276 5440 22332
rect 5376 22272 5440 22276
rect 35856 22332 35920 22336
rect 35856 22276 35860 22332
rect 35860 22276 35916 22332
rect 35916 22276 35920 22332
rect 35856 22272 35920 22276
rect 35936 22332 36000 22336
rect 35936 22276 35940 22332
rect 35940 22276 35996 22332
rect 35996 22276 36000 22332
rect 35936 22272 36000 22276
rect 36016 22332 36080 22336
rect 36016 22276 36020 22332
rect 36020 22276 36076 22332
rect 36076 22276 36080 22332
rect 36016 22272 36080 22276
rect 36096 22332 36160 22336
rect 36096 22276 36100 22332
rect 36100 22276 36156 22332
rect 36156 22276 36160 22332
rect 36096 22272 36160 22276
rect 66576 22332 66640 22336
rect 66576 22276 66580 22332
rect 66580 22276 66636 22332
rect 66636 22276 66640 22332
rect 66576 22272 66640 22276
rect 66656 22332 66720 22336
rect 66656 22276 66660 22332
rect 66660 22276 66716 22332
rect 66716 22276 66720 22332
rect 66656 22272 66720 22276
rect 66736 22332 66800 22336
rect 66736 22276 66740 22332
rect 66740 22276 66796 22332
rect 66796 22276 66800 22332
rect 66736 22272 66800 22276
rect 66816 22332 66880 22336
rect 66816 22276 66820 22332
rect 66820 22276 66876 22332
rect 66876 22276 66880 22332
rect 66816 22272 66880 22276
rect 5796 21788 5860 21792
rect 5796 21732 5800 21788
rect 5800 21732 5856 21788
rect 5856 21732 5860 21788
rect 5796 21728 5860 21732
rect 5876 21788 5940 21792
rect 5876 21732 5880 21788
rect 5880 21732 5936 21788
rect 5936 21732 5940 21788
rect 5876 21728 5940 21732
rect 5956 21788 6020 21792
rect 5956 21732 5960 21788
rect 5960 21732 6016 21788
rect 6016 21732 6020 21788
rect 5956 21728 6020 21732
rect 6036 21788 6100 21792
rect 6036 21732 6040 21788
rect 6040 21732 6096 21788
rect 6096 21732 6100 21788
rect 6036 21728 6100 21732
rect 36516 21788 36580 21792
rect 36516 21732 36520 21788
rect 36520 21732 36576 21788
rect 36576 21732 36580 21788
rect 36516 21728 36580 21732
rect 36596 21788 36660 21792
rect 36596 21732 36600 21788
rect 36600 21732 36656 21788
rect 36656 21732 36660 21788
rect 36596 21728 36660 21732
rect 36676 21788 36740 21792
rect 36676 21732 36680 21788
rect 36680 21732 36736 21788
rect 36736 21732 36740 21788
rect 36676 21728 36740 21732
rect 36756 21788 36820 21792
rect 36756 21732 36760 21788
rect 36760 21732 36816 21788
rect 36816 21732 36820 21788
rect 36756 21728 36820 21732
rect 67236 21788 67300 21792
rect 67236 21732 67240 21788
rect 67240 21732 67296 21788
rect 67296 21732 67300 21788
rect 67236 21728 67300 21732
rect 67316 21788 67380 21792
rect 67316 21732 67320 21788
rect 67320 21732 67376 21788
rect 67376 21732 67380 21788
rect 67316 21728 67380 21732
rect 67396 21788 67460 21792
rect 67396 21732 67400 21788
rect 67400 21732 67456 21788
rect 67456 21732 67460 21788
rect 67396 21728 67460 21732
rect 67476 21788 67540 21792
rect 67476 21732 67480 21788
rect 67480 21732 67536 21788
rect 67536 21732 67540 21788
rect 67476 21728 67540 21732
rect 5136 21244 5200 21248
rect 5136 21188 5140 21244
rect 5140 21188 5196 21244
rect 5196 21188 5200 21244
rect 5136 21184 5200 21188
rect 5216 21244 5280 21248
rect 5216 21188 5220 21244
rect 5220 21188 5276 21244
rect 5276 21188 5280 21244
rect 5216 21184 5280 21188
rect 5296 21244 5360 21248
rect 5296 21188 5300 21244
rect 5300 21188 5356 21244
rect 5356 21188 5360 21244
rect 5296 21184 5360 21188
rect 5376 21244 5440 21248
rect 5376 21188 5380 21244
rect 5380 21188 5436 21244
rect 5436 21188 5440 21244
rect 5376 21184 5440 21188
rect 35856 21244 35920 21248
rect 35856 21188 35860 21244
rect 35860 21188 35916 21244
rect 35916 21188 35920 21244
rect 35856 21184 35920 21188
rect 35936 21244 36000 21248
rect 35936 21188 35940 21244
rect 35940 21188 35996 21244
rect 35996 21188 36000 21244
rect 35936 21184 36000 21188
rect 36016 21244 36080 21248
rect 36016 21188 36020 21244
rect 36020 21188 36076 21244
rect 36076 21188 36080 21244
rect 36016 21184 36080 21188
rect 36096 21244 36160 21248
rect 36096 21188 36100 21244
rect 36100 21188 36156 21244
rect 36156 21188 36160 21244
rect 36096 21184 36160 21188
rect 66576 21244 66640 21248
rect 66576 21188 66580 21244
rect 66580 21188 66636 21244
rect 66636 21188 66640 21244
rect 66576 21184 66640 21188
rect 66656 21244 66720 21248
rect 66656 21188 66660 21244
rect 66660 21188 66716 21244
rect 66716 21188 66720 21244
rect 66656 21184 66720 21188
rect 66736 21244 66800 21248
rect 66736 21188 66740 21244
rect 66740 21188 66796 21244
rect 66796 21188 66800 21244
rect 66736 21184 66800 21188
rect 66816 21244 66880 21248
rect 66816 21188 66820 21244
rect 66820 21188 66876 21244
rect 66876 21188 66880 21244
rect 66816 21184 66880 21188
rect 5796 20700 5860 20704
rect 5796 20644 5800 20700
rect 5800 20644 5856 20700
rect 5856 20644 5860 20700
rect 5796 20640 5860 20644
rect 5876 20700 5940 20704
rect 5876 20644 5880 20700
rect 5880 20644 5936 20700
rect 5936 20644 5940 20700
rect 5876 20640 5940 20644
rect 5956 20700 6020 20704
rect 5956 20644 5960 20700
rect 5960 20644 6016 20700
rect 6016 20644 6020 20700
rect 5956 20640 6020 20644
rect 6036 20700 6100 20704
rect 6036 20644 6040 20700
rect 6040 20644 6096 20700
rect 6096 20644 6100 20700
rect 6036 20640 6100 20644
rect 36516 20700 36580 20704
rect 36516 20644 36520 20700
rect 36520 20644 36576 20700
rect 36576 20644 36580 20700
rect 36516 20640 36580 20644
rect 36596 20700 36660 20704
rect 36596 20644 36600 20700
rect 36600 20644 36656 20700
rect 36656 20644 36660 20700
rect 36596 20640 36660 20644
rect 36676 20700 36740 20704
rect 36676 20644 36680 20700
rect 36680 20644 36736 20700
rect 36736 20644 36740 20700
rect 36676 20640 36740 20644
rect 36756 20700 36820 20704
rect 36756 20644 36760 20700
rect 36760 20644 36816 20700
rect 36816 20644 36820 20700
rect 36756 20640 36820 20644
rect 67236 20700 67300 20704
rect 67236 20644 67240 20700
rect 67240 20644 67296 20700
rect 67296 20644 67300 20700
rect 67236 20640 67300 20644
rect 67316 20700 67380 20704
rect 67316 20644 67320 20700
rect 67320 20644 67376 20700
rect 67376 20644 67380 20700
rect 67316 20640 67380 20644
rect 67396 20700 67460 20704
rect 67396 20644 67400 20700
rect 67400 20644 67456 20700
rect 67456 20644 67460 20700
rect 67396 20640 67460 20644
rect 67476 20700 67540 20704
rect 67476 20644 67480 20700
rect 67480 20644 67536 20700
rect 67536 20644 67540 20700
rect 67476 20640 67540 20644
rect 5136 20156 5200 20160
rect 5136 20100 5140 20156
rect 5140 20100 5196 20156
rect 5196 20100 5200 20156
rect 5136 20096 5200 20100
rect 5216 20156 5280 20160
rect 5216 20100 5220 20156
rect 5220 20100 5276 20156
rect 5276 20100 5280 20156
rect 5216 20096 5280 20100
rect 5296 20156 5360 20160
rect 5296 20100 5300 20156
rect 5300 20100 5356 20156
rect 5356 20100 5360 20156
rect 5296 20096 5360 20100
rect 5376 20156 5440 20160
rect 5376 20100 5380 20156
rect 5380 20100 5436 20156
rect 5436 20100 5440 20156
rect 5376 20096 5440 20100
rect 35856 20156 35920 20160
rect 35856 20100 35860 20156
rect 35860 20100 35916 20156
rect 35916 20100 35920 20156
rect 35856 20096 35920 20100
rect 35936 20156 36000 20160
rect 35936 20100 35940 20156
rect 35940 20100 35996 20156
rect 35996 20100 36000 20156
rect 35936 20096 36000 20100
rect 36016 20156 36080 20160
rect 36016 20100 36020 20156
rect 36020 20100 36076 20156
rect 36076 20100 36080 20156
rect 36016 20096 36080 20100
rect 36096 20156 36160 20160
rect 36096 20100 36100 20156
rect 36100 20100 36156 20156
rect 36156 20100 36160 20156
rect 36096 20096 36160 20100
rect 66576 20156 66640 20160
rect 66576 20100 66580 20156
rect 66580 20100 66636 20156
rect 66636 20100 66640 20156
rect 66576 20096 66640 20100
rect 66656 20156 66720 20160
rect 66656 20100 66660 20156
rect 66660 20100 66716 20156
rect 66716 20100 66720 20156
rect 66656 20096 66720 20100
rect 66736 20156 66800 20160
rect 66736 20100 66740 20156
rect 66740 20100 66796 20156
rect 66796 20100 66800 20156
rect 66736 20096 66800 20100
rect 66816 20156 66880 20160
rect 66816 20100 66820 20156
rect 66820 20100 66876 20156
rect 66876 20100 66880 20156
rect 66816 20096 66880 20100
rect 5796 19612 5860 19616
rect 5796 19556 5800 19612
rect 5800 19556 5856 19612
rect 5856 19556 5860 19612
rect 5796 19552 5860 19556
rect 5876 19612 5940 19616
rect 5876 19556 5880 19612
rect 5880 19556 5936 19612
rect 5936 19556 5940 19612
rect 5876 19552 5940 19556
rect 5956 19612 6020 19616
rect 5956 19556 5960 19612
rect 5960 19556 6016 19612
rect 6016 19556 6020 19612
rect 5956 19552 6020 19556
rect 6036 19612 6100 19616
rect 6036 19556 6040 19612
rect 6040 19556 6096 19612
rect 6096 19556 6100 19612
rect 6036 19552 6100 19556
rect 36516 19612 36580 19616
rect 36516 19556 36520 19612
rect 36520 19556 36576 19612
rect 36576 19556 36580 19612
rect 36516 19552 36580 19556
rect 36596 19612 36660 19616
rect 36596 19556 36600 19612
rect 36600 19556 36656 19612
rect 36656 19556 36660 19612
rect 36596 19552 36660 19556
rect 36676 19612 36740 19616
rect 36676 19556 36680 19612
rect 36680 19556 36736 19612
rect 36736 19556 36740 19612
rect 36676 19552 36740 19556
rect 36756 19612 36820 19616
rect 36756 19556 36760 19612
rect 36760 19556 36816 19612
rect 36816 19556 36820 19612
rect 36756 19552 36820 19556
rect 67236 19612 67300 19616
rect 67236 19556 67240 19612
rect 67240 19556 67296 19612
rect 67296 19556 67300 19612
rect 67236 19552 67300 19556
rect 67316 19612 67380 19616
rect 67316 19556 67320 19612
rect 67320 19556 67376 19612
rect 67376 19556 67380 19612
rect 67316 19552 67380 19556
rect 67396 19612 67460 19616
rect 67396 19556 67400 19612
rect 67400 19556 67456 19612
rect 67456 19556 67460 19612
rect 67396 19552 67460 19556
rect 67476 19612 67540 19616
rect 67476 19556 67480 19612
rect 67480 19556 67536 19612
rect 67536 19556 67540 19612
rect 67476 19552 67540 19556
rect 5136 19068 5200 19072
rect 5136 19012 5140 19068
rect 5140 19012 5196 19068
rect 5196 19012 5200 19068
rect 5136 19008 5200 19012
rect 5216 19068 5280 19072
rect 5216 19012 5220 19068
rect 5220 19012 5276 19068
rect 5276 19012 5280 19068
rect 5216 19008 5280 19012
rect 5296 19068 5360 19072
rect 5296 19012 5300 19068
rect 5300 19012 5356 19068
rect 5356 19012 5360 19068
rect 5296 19008 5360 19012
rect 5376 19068 5440 19072
rect 5376 19012 5380 19068
rect 5380 19012 5436 19068
rect 5436 19012 5440 19068
rect 5376 19008 5440 19012
rect 35856 19068 35920 19072
rect 35856 19012 35860 19068
rect 35860 19012 35916 19068
rect 35916 19012 35920 19068
rect 35856 19008 35920 19012
rect 35936 19068 36000 19072
rect 35936 19012 35940 19068
rect 35940 19012 35996 19068
rect 35996 19012 36000 19068
rect 35936 19008 36000 19012
rect 36016 19068 36080 19072
rect 36016 19012 36020 19068
rect 36020 19012 36076 19068
rect 36076 19012 36080 19068
rect 36016 19008 36080 19012
rect 36096 19068 36160 19072
rect 36096 19012 36100 19068
rect 36100 19012 36156 19068
rect 36156 19012 36160 19068
rect 36096 19008 36160 19012
rect 66576 19068 66640 19072
rect 66576 19012 66580 19068
rect 66580 19012 66636 19068
rect 66636 19012 66640 19068
rect 66576 19008 66640 19012
rect 66656 19068 66720 19072
rect 66656 19012 66660 19068
rect 66660 19012 66716 19068
rect 66716 19012 66720 19068
rect 66656 19008 66720 19012
rect 66736 19068 66800 19072
rect 66736 19012 66740 19068
rect 66740 19012 66796 19068
rect 66796 19012 66800 19068
rect 66736 19008 66800 19012
rect 66816 19068 66880 19072
rect 66816 19012 66820 19068
rect 66820 19012 66876 19068
rect 66876 19012 66880 19068
rect 66816 19008 66880 19012
rect 5796 18524 5860 18528
rect 5796 18468 5800 18524
rect 5800 18468 5856 18524
rect 5856 18468 5860 18524
rect 5796 18464 5860 18468
rect 5876 18524 5940 18528
rect 5876 18468 5880 18524
rect 5880 18468 5936 18524
rect 5936 18468 5940 18524
rect 5876 18464 5940 18468
rect 5956 18524 6020 18528
rect 5956 18468 5960 18524
rect 5960 18468 6016 18524
rect 6016 18468 6020 18524
rect 5956 18464 6020 18468
rect 6036 18524 6100 18528
rect 6036 18468 6040 18524
rect 6040 18468 6096 18524
rect 6096 18468 6100 18524
rect 6036 18464 6100 18468
rect 36516 18524 36580 18528
rect 36516 18468 36520 18524
rect 36520 18468 36576 18524
rect 36576 18468 36580 18524
rect 36516 18464 36580 18468
rect 36596 18524 36660 18528
rect 36596 18468 36600 18524
rect 36600 18468 36656 18524
rect 36656 18468 36660 18524
rect 36596 18464 36660 18468
rect 36676 18524 36740 18528
rect 36676 18468 36680 18524
rect 36680 18468 36736 18524
rect 36736 18468 36740 18524
rect 36676 18464 36740 18468
rect 36756 18524 36820 18528
rect 36756 18468 36760 18524
rect 36760 18468 36816 18524
rect 36816 18468 36820 18524
rect 36756 18464 36820 18468
rect 67236 18524 67300 18528
rect 67236 18468 67240 18524
rect 67240 18468 67296 18524
rect 67296 18468 67300 18524
rect 67236 18464 67300 18468
rect 67316 18524 67380 18528
rect 67316 18468 67320 18524
rect 67320 18468 67376 18524
rect 67376 18468 67380 18524
rect 67316 18464 67380 18468
rect 67396 18524 67460 18528
rect 67396 18468 67400 18524
rect 67400 18468 67456 18524
rect 67456 18468 67460 18524
rect 67396 18464 67460 18468
rect 67476 18524 67540 18528
rect 67476 18468 67480 18524
rect 67480 18468 67536 18524
rect 67536 18468 67540 18524
rect 67476 18464 67540 18468
rect 5136 17980 5200 17984
rect 5136 17924 5140 17980
rect 5140 17924 5196 17980
rect 5196 17924 5200 17980
rect 5136 17920 5200 17924
rect 5216 17980 5280 17984
rect 5216 17924 5220 17980
rect 5220 17924 5276 17980
rect 5276 17924 5280 17980
rect 5216 17920 5280 17924
rect 5296 17980 5360 17984
rect 5296 17924 5300 17980
rect 5300 17924 5356 17980
rect 5356 17924 5360 17980
rect 5296 17920 5360 17924
rect 5376 17980 5440 17984
rect 5376 17924 5380 17980
rect 5380 17924 5436 17980
rect 5436 17924 5440 17980
rect 5376 17920 5440 17924
rect 35856 17980 35920 17984
rect 35856 17924 35860 17980
rect 35860 17924 35916 17980
rect 35916 17924 35920 17980
rect 35856 17920 35920 17924
rect 35936 17980 36000 17984
rect 35936 17924 35940 17980
rect 35940 17924 35996 17980
rect 35996 17924 36000 17980
rect 35936 17920 36000 17924
rect 36016 17980 36080 17984
rect 36016 17924 36020 17980
rect 36020 17924 36076 17980
rect 36076 17924 36080 17980
rect 36016 17920 36080 17924
rect 36096 17980 36160 17984
rect 36096 17924 36100 17980
rect 36100 17924 36156 17980
rect 36156 17924 36160 17980
rect 36096 17920 36160 17924
rect 66576 17980 66640 17984
rect 66576 17924 66580 17980
rect 66580 17924 66636 17980
rect 66636 17924 66640 17980
rect 66576 17920 66640 17924
rect 66656 17980 66720 17984
rect 66656 17924 66660 17980
rect 66660 17924 66716 17980
rect 66716 17924 66720 17980
rect 66656 17920 66720 17924
rect 66736 17980 66800 17984
rect 66736 17924 66740 17980
rect 66740 17924 66796 17980
rect 66796 17924 66800 17980
rect 66736 17920 66800 17924
rect 66816 17980 66880 17984
rect 66816 17924 66820 17980
rect 66820 17924 66876 17980
rect 66876 17924 66880 17980
rect 66816 17920 66880 17924
rect 5796 17436 5860 17440
rect 5796 17380 5800 17436
rect 5800 17380 5856 17436
rect 5856 17380 5860 17436
rect 5796 17376 5860 17380
rect 5876 17436 5940 17440
rect 5876 17380 5880 17436
rect 5880 17380 5936 17436
rect 5936 17380 5940 17436
rect 5876 17376 5940 17380
rect 5956 17436 6020 17440
rect 5956 17380 5960 17436
rect 5960 17380 6016 17436
rect 6016 17380 6020 17436
rect 5956 17376 6020 17380
rect 6036 17436 6100 17440
rect 6036 17380 6040 17436
rect 6040 17380 6096 17436
rect 6096 17380 6100 17436
rect 6036 17376 6100 17380
rect 36516 17436 36580 17440
rect 36516 17380 36520 17436
rect 36520 17380 36576 17436
rect 36576 17380 36580 17436
rect 36516 17376 36580 17380
rect 36596 17436 36660 17440
rect 36596 17380 36600 17436
rect 36600 17380 36656 17436
rect 36656 17380 36660 17436
rect 36596 17376 36660 17380
rect 36676 17436 36740 17440
rect 36676 17380 36680 17436
rect 36680 17380 36736 17436
rect 36736 17380 36740 17436
rect 36676 17376 36740 17380
rect 36756 17436 36820 17440
rect 36756 17380 36760 17436
rect 36760 17380 36816 17436
rect 36816 17380 36820 17436
rect 36756 17376 36820 17380
rect 67236 17436 67300 17440
rect 67236 17380 67240 17436
rect 67240 17380 67296 17436
rect 67296 17380 67300 17436
rect 67236 17376 67300 17380
rect 67316 17436 67380 17440
rect 67316 17380 67320 17436
rect 67320 17380 67376 17436
rect 67376 17380 67380 17436
rect 67316 17376 67380 17380
rect 67396 17436 67460 17440
rect 67396 17380 67400 17436
rect 67400 17380 67456 17436
rect 67456 17380 67460 17436
rect 67396 17376 67460 17380
rect 67476 17436 67540 17440
rect 67476 17380 67480 17436
rect 67480 17380 67536 17436
rect 67536 17380 67540 17436
rect 67476 17376 67540 17380
rect 5136 16892 5200 16896
rect 5136 16836 5140 16892
rect 5140 16836 5196 16892
rect 5196 16836 5200 16892
rect 5136 16832 5200 16836
rect 5216 16892 5280 16896
rect 5216 16836 5220 16892
rect 5220 16836 5276 16892
rect 5276 16836 5280 16892
rect 5216 16832 5280 16836
rect 5296 16892 5360 16896
rect 5296 16836 5300 16892
rect 5300 16836 5356 16892
rect 5356 16836 5360 16892
rect 5296 16832 5360 16836
rect 5376 16892 5440 16896
rect 5376 16836 5380 16892
rect 5380 16836 5436 16892
rect 5436 16836 5440 16892
rect 5376 16832 5440 16836
rect 35856 16892 35920 16896
rect 35856 16836 35860 16892
rect 35860 16836 35916 16892
rect 35916 16836 35920 16892
rect 35856 16832 35920 16836
rect 35936 16892 36000 16896
rect 35936 16836 35940 16892
rect 35940 16836 35996 16892
rect 35996 16836 36000 16892
rect 35936 16832 36000 16836
rect 36016 16892 36080 16896
rect 36016 16836 36020 16892
rect 36020 16836 36076 16892
rect 36076 16836 36080 16892
rect 36016 16832 36080 16836
rect 36096 16892 36160 16896
rect 36096 16836 36100 16892
rect 36100 16836 36156 16892
rect 36156 16836 36160 16892
rect 36096 16832 36160 16836
rect 66576 16892 66640 16896
rect 66576 16836 66580 16892
rect 66580 16836 66636 16892
rect 66636 16836 66640 16892
rect 66576 16832 66640 16836
rect 66656 16892 66720 16896
rect 66656 16836 66660 16892
rect 66660 16836 66716 16892
rect 66716 16836 66720 16892
rect 66656 16832 66720 16836
rect 66736 16892 66800 16896
rect 66736 16836 66740 16892
rect 66740 16836 66796 16892
rect 66796 16836 66800 16892
rect 66736 16832 66800 16836
rect 66816 16892 66880 16896
rect 66816 16836 66820 16892
rect 66820 16836 66876 16892
rect 66876 16836 66880 16892
rect 66816 16832 66880 16836
rect 5796 16348 5860 16352
rect 5796 16292 5800 16348
rect 5800 16292 5856 16348
rect 5856 16292 5860 16348
rect 5796 16288 5860 16292
rect 5876 16348 5940 16352
rect 5876 16292 5880 16348
rect 5880 16292 5936 16348
rect 5936 16292 5940 16348
rect 5876 16288 5940 16292
rect 5956 16348 6020 16352
rect 5956 16292 5960 16348
rect 5960 16292 6016 16348
rect 6016 16292 6020 16348
rect 5956 16288 6020 16292
rect 6036 16348 6100 16352
rect 6036 16292 6040 16348
rect 6040 16292 6096 16348
rect 6096 16292 6100 16348
rect 6036 16288 6100 16292
rect 36516 16348 36580 16352
rect 36516 16292 36520 16348
rect 36520 16292 36576 16348
rect 36576 16292 36580 16348
rect 36516 16288 36580 16292
rect 36596 16348 36660 16352
rect 36596 16292 36600 16348
rect 36600 16292 36656 16348
rect 36656 16292 36660 16348
rect 36596 16288 36660 16292
rect 36676 16348 36740 16352
rect 36676 16292 36680 16348
rect 36680 16292 36736 16348
rect 36736 16292 36740 16348
rect 36676 16288 36740 16292
rect 36756 16348 36820 16352
rect 36756 16292 36760 16348
rect 36760 16292 36816 16348
rect 36816 16292 36820 16348
rect 36756 16288 36820 16292
rect 67236 16348 67300 16352
rect 67236 16292 67240 16348
rect 67240 16292 67296 16348
rect 67296 16292 67300 16348
rect 67236 16288 67300 16292
rect 67316 16348 67380 16352
rect 67316 16292 67320 16348
rect 67320 16292 67376 16348
rect 67376 16292 67380 16348
rect 67316 16288 67380 16292
rect 67396 16348 67460 16352
rect 67396 16292 67400 16348
rect 67400 16292 67456 16348
rect 67456 16292 67460 16348
rect 67396 16288 67460 16292
rect 67476 16348 67540 16352
rect 67476 16292 67480 16348
rect 67480 16292 67536 16348
rect 67536 16292 67540 16348
rect 67476 16288 67540 16292
rect 5136 15804 5200 15808
rect 5136 15748 5140 15804
rect 5140 15748 5196 15804
rect 5196 15748 5200 15804
rect 5136 15744 5200 15748
rect 5216 15804 5280 15808
rect 5216 15748 5220 15804
rect 5220 15748 5276 15804
rect 5276 15748 5280 15804
rect 5216 15744 5280 15748
rect 5296 15804 5360 15808
rect 5296 15748 5300 15804
rect 5300 15748 5356 15804
rect 5356 15748 5360 15804
rect 5296 15744 5360 15748
rect 5376 15804 5440 15808
rect 5376 15748 5380 15804
rect 5380 15748 5436 15804
rect 5436 15748 5440 15804
rect 5376 15744 5440 15748
rect 35856 15804 35920 15808
rect 35856 15748 35860 15804
rect 35860 15748 35916 15804
rect 35916 15748 35920 15804
rect 35856 15744 35920 15748
rect 35936 15804 36000 15808
rect 35936 15748 35940 15804
rect 35940 15748 35996 15804
rect 35996 15748 36000 15804
rect 35936 15744 36000 15748
rect 36016 15804 36080 15808
rect 36016 15748 36020 15804
rect 36020 15748 36076 15804
rect 36076 15748 36080 15804
rect 36016 15744 36080 15748
rect 36096 15804 36160 15808
rect 36096 15748 36100 15804
rect 36100 15748 36156 15804
rect 36156 15748 36160 15804
rect 36096 15744 36160 15748
rect 66576 15804 66640 15808
rect 66576 15748 66580 15804
rect 66580 15748 66636 15804
rect 66636 15748 66640 15804
rect 66576 15744 66640 15748
rect 66656 15804 66720 15808
rect 66656 15748 66660 15804
rect 66660 15748 66716 15804
rect 66716 15748 66720 15804
rect 66656 15744 66720 15748
rect 66736 15804 66800 15808
rect 66736 15748 66740 15804
rect 66740 15748 66796 15804
rect 66796 15748 66800 15804
rect 66736 15744 66800 15748
rect 66816 15804 66880 15808
rect 66816 15748 66820 15804
rect 66820 15748 66876 15804
rect 66876 15748 66880 15804
rect 66816 15744 66880 15748
rect 5796 15260 5860 15264
rect 5796 15204 5800 15260
rect 5800 15204 5856 15260
rect 5856 15204 5860 15260
rect 5796 15200 5860 15204
rect 5876 15260 5940 15264
rect 5876 15204 5880 15260
rect 5880 15204 5936 15260
rect 5936 15204 5940 15260
rect 5876 15200 5940 15204
rect 5956 15260 6020 15264
rect 5956 15204 5960 15260
rect 5960 15204 6016 15260
rect 6016 15204 6020 15260
rect 5956 15200 6020 15204
rect 6036 15260 6100 15264
rect 6036 15204 6040 15260
rect 6040 15204 6096 15260
rect 6096 15204 6100 15260
rect 6036 15200 6100 15204
rect 36516 15260 36580 15264
rect 36516 15204 36520 15260
rect 36520 15204 36576 15260
rect 36576 15204 36580 15260
rect 36516 15200 36580 15204
rect 36596 15260 36660 15264
rect 36596 15204 36600 15260
rect 36600 15204 36656 15260
rect 36656 15204 36660 15260
rect 36596 15200 36660 15204
rect 36676 15260 36740 15264
rect 36676 15204 36680 15260
rect 36680 15204 36736 15260
rect 36736 15204 36740 15260
rect 36676 15200 36740 15204
rect 36756 15260 36820 15264
rect 36756 15204 36760 15260
rect 36760 15204 36816 15260
rect 36816 15204 36820 15260
rect 36756 15200 36820 15204
rect 67236 15260 67300 15264
rect 67236 15204 67240 15260
rect 67240 15204 67296 15260
rect 67296 15204 67300 15260
rect 67236 15200 67300 15204
rect 67316 15260 67380 15264
rect 67316 15204 67320 15260
rect 67320 15204 67376 15260
rect 67376 15204 67380 15260
rect 67316 15200 67380 15204
rect 67396 15260 67460 15264
rect 67396 15204 67400 15260
rect 67400 15204 67456 15260
rect 67456 15204 67460 15260
rect 67396 15200 67460 15204
rect 67476 15260 67540 15264
rect 67476 15204 67480 15260
rect 67480 15204 67536 15260
rect 67536 15204 67540 15260
rect 67476 15200 67540 15204
rect 5136 14716 5200 14720
rect 5136 14660 5140 14716
rect 5140 14660 5196 14716
rect 5196 14660 5200 14716
rect 5136 14656 5200 14660
rect 5216 14716 5280 14720
rect 5216 14660 5220 14716
rect 5220 14660 5276 14716
rect 5276 14660 5280 14716
rect 5216 14656 5280 14660
rect 5296 14716 5360 14720
rect 5296 14660 5300 14716
rect 5300 14660 5356 14716
rect 5356 14660 5360 14716
rect 5296 14656 5360 14660
rect 5376 14716 5440 14720
rect 5376 14660 5380 14716
rect 5380 14660 5436 14716
rect 5436 14660 5440 14716
rect 5376 14656 5440 14660
rect 35856 14716 35920 14720
rect 35856 14660 35860 14716
rect 35860 14660 35916 14716
rect 35916 14660 35920 14716
rect 35856 14656 35920 14660
rect 35936 14716 36000 14720
rect 35936 14660 35940 14716
rect 35940 14660 35996 14716
rect 35996 14660 36000 14716
rect 35936 14656 36000 14660
rect 36016 14716 36080 14720
rect 36016 14660 36020 14716
rect 36020 14660 36076 14716
rect 36076 14660 36080 14716
rect 36016 14656 36080 14660
rect 36096 14716 36160 14720
rect 36096 14660 36100 14716
rect 36100 14660 36156 14716
rect 36156 14660 36160 14716
rect 36096 14656 36160 14660
rect 66576 14716 66640 14720
rect 66576 14660 66580 14716
rect 66580 14660 66636 14716
rect 66636 14660 66640 14716
rect 66576 14656 66640 14660
rect 66656 14716 66720 14720
rect 66656 14660 66660 14716
rect 66660 14660 66716 14716
rect 66716 14660 66720 14716
rect 66656 14656 66720 14660
rect 66736 14716 66800 14720
rect 66736 14660 66740 14716
rect 66740 14660 66796 14716
rect 66796 14660 66800 14716
rect 66736 14656 66800 14660
rect 66816 14716 66880 14720
rect 66816 14660 66820 14716
rect 66820 14660 66876 14716
rect 66876 14660 66880 14716
rect 66816 14656 66880 14660
rect 5796 14172 5860 14176
rect 5796 14116 5800 14172
rect 5800 14116 5856 14172
rect 5856 14116 5860 14172
rect 5796 14112 5860 14116
rect 5876 14172 5940 14176
rect 5876 14116 5880 14172
rect 5880 14116 5936 14172
rect 5936 14116 5940 14172
rect 5876 14112 5940 14116
rect 5956 14172 6020 14176
rect 5956 14116 5960 14172
rect 5960 14116 6016 14172
rect 6016 14116 6020 14172
rect 5956 14112 6020 14116
rect 6036 14172 6100 14176
rect 6036 14116 6040 14172
rect 6040 14116 6096 14172
rect 6096 14116 6100 14172
rect 6036 14112 6100 14116
rect 36516 14172 36580 14176
rect 36516 14116 36520 14172
rect 36520 14116 36576 14172
rect 36576 14116 36580 14172
rect 36516 14112 36580 14116
rect 36596 14172 36660 14176
rect 36596 14116 36600 14172
rect 36600 14116 36656 14172
rect 36656 14116 36660 14172
rect 36596 14112 36660 14116
rect 36676 14172 36740 14176
rect 36676 14116 36680 14172
rect 36680 14116 36736 14172
rect 36736 14116 36740 14172
rect 36676 14112 36740 14116
rect 36756 14172 36820 14176
rect 36756 14116 36760 14172
rect 36760 14116 36816 14172
rect 36816 14116 36820 14172
rect 36756 14112 36820 14116
rect 67236 14172 67300 14176
rect 67236 14116 67240 14172
rect 67240 14116 67296 14172
rect 67296 14116 67300 14172
rect 67236 14112 67300 14116
rect 67316 14172 67380 14176
rect 67316 14116 67320 14172
rect 67320 14116 67376 14172
rect 67376 14116 67380 14172
rect 67316 14112 67380 14116
rect 67396 14172 67460 14176
rect 67396 14116 67400 14172
rect 67400 14116 67456 14172
rect 67456 14116 67460 14172
rect 67396 14112 67460 14116
rect 67476 14172 67540 14176
rect 67476 14116 67480 14172
rect 67480 14116 67536 14172
rect 67536 14116 67540 14172
rect 67476 14112 67540 14116
rect 5136 13628 5200 13632
rect 5136 13572 5140 13628
rect 5140 13572 5196 13628
rect 5196 13572 5200 13628
rect 5136 13568 5200 13572
rect 5216 13628 5280 13632
rect 5216 13572 5220 13628
rect 5220 13572 5276 13628
rect 5276 13572 5280 13628
rect 5216 13568 5280 13572
rect 5296 13628 5360 13632
rect 5296 13572 5300 13628
rect 5300 13572 5356 13628
rect 5356 13572 5360 13628
rect 5296 13568 5360 13572
rect 5376 13628 5440 13632
rect 5376 13572 5380 13628
rect 5380 13572 5436 13628
rect 5436 13572 5440 13628
rect 5376 13568 5440 13572
rect 35856 13628 35920 13632
rect 35856 13572 35860 13628
rect 35860 13572 35916 13628
rect 35916 13572 35920 13628
rect 35856 13568 35920 13572
rect 35936 13628 36000 13632
rect 35936 13572 35940 13628
rect 35940 13572 35996 13628
rect 35996 13572 36000 13628
rect 35936 13568 36000 13572
rect 36016 13628 36080 13632
rect 36016 13572 36020 13628
rect 36020 13572 36076 13628
rect 36076 13572 36080 13628
rect 36016 13568 36080 13572
rect 36096 13628 36160 13632
rect 36096 13572 36100 13628
rect 36100 13572 36156 13628
rect 36156 13572 36160 13628
rect 36096 13568 36160 13572
rect 66576 13628 66640 13632
rect 66576 13572 66580 13628
rect 66580 13572 66636 13628
rect 66636 13572 66640 13628
rect 66576 13568 66640 13572
rect 66656 13628 66720 13632
rect 66656 13572 66660 13628
rect 66660 13572 66716 13628
rect 66716 13572 66720 13628
rect 66656 13568 66720 13572
rect 66736 13628 66800 13632
rect 66736 13572 66740 13628
rect 66740 13572 66796 13628
rect 66796 13572 66800 13628
rect 66736 13568 66800 13572
rect 66816 13628 66880 13632
rect 66816 13572 66820 13628
rect 66820 13572 66876 13628
rect 66876 13572 66880 13628
rect 66816 13568 66880 13572
rect 5796 13084 5860 13088
rect 5796 13028 5800 13084
rect 5800 13028 5856 13084
rect 5856 13028 5860 13084
rect 5796 13024 5860 13028
rect 5876 13084 5940 13088
rect 5876 13028 5880 13084
rect 5880 13028 5936 13084
rect 5936 13028 5940 13084
rect 5876 13024 5940 13028
rect 5956 13084 6020 13088
rect 5956 13028 5960 13084
rect 5960 13028 6016 13084
rect 6016 13028 6020 13084
rect 5956 13024 6020 13028
rect 6036 13084 6100 13088
rect 6036 13028 6040 13084
rect 6040 13028 6096 13084
rect 6096 13028 6100 13084
rect 6036 13024 6100 13028
rect 36516 13084 36580 13088
rect 36516 13028 36520 13084
rect 36520 13028 36576 13084
rect 36576 13028 36580 13084
rect 36516 13024 36580 13028
rect 36596 13084 36660 13088
rect 36596 13028 36600 13084
rect 36600 13028 36656 13084
rect 36656 13028 36660 13084
rect 36596 13024 36660 13028
rect 36676 13084 36740 13088
rect 36676 13028 36680 13084
rect 36680 13028 36736 13084
rect 36736 13028 36740 13084
rect 36676 13024 36740 13028
rect 36756 13084 36820 13088
rect 36756 13028 36760 13084
rect 36760 13028 36816 13084
rect 36816 13028 36820 13084
rect 36756 13024 36820 13028
rect 67236 13084 67300 13088
rect 67236 13028 67240 13084
rect 67240 13028 67296 13084
rect 67296 13028 67300 13084
rect 67236 13024 67300 13028
rect 67316 13084 67380 13088
rect 67316 13028 67320 13084
rect 67320 13028 67376 13084
rect 67376 13028 67380 13084
rect 67316 13024 67380 13028
rect 67396 13084 67460 13088
rect 67396 13028 67400 13084
rect 67400 13028 67456 13084
rect 67456 13028 67460 13084
rect 67396 13024 67460 13028
rect 67476 13084 67540 13088
rect 67476 13028 67480 13084
rect 67480 13028 67536 13084
rect 67536 13028 67540 13084
rect 67476 13024 67540 13028
rect 5136 12540 5200 12544
rect 5136 12484 5140 12540
rect 5140 12484 5196 12540
rect 5196 12484 5200 12540
rect 5136 12480 5200 12484
rect 5216 12540 5280 12544
rect 5216 12484 5220 12540
rect 5220 12484 5276 12540
rect 5276 12484 5280 12540
rect 5216 12480 5280 12484
rect 5296 12540 5360 12544
rect 5296 12484 5300 12540
rect 5300 12484 5356 12540
rect 5356 12484 5360 12540
rect 5296 12480 5360 12484
rect 5376 12540 5440 12544
rect 5376 12484 5380 12540
rect 5380 12484 5436 12540
rect 5436 12484 5440 12540
rect 5376 12480 5440 12484
rect 35856 12540 35920 12544
rect 35856 12484 35860 12540
rect 35860 12484 35916 12540
rect 35916 12484 35920 12540
rect 35856 12480 35920 12484
rect 35936 12540 36000 12544
rect 35936 12484 35940 12540
rect 35940 12484 35996 12540
rect 35996 12484 36000 12540
rect 35936 12480 36000 12484
rect 36016 12540 36080 12544
rect 36016 12484 36020 12540
rect 36020 12484 36076 12540
rect 36076 12484 36080 12540
rect 36016 12480 36080 12484
rect 36096 12540 36160 12544
rect 36096 12484 36100 12540
rect 36100 12484 36156 12540
rect 36156 12484 36160 12540
rect 36096 12480 36160 12484
rect 66576 12540 66640 12544
rect 66576 12484 66580 12540
rect 66580 12484 66636 12540
rect 66636 12484 66640 12540
rect 66576 12480 66640 12484
rect 66656 12540 66720 12544
rect 66656 12484 66660 12540
rect 66660 12484 66716 12540
rect 66716 12484 66720 12540
rect 66656 12480 66720 12484
rect 66736 12540 66800 12544
rect 66736 12484 66740 12540
rect 66740 12484 66796 12540
rect 66796 12484 66800 12540
rect 66736 12480 66800 12484
rect 66816 12540 66880 12544
rect 66816 12484 66820 12540
rect 66820 12484 66876 12540
rect 66876 12484 66880 12540
rect 66816 12480 66880 12484
rect 5796 11996 5860 12000
rect 5796 11940 5800 11996
rect 5800 11940 5856 11996
rect 5856 11940 5860 11996
rect 5796 11936 5860 11940
rect 5876 11996 5940 12000
rect 5876 11940 5880 11996
rect 5880 11940 5936 11996
rect 5936 11940 5940 11996
rect 5876 11936 5940 11940
rect 5956 11996 6020 12000
rect 5956 11940 5960 11996
rect 5960 11940 6016 11996
rect 6016 11940 6020 11996
rect 5956 11936 6020 11940
rect 6036 11996 6100 12000
rect 6036 11940 6040 11996
rect 6040 11940 6096 11996
rect 6096 11940 6100 11996
rect 6036 11936 6100 11940
rect 36516 11996 36580 12000
rect 36516 11940 36520 11996
rect 36520 11940 36576 11996
rect 36576 11940 36580 11996
rect 36516 11936 36580 11940
rect 36596 11996 36660 12000
rect 36596 11940 36600 11996
rect 36600 11940 36656 11996
rect 36656 11940 36660 11996
rect 36596 11936 36660 11940
rect 36676 11996 36740 12000
rect 36676 11940 36680 11996
rect 36680 11940 36736 11996
rect 36736 11940 36740 11996
rect 36676 11936 36740 11940
rect 36756 11996 36820 12000
rect 36756 11940 36760 11996
rect 36760 11940 36816 11996
rect 36816 11940 36820 11996
rect 36756 11936 36820 11940
rect 67236 11996 67300 12000
rect 67236 11940 67240 11996
rect 67240 11940 67296 11996
rect 67296 11940 67300 11996
rect 67236 11936 67300 11940
rect 67316 11996 67380 12000
rect 67316 11940 67320 11996
rect 67320 11940 67376 11996
rect 67376 11940 67380 11996
rect 67316 11936 67380 11940
rect 67396 11996 67460 12000
rect 67396 11940 67400 11996
rect 67400 11940 67456 11996
rect 67456 11940 67460 11996
rect 67396 11936 67460 11940
rect 67476 11996 67540 12000
rect 67476 11940 67480 11996
rect 67480 11940 67536 11996
rect 67536 11940 67540 11996
rect 67476 11936 67540 11940
rect 20668 11868 20732 11932
rect 17540 11596 17604 11660
rect 15700 11460 15764 11524
rect 5136 11452 5200 11456
rect 5136 11396 5140 11452
rect 5140 11396 5196 11452
rect 5196 11396 5200 11452
rect 5136 11392 5200 11396
rect 5216 11452 5280 11456
rect 5216 11396 5220 11452
rect 5220 11396 5276 11452
rect 5276 11396 5280 11452
rect 5216 11392 5280 11396
rect 5296 11452 5360 11456
rect 5296 11396 5300 11452
rect 5300 11396 5356 11452
rect 5356 11396 5360 11452
rect 5296 11392 5360 11396
rect 5376 11452 5440 11456
rect 5376 11396 5380 11452
rect 5380 11396 5436 11452
rect 5436 11396 5440 11452
rect 5376 11392 5440 11396
rect 35856 11452 35920 11456
rect 35856 11396 35860 11452
rect 35860 11396 35916 11452
rect 35916 11396 35920 11452
rect 35856 11392 35920 11396
rect 35936 11452 36000 11456
rect 35936 11396 35940 11452
rect 35940 11396 35996 11452
rect 35996 11396 36000 11452
rect 35936 11392 36000 11396
rect 36016 11452 36080 11456
rect 36016 11396 36020 11452
rect 36020 11396 36076 11452
rect 36076 11396 36080 11452
rect 36016 11392 36080 11396
rect 36096 11452 36160 11456
rect 36096 11396 36100 11452
rect 36100 11396 36156 11452
rect 36156 11396 36160 11452
rect 36096 11392 36160 11396
rect 66576 11452 66640 11456
rect 66576 11396 66580 11452
rect 66580 11396 66636 11452
rect 66636 11396 66640 11452
rect 66576 11392 66640 11396
rect 66656 11452 66720 11456
rect 66656 11396 66660 11452
rect 66660 11396 66716 11452
rect 66716 11396 66720 11452
rect 66656 11392 66720 11396
rect 66736 11452 66800 11456
rect 66736 11396 66740 11452
rect 66740 11396 66796 11452
rect 66796 11396 66800 11452
rect 66736 11392 66800 11396
rect 66816 11452 66880 11456
rect 66816 11396 66820 11452
rect 66820 11396 66876 11452
rect 66876 11396 66880 11452
rect 66816 11392 66880 11396
rect 11468 11324 11532 11388
rect 11652 11188 11716 11252
rect 23428 11188 23492 11252
rect 26188 11248 26252 11252
rect 26188 11192 26238 11248
rect 26238 11192 26252 11248
rect 26188 11188 26252 11192
rect 12204 11052 12268 11116
rect 24532 11052 24596 11116
rect 15884 10916 15948 10980
rect 5796 10908 5860 10912
rect 5796 10852 5800 10908
rect 5800 10852 5856 10908
rect 5856 10852 5860 10908
rect 5796 10848 5860 10852
rect 5876 10908 5940 10912
rect 5876 10852 5880 10908
rect 5880 10852 5936 10908
rect 5936 10852 5940 10908
rect 5876 10848 5940 10852
rect 5956 10908 6020 10912
rect 5956 10852 5960 10908
rect 5960 10852 6016 10908
rect 6016 10852 6020 10908
rect 5956 10848 6020 10852
rect 6036 10908 6100 10912
rect 6036 10852 6040 10908
rect 6040 10852 6096 10908
rect 6096 10852 6100 10908
rect 6036 10848 6100 10852
rect 36516 10908 36580 10912
rect 36516 10852 36520 10908
rect 36520 10852 36576 10908
rect 36576 10852 36580 10908
rect 36516 10848 36580 10852
rect 36596 10908 36660 10912
rect 36596 10852 36600 10908
rect 36600 10852 36656 10908
rect 36656 10852 36660 10908
rect 36596 10848 36660 10852
rect 36676 10908 36740 10912
rect 36676 10852 36680 10908
rect 36680 10852 36736 10908
rect 36736 10852 36740 10908
rect 36676 10848 36740 10852
rect 36756 10908 36820 10912
rect 36756 10852 36760 10908
rect 36760 10852 36816 10908
rect 36816 10852 36820 10908
rect 36756 10848 36820 10852
rect 67236 10908 67300 10912
rect 67236 10852 67240 10908
rect 67240 10852 67296 10908
rect 67296 10852 67300 10908
rect 67236 10848 67300 10852
rect 67316 10908 67380 10912
rect 67316 10852 67320 10908
rect 67320 10852 67376 10908
rect 67376 10852 67380 10908
rect 67316 10848 67380 10852
rect 67396 10908 67460 10912
rect 67396 10852 67400 10908
rect 67400 10852 67456 10908
rect 67456 10852 67460 10908
rect 67396 10848 67460 10852
rect 67476 10908 67540 10912
rect 67476 10852 67480 10908
rect 67480 10852 67536 10908
rect 67536 10852 67540 10908
rect 67476 10848 67540 10852
rect 25820 10780 25884 10844
rect 37412 10508 37476 10572
rect 8156 10372 8220 10436
rect 26004 10372 26068 10436
rect 5136 10364 5200 10368
rect 5136 10308 5140 10364
rect 5140 10308 5196 10364
rect 5196 10308 5200 10364
rect 5136 10304 5200 10308
rect 5216 10364 5280 10368
rect 5216 10308 5220 10364
rect 5220 10308 5276 10364
rect 5276 10308 5280 10364
rect 5216 10304 5280 10308
rect 5296 10364 5360 10368
rect 5296 10308 5300 10364
rect 5300 10308 5356 10364
rect 5356 10308 5360 10364
rect 5296 10304 5360 10308
rect 5376 10364 5440 10368
rect 5376 10308 5380 10364
rect 5380 10308 5436 10364
rect 5436 10308 5440 10364
rect 5376 10304 5440 10308
rect 35856 10364 35920 10368
rect 35856 10308 35860 10364
rect 35860 10308 35916 10364
rect 35916 10308 35920 10364
rect 35856 10304 35920 10308
rect 35936 10364 36000 10368
rect 35936 10308 35940 10364
rect 35940 10308 35996 10364
rect 35996 10308 36000 10364
rect 35936 10304 36000 10308
rect 36016 10364 36080 10368
rect 36016 10308 36020 10364
rect 36020 10308 36076 10364
rect 36076 10308 36080 10364
rect 36016 10304 36080 10308
rect 36096 10364 36160 10368
rect 36096 10308 36100 10364
rect 36100 10308 36156 10364
rect 36156 10308 36160 10364
rect 36096 10304 36160 10308
rect 66576 10364 66640 10368
rect 66576 10308 66580 10364
rect 66580 10308 66636 10364
rect 66636 10308 66640 10364
rect 66576 10304 66640 10308
rect 66656 10364 66720 10368
rect 66656 10308 66660 10364
rect 66660 10308 66716 10364
rect 66716 10308 66720 10364
rect 66656 10304 66720 10308
rect 66736 10364 66800 10368
rect 66736 10308 66740 10364
rect 66740 10308 66796 10364
rect 66796 10308 66800 10364
rect 66736 10304 66800 10308
rect 66816 10364 66880 10368
rect 66816 10308 66820 10364
rect 66820 10308 66876 10364
rect 66876 10308 66880 10364
rect 66816 10304 66880 10308
rect 21220 10296 21284 10300
rect 21220 10240 21234 10296
rect 21234 10240 21284 10296
rect 21220 10236 21284 10240
rect 30788 10100 30852 10164
rect 37228 10100 37292 10164
rect 10180 9964 10244 10028
rect 20852 9964 20916 10028
rect 28028 9964 28092 10028
rect 10732 9828 10796 9892
rect 5796 9820 5860 9824
rect 5796 9764 5800 9820
rect 5800 9764 5856 9820
rect 5856 9764 5860 9820
rect 5796 9760 5860 9764
rect 5876 9820 5940 9824
rect 5876 9764 5880 9820
rect 5880 9764 5936 9820
rect 5936 9764 5940 9820
rect 5876 9760 5940 9764
rect 5956 9820 6020 9824
rect 5956 9764 5960 9820
rect 5960 9764 6016 9820
rect 6016 9764 6020 9820
rect 5956 9760 6020 9764
rect 6036 9820 6100 9824
rect 6036 9764 6040 9820
rect 6040 9764 6096 9820
rect 6096 9764 6100 9820
rect 6036 9760 6100 9764
rect 19748 9692 19812 9756
rect 20484 9692 20548 9756
rect 21404 9692 21468 9756
rect 24164 9692 24228 9756
rect 26188 9692 26252 9756
rect 29132 9692 29196 9756
rect 36516 9820 36580 9824
rect 36516 9764 36520 9820
rect 36520 9764 36576 9820
rect 36576 9764 36580 9820
rect 36516 9760 36580 9764
rect 36596 9820 36660 9824
rect 36596 9764 36600 9820
rect 36600 9764 36656 9820
rect 36656 9764 36660 9820
rect 36596 9760 36660 9764
rect 36676 9820 36740 9824
rect 36676 9764 36680 9820
rect 36680 9764 36736 9820
rect 36736 9764 36740 9820
rect 36676 9760 36740 9764
rect 36756 9820 36820 9824
rect 36756 9764 36760 9820
rect 36760 9764 36816 9820
rect 36816 9764 36820 9820
rect 36756 9760 36820 9764
rect 67236 9820 67300 9824
rect 67236 9764 67240 9820
rect 67240 9764 67296 9820
rect 67296 9764 67300 9820
rect 67236 9760 67300 9764
rect 67316 9820 67380 9824
rect 67316 9764 67320 9820
rect 67320 9764 67376 9820
rect 67376 9764 67380 9820
rect 67316 9760 67380 9764
rect 67396 9820 67460 9824
rect 67396 9764 67400 9820
rect 67400 9764 67456 9820
rect 67456 9764 67460 9820
rect 67396 9760 67460 9764
rect 67476 9820 67540 9824
rect 67476 9764 67480 9820
rect 67480 9764 67536 9820
rect 67536 9764 67540 9820
rect 67476 9760 67540 9764
rect 24348 9556 24412 9620
rect 29316 9556 29380 9620
rect 29684 9556 29748 9620
rect 34284 9752 34348 9756
rect 34284 9696 34298 9752
rect 34298 9696 34348 9752
rect 34284 9692 34348 9696
rect 31156 9556 31220 9620
rect 32628 9556 32692 9620
rect 13676 9420 13740 9484
rect 30972 9420 31036 9484
rect 32444 9420 32508 9484
rect 27108 9284 27172 9348
rect 5136 9276 5200 9280
rect 5136 9220 5140 9276
rect 5140 9220 5196 9276
rect 5196 9220 5200 9276
rect 5136 9216 5200 9220
rect 5216 9276 5280 9280
rect 5216 9220 5220 9276
rect 5220 9220 5276 9276
rect 5276 9220 5280 9276
rect 5216 9216 5280 9220
rect 5296 9276 5360 9280
rect 5296 9220 5300 9276
rect 5300 9220 5356 9276
rect 5356 9220 5360 9276
rect 5296 9216 5360 9220
rect 5376 9276 5440 9280
rect 5376 9220 5380 9276
rect 5380 9220 5436 9276
rect 5436 9220 5440 9276
rect 5376 9216 5440 9220
rect 35856 9276 35920 9280
rect 35856 9220 35860 9276
rect 35860 9220 35916 9276
rect 35916 9220 35920 9276
rect 35856 9216 35920 9220
rect 35936 9276 36000 9280
rect 35936 9220 35940 9276
rect 35940 9220 35996 9276
rect 35996 9220 36000 9276
rect 35936 9216 36000 9220
rect 36016 9276 36080 9280
rect 36016 9220 36020 9276
rect 36020 9220 36076 9276
rect 36076 9220 36080 9276
rect 36016 9216 36080 9220
rect 36096 9276 36160 9280
rect 36096 9220 36100 9276
rect 36100 9220 36156 9276
rect 36156 9220 36160 9276
rect 36096 9216 36160 9220
rect 66576 9276 66640 9280
rect 66576 9220 66580 9276
rect 66580 9220 66636 9276
rect 66636 9220 66640 9276
rect 66576 9216 66640 9220
rect 66656 9276 66720 9280
rect 66656 9220 66660 9276
rect 66660 9220 66716 9276
rect 66716 9220 66720 9276
rect 66656 9216 66720 9220
rect 66736 9276 66800 9280
rect 66736 9220 66740 9276
rect 66740 9220 66796 9276
rect 66796 9220 66800 9276
rect 66736 9216 66800 9220
rect 66816 9276 66880 9280
rect 66816 9220 66820 9276
rect 66820 9220 66876 9276
rect 66876 9220 66880 9276
rect 66816 9216 66880 9220
rect 17172 9148 17236 9212
rect 19196 9208 19260 9212
rect 19196 9152 19246 9208
rect 19246 9152 19260 9208
rect 19196 9148 19260 9152
rect 27292 9148 27356 9212
rect 33916 9208 33980 9212
rect 33916 9152 33966 9208
rect 33966 9152 33980 9208
rect 33916 9148 33980 9152
rect 16804 9012 16868 9076
rect 36308 9012 36372 9076
rect 24900 8876 24964 8940
rect 27476 8876 27540 8940
rect 35204 8936 35268 8940
rect 35204 8880 35254 8936
rect 35254 8880 35268 8936
rect 35204 8876 35268 8880
rect 18092 8740 18156 8804
rect 5796 8732 5860 8736
rect 5796 8676 5800 8732
rect 5800 8676 5856 8732
rect 5856 8676 5860 8732
rect 5796 8672 5860 8676
rect 5876 8732 5940 8736
rect 5876 8676 5880 8732
rect 5880 8676 5936 8732
rect 5936 8676 5940 8732
rect 5876 8672 5940 8676
rect 5956 8732 6020 8736
rect 5956 8676 5960 8732
rect 5960 8676 6016 8732
rect 6016 8676 6020 8732
rect 5956 8672 6020 8676
rect 6036 8732 6100 8736
rect 6036 8676 6040 8732
rect 6040 8676 6096 8732
rect 6096 8676 6100 8732
rect 6036 8672 6100 8676
rect 36516 8732 36580 8736
rect 36516 8676 36520 8732
rect 36520 8676 36576 8732
rect 36576 8676 36580 8732
rect 36516 8672 36580 8676
rect 36596 8732 36660 8736
rect 36596 8676 36600 8732
rect 36600 8676 36656 8732
rect 36656 8676 36660 8732
rect 36596 8672 36660 8676
rect 36676 8732 36740 8736
rect 36676 8676 36680 8732
rect 36680 8676 36736 8732
rect 36736 8676 36740 8732
rect 36676 8672 36740 8676
rect 36756 8732 36820 8736
rect 36756 8676 36760 8732
rect 36760 8676 36816 8732
rect 36816 8676 36820 8732
rect 36756 8672 36820 8676
rect 67236 8732 67300 8736
rect 67236 8676 67240 8732
rect 67240 8676 67296 8732
rect 67296 8676 67300 8732
rect 67236 8672 67300 8676
rect 67316 8732 67380 8736
rect 67316 8676 67320 8732
rect 67320 8676 67376 8732
rect 67376 8676 67380 8732
rect 67316 8672 67380 8676
rect 67396 8732 67460 8736
rect 67396 8676 67400 8732
rect 67400 8676 67456 8732
rect 67456 8676 67460 8732
rect 67396 8672 67460 8676
rect 67476 8732 67540 8736
rect 67476 8676 67480 8732
rect 67480 8676 67536 8732
rect 67536 8676 67540 8732
rect 67476 8672 67540 8676
rect 27660 8604 27724 8668
rect 35572 8604 35636 8668
rect 20116 8468 20180 8532
rect 23060 8468 23124 8532
rect 30604 8468 30668 8532
rect 33364 8468 33428 8532
rect 9996 8332 10060 8396
rect 19564 8332 19628 8396
rect 28212 8332 28276 8396
rect 32996 8332 33060 8396
rect 34836 8332 34900 8396
rect 18276 8196 18340 8260
rect 5136 8188 5200 8192
rect 5136 8132 5140 8188
rect 5140 8132 5196 8188
rect 5196 8132 5200 8188
rect 5136 8128 5200 8132
rect 5216 8188 5280 8192
rect 5216 8132 5220 8188
rect 5220 8132 5276 8188
rect 5276 8132 5280 8188
rect 5216 8128 5280 8132
rect 5296 8188 5360 8192
rect 5296 8132 5300 8188
rect 5300 8132 5356 8188
rect 5356 8132 5360 8188
rect 5296 8128 5360 8132
rect 5376 8188 5440 8192
rect 5376 8132 5380 8188
rect 5380 8132 5436 8188
rect 5436 8132 5440 8188
rect 5376 8128 5440 8132
rect 35856 8188 35920 8192
rect 35856 8132 35860 8188
rect 35860 8132 35916 8188
rect 35916 8132 35920 8188
rect 35856 8128 35920 8132
rect 35936 8188 36000 8192
rect 35936 8132 35940 8188
rect 35940 8132 35996 8188
rect 35996 8132 36000 8188
rect 35936 8128 36000 8132
rect 36016 8188 36080 8192
rect 36016 8132 36020 8188
rect 36020 8132 36076 8188
rect 36076 8132 36080 8188
rect 36016 8128 36080 8132
rect 36096 8188 36160 8192
rect 36096 8132 36100 8188
rect 36100 8132 36156 8188
rect 36156 8132 36160 8188
rect 36096 8128 36160 8132
rect 66576 8188 66640 8192
rect 66576 8132 66580 8188
rect 66580 8132 66636 8188
rect 66636 8132 66640 8188
rect 66576 8128 66640 8132
rect 66656 8188 66720 8192
rect 66656 8132 66660 8188
rect 66660 8132 66716 8188
rect 66716 8132 66720 8188
rect 66656 8128 66720 8132
rect 66736 8188 66800 8192
rect 66736 8132 66740 8188
rect 66740 8132 66796 8188
rect 66796 8132 66800 8188
rect 66736 8128 66800 8132
rect 66816 8188 66880 8192
rect 66816 8132 66820 8188
rect 66820 8132 66876 8188
rect 66876 8132 66880 8188
rect 66816 8128 66880 8132
rect 22508 8060 22572 8124
rect 24348 8060 24412 8124
rect 33180 8060 33244 8124
rect 14964 7848 15028 7852
rect 14964 7792 15014 7848
rect 15014 7792 15028 7848
rect 14964 7788 15028 7792
rect 25084 7788 25148 7852
rect 41460 7788 41524 7852
rect 5796 7644 5860 7648
rect 5796 7588 5800 7644
rect 5800 7588 5856 7644
rect 5856 7588 5860 7644
rect 5796 7584 5860 7588
rect 5876 7644 5940 7648
rect 5876 7588 5880 7644
rect 5880 7588 5936 7644
rect 5936 7588 5940 7644
rect 5876 7584 5940 7588
rect 5956 7644 6020 7648
rect 5956 7588 5960 7644
rect 5960 7588 6016 7644
rect 6016 7588 6020 7644
rect 5956 7584 6020 7588
rect 6036 7644 6100 7648
rect 6036 7588 6040 7644
rect 6040 7588 6096 7644
rect 6096 7588 6100 7644
rect 6036 7584 6100 7588
rect 17908 7516 17972 7580
rect 22508 7516 22572 7580
rect 36516 7644 36580 7648
rect 36516 7588 36520 7644
rect 36520 7588 36576 7644
rect 36576 7588 36580 7644
rect 36516 7584 36580 7588
rect 36596 7644 36660 7648
rect 36596 7588 36600 7644
rect 36600 7588 36656 7644
rect 36656 7588 36660 7644
rect 36596 7584 36660 7588
rect 36676 7644 36740 7648
rect 36676 7588 36680 7644
rect 36680 7588 36736 7644
rect 36736 7588 36740 7644
rect 36676 7584 36740 7588
rect 36756 7644 36820 7648
rect 36756 7588 36760 7644
rect 36760 7588 36816 7644
rect 36816 7588 36820 7644
rect 36756 7584 36820 7588
rect 67236 7644 67300 7648
rect 67236 7588 67240 7644
rect 67240 7588 67296 7644
rect 67296 7588 67300 7644
rect 67236 7584 67300 7588
rect 67316 7644 67380 7648
rect 67316 7588 67320 7644
rect 67320 7588 67376 7644
rect 67376 7588 67380 7644
rect 67316 7584 67380 7588
rect 67396 7644 67460 7648
rect 67396 7588 67400 7644
rect 67400 7588 67456 7644
rect 67456 7588 67460 7644
rect 67396 7584 67460 7588
rect 67476 7644 67540 7648
rect 67476 7588 67480 7644
rect 67480 7588 67536 7644
rect 67536 7588 67540 7644
rect 67476 7584 67540 7588
rect 31524 7516 31588 7580
rect 35388 7516 35452 7580
rect 25820 7380 25884 7444
rect 32812 7380 32876 7444
rect 26004 7108 26068 7172
rect 28212 7108 28276 7172
rect 33916 7168 33980 7172
rect 33916 7112 33930 7168
rect 33930 7112 33980 7168
rect 33916 7108 33980 7112
rect 5136 7100 5200 7104
rect 5136 7044 5140 7100
rect 5140 7044 5196 7100
rect 5196 7044 5200 7100
rect 5136 7040 5200 7044
rect 5216 7100 5280 7104
rect 5216 7044 5220 7100
rect 5220 7044 5276 7100
rect 5276 7044 5280 7100
rect 5216 7040 5280 7044
rect 5296 7100 5360 7104
rect 5296 7044 5300 7100
rect 5300 7044 5356 7100
rect 5356 7044 5360 7100
rect 5296 7040 5360 7044
rect 5376 7100 5440 7104
rect 5376 7044 5380 7100
rect 5380 7044 5436 7100
rect 5436 7044 5440 7100
rect 5376 7040 5440 7044
rect 35856 7100 35920 7104
rect 35856 7044 35860 7100
rect 35860 7044 35916 7100
rect 35916 7044 35920 7100
rect 35856 7040 35920 7044
rect 35936 7100 36000 7104
rect 35936 7044 35940 7100
rect 35940 7044 35996 7100
rect 35996 7044 36000 7100
rect 35936 7040 36000 7044
rect 36016 7100 36080 7104
rect 36016 7044 36020 7100
rect 36020 7044 36076 7100
rect 36076 7044 36080 7100
rect 36016 7040 36080 7044
rect 36096 7100 36160 7104
rect 36096 7044 36100 7100
rect 36100 7044 36156 7100
rect 36156 7044 36160 7100
rect 36096 7040 36160 7044
rect 66576 7100 66640 7104
rect 66576 7044 66580 7100
rect 66580 7044 66636 7100
rect 66636 7044 66640 7100
rect 66576 7040 66640 7044
rect 66656 7100 66720 7104
rect 66656 7044 66660 7100
rect 66660 7044 66716 7100
rect 66716 7044 66720 7100
rect 66656 7040 66720 7044
rect 66736 7100 66800 7104
rect 66736 7044 66740 7100
rect 66740 7044 66796 7100
rect 66796 7044 66800 7100
rect 66736 7040 66800 7044
rect 66816 7100 66880 7104
rect 66816 7044 66820 7100
rect 66820 7044 66876 7100
rect 66876 7044 66880 7100
rect 66816 7040 66880 7044
rect 15148 6972 15212 7036
rect 22508 6896 22572 6900
rect 22508 6840 22558 6896
rect 22558 6840 22572 6896
rect 22508 6836 22572 6840
rect 27292 6836 27356 6900
rect 25636 6700 25700 6764
rect 32628 6700 32692 6764
rect 5796 6556 5860 6560
rect 5796 6500 5800 6556
rect 5800 6500 5856 6556
rect 5856 6500 5860 6556
rect 5796 6496 5860 6500
rect 5876 6556 5940 6560
rect 5876 6500 5880 6556
rect 5880 6500 5936 6556
rect 5936 6500 5940 6556
rect 5876 6496 5940 6500
rect 5956 6556 6020 6560
rect 5956 6500 5960 6556
rect 5960 6500 6016 6556
rect 6016 6500 6020 6556
rect 5956 6496 6020 6500
rect 6036 6556 6100 6560
rect 6036 6500 6040 6556
rect 6040 6500 6096 6556
rect 6096 6500 6100 6556
rect 6036 6496 6100 6500
rect 29316 6564 29380 6628
rect 36516 6556 36580 6560
rect 36516 6500 36520 6556
rect 36520 6500 36576 6556
rect 36576 6500 36580 6556
rect 36516 6496 36580 6500
rect 36596 6556 36660 6560
rect 36596 6500 36600 6556
rect 36600 6500 36656 6556
rect 36656 6500 36660 6556
rect 36596 6496 36660 6500
rect 36676 6556 36740 6560
rect 36676 6500 36680 6556
rect 36680 6500 36736 6556
rect 36736 6500 36740 6556
rect 36676 6496 36740 6500
rect 36756 6556 36820 6560
rect 36756 6500 36760 6556
rect 36760 6500 36816 6556
rect 36816 6500 36820 6556
rect 36756 6496 36820 6500
rect 67236 6556 67300 6560
rect 67236 6500 67240 6556
rect 67240 6500 67296 6556
rect 67296 6500 67300 6556
rect 67236 6496 67300 6500
rect 67316 6556 67380 6560
rect 67316 6500 67320 6556
rect 67320 6500 67376 6556
rect 67376 6500 67380 6556
rect 67316 6496 67380 6500
rect 67396 6556 67460 6560
rect 67396 6500 67400 6556
rect 67400 6500 67456 6556
rect 67456 6500 67460 6556
rect 67396 6496 67460 6500
rect 67476 6556 67540 6560
rect 67476 6500 67480 6556
rect 67480 6500 67536 6556
rect 67536 6500 67540 6556
rect 67476 6496 67540 6500
rect 14596 6292 14660 6356
rect 24532 6428 24596 6492
rect 31156 6428 31220 6492
rect 21220 6156 21284 6220
rect 5136 6012 5200 6016
rect 5136 5956 5140 6012
rect 5140 5956 5196 6012
rect 5196 5956 5200 6012
rect 5136 5952 5200 5956
rect 5216 6012 5280 6016
rect 5216 5956 5220 6012
rect 5220 5956 5276 6012
rect 5276 5956 5280 6012
rect 5216 5952 5280 5956
rect 5296 6012 5360 6016
rect 5296 5956 5300 6012
rect 5300 5956 5356 6012
rect 5356 5956 5360 6012
rect 5296 5952 5360 5956
rect 5376 6012 5440 6016
rect 5376 5956 5380 6012
rect 5380 5956 5436 6012
rect 5436 5956 5440 6012
rect 5376 5952 5440 5956
rect 35856 6012 35920 6016
rect 35856 5956 35860 6012
rect 35860 5956 35916 6012
rect 35916 5956 35920 6012
rect 35856 5952 35920 5956
rect 35936 6012 36000 6016
rect 35936 5956 35940 6012
rect 35940 5956 35996 6012
rect 35996 5956 36000 6012
rect 35936 5952 36000 5956
rect 36016 6012 36080 6016
rect 36016 5956 36020 6012
rect 36020 5956 36076 6012
rect 36076 5956 36080 6012
rect 36016 5952 36080 5956
rect 36096 6012 36160 6016
rect 36096 5956 36100 6012
rect 36100 5956 36156 6012
rect 36156 5956 36160 6012
rect 36096 5952 36160 5956
rect 66576 6012 66640 6016
rect 66576 5956 66580 6012
rect 66580 5956 66636 6012
rect 66636 5956 66640 6012
rect 66576 5952 66640 5956
rect 66656 6012 66720 6016
rect 66656 5956 66660 6012
rect 66660 5956 66716 6012
rect 66716 5956 66720 6012
rect 66656 5952 66720 5956
rect 66736 6012 66800 6016
rect 66736 5956 66740 6012
rect 66740 5956 66796 6012
rect 66796 5956 66800 6012
rect 66736 5952 66800 5956
rect 66816 6012 66880 6016
rect 66816 5956 66820 6012
rect 66820 5956 66876 6012
rect 66876 5956 66880 6012
rect 66816 5952 66880 5956
rect 26924 5884 26988 5948
rect 27476 5748 27540 5812
rect 19196 5672 19260 5676
rect 19196 5616 19246 5672
rect 19246 5616 19260 5672
rect 19196 5612 19260 5616
rect 20852 5672 20916 5676
rect 20852 5616 20866 5672
rect 20866 5616 20916 5672
rect 20852 5612 20916 5616
rect 23060 5672 23124 5676
rect 23060 5616 23074 5672
rect 23074 5616 23124 5672
rect 23060 5612 23124 5616
rect 24164 5672 24228 5676
rect 24164 5616 24178 5672
rect 24178 5616 24228 5672
rect 24164 5612 24228 5616
rect 25084 5672 25148 5676
rect 25084 5616 25134 5672
rect 25134 5616 25148 5672
rect 25084 5612 25148 5616
rect 29132 5612 29196 5676
rect 15700 5476 15764 5540
rect 31524 5748 31588 5812
rect 35388 5536 35452 5540
rect 35388 5480 35438 5536
rect 35438 5480 35452 5536
rect 35388 5476 35452 5480
rect 5796 5468 5860 5472
rect 5796 5412 5800 5468
rect 5800 5412 5856 5468
rect 5856 5412 5860 5468
rect 5796 5408 5860 5412
rect 5876 5468 5940 5472
rect 5876 5412 5880 5468
rect 5880 5412 5936 5468
rect 5936 5412 5940 5468
rect 5876 5408 5940 5412
rect 5956 5468 6020 5472
rect 5956 5412 5960 5468
rect 5960 5412 6016 5468
rect 6016 5412 6020 5468
rect 5956 5408 6020 5412
rect 6036 5468 6100 5472
rect 6036 5412 6040 5468
rect 6040 5412 6096 5468
rect 6096 5412 6100 5468
rect 6036 5408 6100 5412
rect 36516 5468 36580 5472
rect 36516 5412 36520 5468
rect 36520 5412 36576 5468
rect 36576 5412 36580 5468
rect 36516 5408 36580 5412
rect 36596 5468 36660 5472
rect 36596 5412 36600 5468
rect 36600 5412 36656 5468
rect 36656 5412 36660 5468
rect 36596 5408 36660 5412
rect 36676 5468 36740 5472
rect 36676 5412 36680 5468
rect 36680 5412 36736 5468
rect 36736 5412 36740 5468
rect 36676 5408 36740 5412
rect 36756 5468 36820 5472
rect 36756 5412 36760 5468
rect 36760 5412 36816 5468
rect 36816 5412 36820 5468
rect 36756 5408 36820 5412
rect 67236 5468 67300 5472
rect 67236 5412 67240 5468
rect 67240 5412 67296 5468
rect 67296 5412 67300 5468
rect 67236 5408 67300 5412
rect 67316 5468 67380 5472
rect 67316 5412 67320 5468
rect 67320 5412 67376 5468
rect 67376 5412 67380 5468
rect 67316 5408 67380 5412
rect 67396 5468 67460 5472
rect 67396 5412 67400 5468
rect 67400 5412 67456 5468
rect 67456 5412 67460 5468
rect 67396 5408 67460 5412
rect 67476 5468 67540 5472
rect 67476 5412 67480 5468
rect 67480 5412 67536 5468
rect 67536 5412 67540 5468
rect 67476 5408 67540 5412
rect 17908 5340 17972 5404
rect 32444 5340 32508 5404
rect 27660 5204 27724 5268
rect 30604 5204 30668 5268
rect 14780 5068 14844 5132
rect 34836 5128 34900 5132
rect 34836 5072 34850 5128
rect 34850 5072 34900 5128
rect 34836 5068 34900 5072
rect 35572 5068 35636 5132
rect 40356 5068 40420 5132
rect 5136 4924 5200 4928
rect 5136 4868 5140 4924
rect 5140 4868 5196 4924
rect 5196 4868 5200 4924
rect 5136 4864 5200 4868
rect 5216 4924 5280 4928
rect 5216 4868 5220 4924
rect 5220 4868 5276 4924
rect 5276 4868 5280 4924
rect 5216 4864 5280 4868
rect 5296 4924 5360 4928
rect 5296 4868 5300 4924
rect 5300 4868 5356 4924
rect 5356 4868 5360 4924
rect 5296 4864 5360 4868
rect 5376 4924 5440 4928
rect 5376 4868 5380 4924
rect 5380 4868 5436 4924
rect 5436 4868 5440 4924
rect 5376 4864 5440 4868
rect 35856 4924 35920 4928
rect 35856 4868 35860 4924
rect 35860 4868 35916 4924
rect 35916 4868 35920 4924
rect 35856 4864 35920 4868
rect 35936 4924 36000 4928
rect 35936 4868 35940 4924
rect 35940 4868 35996 4924
rect 35996 4868 36000 4924
rect 35936 4864 36000 4868
rect 36016 4924 36080 4928
rect 36016 4868 36020 4924
rect 36020 4868 36076 4924
rect 36076 4868 36080 4924
rect 36016 4864 36080 4868
rect 36096 4924 36160 4928
rect 36096 4868 36100 4924
rect 36100 4868 36156 4924
rect 36156 4868 36160 4924
rect 36096 4864 36160 4868
rect 66576 4924 66640 4928
rect 66576 4868 66580 4924
rect 66580 4868 66636 4924
rect 66636 4868 66640 4924
rect 66576 4864 66640 4868
rect 66656 4924 66720 4928
rect 66656 4868 66660 4924
rect 66660 4868 66716 4924
rect 66716 4868 66720 4924
rect 66656 4864 66720 4868
rect 66736 4924 66800 4928
rect 66736 4868 66740 4924
rect 66740 4868 66796 4924
rect 66796 4868 66800 4924
rect 66736 4864 66800 4868
rect 66816 4924 66880 4928
rect 66816 4868 66820 4924
rect 66820 4868 66876 4924
rect 66876 4868 66880 4924
rect 66816 4864 66880 4868
rect 30972 4796 31036 4860
rect 10732 4660 10796 4724
rect 11468 4660 11532 4724
rect 12204 4660 12268 4724
rect 13676 4660 13740 4724
rect 5796 4380 5860 4384
rect 5796 4324 5800 4380
rect 5800 4324 5856 4380
rect 5856 4324 5860 4380
rect 5796 4320 5860 4324
rect 5876 4380 5940 4384
rect 5876 4324 5880 4380
rect 5880 4324 5936 4380
rect 5936 4324 5940 4380
rect 5876 4320 5940 4324
rect 5956 4380 6020 4384
rect 5956 4324 5960 4380
rect 5960 4324 6016 4380
rect 6016 4324 6020 4380
rect 5956 4320 6020 4324
rect 6036 4380 6100 4384
rect 6036 4324 6040 4380
rect 6040 4324 6096 4380
rect 6096 4324 6100 4380
rect 6036 4320 6100 4324
rect 17540 4252 17604 4316
rect 23428 4660 23492 4724
rect 28028 4584 28092 4588
rect 28028 4528 28042 4584
rect 28042 4528 28092 4584
rect 28028 4524 28092 4528
rect 28948 4584 29012 4588
rect 28948 4528 28998 4584
rect 28998 4528 29012 4584
rect 28948 4524 29012 4528
rect 26924 4388 26988 4452
rect 35572 4388 35636 4452
rect 36516 4380 36580 4384
rect 36516 4324 36520 4380
rect 36520 4324 36576 4380
rect 36576 4324 36580 4380
rect 36516 4320 36580 4324
rect 36596 4380 36660 4384
rect 36596 4324 36600 4380
rect 36600 4324 36656 4380
rect 36656 4324 36660 4380
rect 36596 4320 36660 4324
rect 36676 4380 36740 4384
rect 36676 4324 36680 4380
rect 36680 4324 36736 4380
rect 36736 4324 36740 4380
rect 36676 4320 36740 4324
rect 36756 4380 36820 4384
rect 36756 4324 36760 4380
rect 36760 4324 36816 4380
rect 36816 4324 36820 4380
rect 36756 4320 36820 4324
rect 67236 4380 67300 4384
rect 67236 4324 67240 4380
rect 67240 4324 67296 4380
rect 67296 4324 67300 4380
rect 67236 4320 67300 4324
rect 67316 4380 67380 4384
rect 67316 4324 67320 4380
rect 67320 4324 67376 4380
rect 67376 4324 67380 4380
rect 67316 4320 67380 4324
rect 67396 4380 67460 4384
rect 67396 4324 67400 4380
rect 67400 4324 67456 4380
rect 67456 4324 67460 4380
rect 67396 4320 67460 4324
rect 67476 4380 67540 4384
rect 67476 4324 67480 4380
rect 67480 4324 67536 4380
rect 67536 4324 67540 4380
rect 67476 4320 67540 4324
rect 24900 4116 24964 4180
rect 10180 3980 10244 4044
rect 16804 4040 16868 4044
rect 16804 3984 16818 4040
rect 16818 3984 16868 4040
rect 16804 3980 16868 3984
rect 20668 3980 20732 4044
rect 21404 4040 21468 4044
rect 21404 3984 21418 4040
rect 21418 3984 21468 4040
rect 21404 3980 21468 3984
rect 15884 3844 15948 3908
rect 5136 3836 5200 3840
rect 5136 3780 5140 3836
rect 5140 3780 5196 3836
rect 5196 3780 5200 3836
rect 5136 3776 5200 3780
rect 5216 3836 5280 3840
rect 5216 3780 5220 3836
rect 5220 3780 5276 3836
rect 5276 3780 5280 3836
rect 5216 3776 5280 3780
rect 5296 3836 5360 3840
rect 5296 3780 5300 3836
rect 5300 3780 5356 3836
rect 5356 3780 5360 3836
rect 5296 3776 5360 3780
rect 5376 3836 5440 3840
rect 5376 3780 5380 3836
rect 5380 3780 5436 3836
rect 5436 3780 5440 3836
rect 5376 3776 5440 3780
rect 11652 3708 11716 3772
rect 18276 3708 18340 3772
rect 20484 3708 20548 3772
rect 14228 3572 14292 3636
rect 14964 3572 15028 3636
rect 26188 3904 26252 3908
rect 26188 3848 26202 3904
rect 26202 3848 26252 3904
rect 25636 3768 25700 3772
rect 25636 3712 25650 3768
rect 25650 3712 25700 3768
rect 25636 3708 25700 3712
rect 26188 3844 26252 3848
rect 35856 3836 35920 3840
rect 35856 3780 35860 3836
rect 35860 3780 35916 3836
rect 35916 3780 35920 3836
rect 35856 3776 35920 3780
rect 35936 3836 36000 3840
rect 35936 3780 35940 3836
rect 35940 3780 35996 3836
rect 35996 3780 36000 3836
rect 35936 3776 36000 3780
rect 36016 3836 36080 3840
rect 36016 3780 36020 3836
rect 36020 3780 36076 3836
rect 36076 3780 36080 3836
rect 36016 3776 36080 3780
rect 36096 3836 36160 3840
rect 36096 3780 36100 3836
rect 36100 3780 36156 3836
rect 36156 3780 36160 3836
rect 36096 3776 36160 3780
rect 66576 3836 66640 3840
rect 66576 3780 66580 3836
rect 66580 3780 66636 3836
rect 66636 3780 66640 3836
rect 66576 3776 66640 3780
rect 66656 3836 66720 3840
rect 66656 3780 66660 3836
rect 66660 3780 66716 3836
rect 66716 3780 66720 3836
rect 66656 3776 66720 3780
rect 66736 3836 66800 3840
rect 66736 3780 66740 3836
rect 66740 3780 66796 3836
rect 66796 3780 66800 3836
rect 66736 3776 66800 3780
rect 66816 3836 66880 3840
rect 66816 3780 66820 3836
rect 66820 3780 66876 3836
rect 66876 3780 66880 3836
rect 66816 3776 66880 3780
rect 17172 3300 17236 3364
rect 26924 3360 26988 3364
rect 26924 3304 26974 3360
rect 26974 3304 26988 3360
rect 26924 3300 26988 3304
rect 32812 3300 32876 3364
rect 35204 3300 35268 3364
rect 5796 3292 5860 3296
rect 5796 3236 5800 3292
rect 5800 3236 5856 3292
rect 5856 3236 5860 3292
rect 5796 3232 5860 3236
rect 5876 3292 5940 3296
rect 5876 3236 5880 3292
rect 5880 3236 5936 3292
rect 5936 3236 5940 3292
rect 5876 3232 5940 3236
rect 5956 3292 6020 3296
rect 5956 3236 5960 3292
rect 5960 3236 6016 3292
rect 6016 3236 6020 3292
rect 5956 3232 6020 3236
rect 6036 3292 6100 3296
rect 6036 3236 6040 3292
rect 6040 3236 6096 3292
rect 6096 3236 6100 3292
rect 6036 3232 6100 3236
rect 36516 3292 36580 3296
rect 36516 3236 36520 3292
rect 36520 3236 36576 3292
rect 36576 3236 36580 3292
rect 36516 3232 36580 3236
rect 36596 3292 36660 3296
rect 36596 3236 36600 3292
rect 36600 3236 36656 3292
rect 36656 3236 36660 3292
rect 36596 3232 36660 3236
rect 36676 3292 36740 3296
rect 36676 3236 36680 3292
rect 36680 3236 36736 3292
rect 36736 3236 36740 3292
rect 36676 3232 36740 3236
rect 36756 3292 36820 3296
rect 36756 3236 36760 3292
rect 36760 3236 36816 3292
rect 36816 3236 36820 3292
rect 36756 3232 36820 3236
rect 67236 3292 67300 3296
rect 67236 3236 67240 3292
rect 67240 3236 67296 3292
rect 67296 3236 67300 3292
rect 67236 3232 67300 3236
rect 67316 3292 67380 3296
rect 67316 3236 67320 3292
rect 67320 3236 67376 3292
rect 67376 3236 67380 3292
rect 67316 3232 67380 3236
rect 67396 3292 67460 3296
rect 67396 3236 67400 3292
rect 67400 3236 67456 3292
rect 67456 3236 67460 3292
rect 67396 3232 67460 3236
rect 67476 3292 67540 3296
rect 67476 3236 67480 3292
rect 67480 3236 67536 3292
rect 67536 3236 67540 3292
rect 67476 3232 67540 3236
rect 8156 3224 8220 3228
rect 8156 3168 8206 3224
rect 8206 3168 8220 3224
rect 8156 3164 8220 3168
rect 33364 3164 33428 3228
rect 9996 3088 10060 3092
rect 9996 3032 10010 3088
rect 10010 3032 10060 3088
rect 9996 3028 10060 3032
rect 37412 3028 37476 3092
rect 27108 2892 27172 2956
rect 32996 2952 33060 2956
rect 32996 2896 33046 2952
rect 33046 2896 33060 2952
rect 32996 2892 33060 2896
rect 5136 2748 5200 2752
rect 5136 2692 5140 2748
rect 5140 2692 5196 2748
rect 5196 2692 5200 2748
rect 5136 2688 5200 2692
rect 5216 2748 5280 2752
rect 5216 2692 5220 2748
rect 5220 2692 5276 2748
rect 5276 2692 5280 2748
rect 5216 2688 5280 2692
rect 5296 2748 5360 2752
rect 5296 2692 5300 2748
rect 5300 2692 5356 2748
rect 5356 2692 5360 2748
rect 5296 2688 5360 2692
rect 5376 2748 5440 2752
rect 5376 2692 5380 2748
rect 5380 2692 5436 2748
rect 5436 2692 5440 2748
rect 5376 2688 5440 2692
rect 15148 2620 15212 2684
rect 35856 2748 35920 2752
rect 35856 2692 35860 2748
rect 35860 2692 35916 2748
rect 35916 2692 35920 2748
rect 35856 2688 35920 2692
rect 35936 2748 36000 2752
rect 35936 2692 35940 2748
rect 35940 2692 35996 2748
rect 35996 2692 36000 2748
rect 35936 2688 36000 2692
rect 36016 2748 36080 2752
rect 36016 2692 36020 2748
rect 36020 2692 36076 2748
rect 36076 2692 36080 2748
rect 36016 2688 36080 2692
rect 36096 2748 36160 2752
rect 36096 2692 36100 2748
rect 36100 2692 36156 2748
rect 36156 2692 36160 2748
rect 36096 2688 36160 2692
rect 66576 2748 66640 2752
rect 66576 2692 66580 2748
rect 66580 2692 66636 2748
rect 66636 2692 66640 2748
rect 66576 2688 66640 2692
rect 66656 2748 66720 2752
rect 66656 2692 66660 2748
rect 66660 2692 66716 2748
rect 66716 2692 66720 2748
rect 66656 2688 66720 2692
rect 66736 2748 66800 2752
rect 66736 2692 66740 2748
rect 66740 2692 66796 2748
rect 66796 2692 66800 2748
rect 66736 2688 66800 2692
rect 66816 2748 66880 2752
rect 66816 2692 66820 2748
rect 66820 2692 66876 2748
rect 66876 2692 66880 2748
rect 66816 2688 66880 2692
rect 22508 2620 22572 2684
rect 19748 2484 19812 2548
rect 37228 2484 37292 2548
rect 19564 2348 19628 2412
rect 36308 2348 36372 2412
rect 18092 2212 18156 2276
rect 29684 2212 29748 2276
rect 5796 2204 5860 2208
rect 5796 2148 5800 2204
rect 5800 2148 5856 2204
rect 5856 2148 5860 2204
rect 5796 2144 5860 2148
rect 5876 2204 5940 2208
rect 5876 2148 5880 2204
rect 5880 2148 5936 2204
rect 5936 2148 5940 2204
rect 5876 2144 5940 2148
rect 5956 2204 6020 2208
rect 5956 2148 5960 2204
rect 5960 2148 6016 2204
rect 6016 2148 6020 2204
rect 5956 2144 6020 2148
rect 6036 2204 6100 2208
rect 6036 2148 6040 2204
rect 6040 2148 6096 2204
rect 6096 2148 6100 2204
rect 6036 2144 6100 2148
rect 36516 2204 36580 2208
rect 36516 2148 36520 2204
rect 36520 2148 36576 2204
rect 36576 2148 36580 2204
rect 36516 2144 36580 2148
rect 36596 2204 36660 2208
rect 36596 2148 36600 2204
rect 36600 2148 36656 2204
rect 36656 2148 36660 2204
rect 36596 2144 36660 2148
rect 36676 2204 36740 2208
rect 36676 2148 36680 2204
rect 36680 2148 36736 2204
rect 36736 2148 36740 2204
rect 36676 2144 36740 2148
rect 36756 2204 36820 2208
rect 36756 2148 36760 2204
rect 36760 2148 36816 2204
rect 36816 2148 36820 2204
rect 36756 2144 36820 2148
rect 67236 2204 67300 2208
rect 67236 2148 67240 2204
rect 67240 2148 67296 2204
rect 67296 2148 67300 2204
rect 67236 2144 67300 2148
rect 67316 2204 67380 2208
rect 67316 2148 67320 2204
rect 67320 2148 67376 2204
rect 67376 2148 67380 2204
rect 67316 2144 67380 2148
rect 67396 2204 67460 2208
rect 67396 2148 67400 2204
rect 67400 2148 67456 2204
rect 67456 2148 67460 2204
rect 67396 2144 67460 2148
rect 67476 2204 67540 2208
rect 67476 2148 67480 2204
rect 67480 2148 67536 2204
rect 67536 2148 67540 2204
rect 67476 2144 67540 2148
rect 24900 2076 24964 2140
rect 34284 2076 34348 2140
rect 18276 1804 18340 1868
rect 30788 1532 30852 1596
rect 31524 1260 31588 1324
rect 14780 172 14844 236
rect 28948 36 29012 100
<< metal4 >>
rect 5128 37568 5448 37584
rect 5128 37504 5136 37568
rect 5200 37504 5216 37568
rect 5280 37504 5296 37568
rect 5360 37504 5376 37568
rect 5440 37504 5448 37568
rect 5128 36480 5448 37504
rect 5128 36416 5136 36480
rect 5200 36416 5216 36480
rect 5280 36416 5296 36480
rect 5360 36416 5376 36480
rect 5440 36416 5448 36480
rect 5128 35392 5448 36416
rect 5128 35328 5136 35392
rect 5200 35328 5216 35392
rect 5280 35328 5296 35392
rect 5360 35328 5376 35392
rect 5440 35328 5448 35392
rect 5128 34304 5448 35328
rect 5128 34240 5136 34304
rect 5200 34240 5216 34304
rect 5280 34240 5296 34304
rect 5360 34240 5376 34304
rect 5440 34240 5448 34304
rect 5128 33216 5448 34240
rect 5128 33152 5136 33216
rect 5200 33152 5216 33216
rect 5280 33152 5296 33216
rect 5360 33152 5376 33216
rect 5440 33152 5448 33216
rect 5128 32128 5448 33152
rect 5128 32064 5136 32128
rect 5200 32064 5216 32128
rect 5280 32064 5296 32128
rect 5360 32064 5376 32128
rect 5440 32064 5448 32128
rect 5128 31040 5448 32064
rect 5128 30976 5136 31040
rect 5200 30976 5216 31040
rect 5280 30976 5296 31040
rect 5360 30976 5376 31040
rect 5440 30976 5448 31040
rect 5128 29952 5448 30976
rect 5128 29888 5136 29952
rect 5200 29888 5216 29952
rect 5280 29888 5296 29952
rect 5360 29888 5376 29952
rect 5440 29888 5448 29952
rect 5128 28864 5448 29888
rect 5128 28800 5136 28864
rect 5200 28800 5216 28864
rect 5280 28800 5296 28864
rect 5360 28800 5376 28864
rect 5440 28800 5448 28864
rect 5128 27776 5448 28800
rect 5128 27712 5136 27776
rect 5200 27712 5216 27776
rect 5280 27712 5296 27776
rect 5360 27712 5376 27776
rect 5440 27712 5448 27776
rect 5128 26688 5448 27712
rect 5128 26624 5136 26688
rect 5200 26624 5216 26688
rect 5280 26624 5296 26688
rect 5360 26624 5376 26688
rect 5440 26624 5448 26688
rect 5128 25600 5448 26624
rect 5128 25536 5136 25600
rect 5200 25536 5216 25600
rect 5280 25536 5296 25600
rect 5360 25536 5376 25600
rect 5440 25536 5448 25600
rect 5128 24512 5448 25536
rect 5128 24448 5136 24512
rect 5200 24448 5216 24512
rect 5280 24448 5296 24512
rect 5360 24448 5376 24512
rect 5440 24448 5448 24512
rect 5128 23424 5448 24448
rect 5128 23360 5136 23424
rect 5200 23360 5216 23424
rect 5280 23360 5296 23424
rect 5360 23360 5376 23424
rect 5440 23360 5448 23424
rect 5128 22336 5448 23360
rect 5128 22272 5136 22336
rect 5200 22272 5216 22336
rect 5280 22272 5296 22336
rect 5360 22272 5376 22336
rect 5440 22272 5448 22336
rect 5128 21248 5448 22272
rect 5128 21184 5136 21248
rect 5200 21184 5216 21248
rect 5280 21184 5296 21248
rect 5360 21184 5376 21248
rect 5440 21184 5448 21248
rect 5128 20160 5448 21184
rect 5128 20096 5136 20160
rect 5200 20096 5216 20160
rect 5280 20096 5296 20160
rect 5360 20096 5376 20160
rect 5440 20096 5448 20160
rect 5128 19072 5448 20096
rect 5128 19008 5136 19072
rect 5200 19008 5216 19072
rect 5280 19008 5296 19072
rect 5360 19008 5376 19072
rect 5440 19008 5448 19072
rect 5128 17984 5448 19008
rect 5128 17920 5136 17984
rect 5200 17920 5216 17984
rect 5280 17920 5296 17984
rect 5360 17920 5376 17984
rect 5440 17920 5448 17984
rect 5128 16896 5448 17920
rect 5128 16832 5136 16896
rect 5200 16832 5216 16896
rect 5280 16832 5296 16896
rect 5360 16832 5376 16896
rect 5440 16832 5448 16896
rect 5128 15808 5448 16832
rect 5128 15744 5136 15808
rect 5200 15744 5216 15808
rect 5280 15744 5296 15808
rect 5360 15744 5376 15808
rect 5440 15744 5448 15808
rect 5128 14720 5448 15744
rect 5128 14656 5136 14720
rect 5200 14656 5216 14720
rect 5280 14656 5296 14720
rect 5360 14656 5376 14720
rect 5440 14656 5448 14720
rect 5128 13632 5448 14656
rect 5128 13568 5136 13632
rect 5200 13568 5216 13632
rect 5280 13568 5296 13632
rect 5360 13568 5376 13632
rect 5440 13568 5448 13632
rect 5128 12544 5448 13568
rect 5128 12480 5136 12544
rect 5200 12480 5216 12544
rect 5280 12480 5296 12544
rect 5360 12480 5376 12544
rect 5440 12480 5448 12544
rect 5128 11456 5448 12480
rect 5128 11392 5136 11456
rect 5200 11392 5216 11456
rect 5280 11392 5296 11456
rect 5360 11392 5376 11456
rect 5440 11392 5448 11456
rect 5128 10368 5448 11392
rect 5128 10304 5136 10368
rect 5200 10304 5216 10368
rect 5280 10304 5296 10368
rect 5360 10304 5376 10368
rect 5440 10304 5448 10368
rect 5128 9280 5448 10304
rect 5128 9216 5136 9280
rect 5200 9216 5216 9280
rect 5280 9216 5296 9280
rect 5360 9216 5376 9280
rect 5440 9216 5448 9280
rect 5128 8192 5448 9216
rect 5128 8128 5136 8192
rect 5200 8128 5216 8192
rect 5280 8128 5296 8192
rect 5360 8128 5376 8192
rect 5440 8128 5448 8192
rect 5128 7104 5448 8128
rect 5128 7040 5136 7104
rect 5200 7040 5216 7104
rect 5280 7040 5296 7104
rect 5360 7040 5376 7104
rect 5440 7040 5448 7104
rect 5128 6016 5448 7040
rect 5128 5952 5136 6016
rect 5200 5952 5216 6016
rect 5280 5952 5296 6016
rect 5360 5952 5376 6016
rect 5440 5952 5448 6016
rect 5128 4928 5448 5952
rect 5128 4864 5136 4928
rect 5200 4864 5216 4928
rect 5280 4864 5296 4928
rect 5360 4864 5376 4928
rect 5440 4864 5448 4928
rect 5128 3840 5448 4864
rect 5128 3776 5136 3840
rect 5200 3776 5216 3840
rect 5280 3776 5296 3840
rect 5360 3776 5376 3840
rect 5440 3776 5448 3840
rect 5128 2752 5448 3776
rect 5128 2688 5136 2752
rect 5200 2688 5216 2752
rect 5280 2688 5296 2752
rect 5360 2688 5376 2752
rect 5440 2688 5448 2752
rect 5128 2128 5448 2688
rect 5788 37024 6108 37584
rect 5788 36960 5796 37024
rect 5860 36960 5876 37024
rect 5940 36960 5956 37024
rect 6020 36960 6036 37024
rect 6100 36960 6108 37024
rect 5788 35936 6108 36960
rect 35848 37568 36168 37584
rect 35848 37504 35856 37568
rect 35920 37504 35936 37568
rect 36000 37504 36016 37568
rect 36080 37504 36096 37568
rect 36160 37504 36168 37568
rect 14595 36548 14661 36549
rect 14595 36484 14596 36548
rect 14660 36484 14661 36548
rect 14595 36483 14661 36484
rect 5788 35872 5796 35936
rect 5860 35872 5876 35936
rect 5940 35872 5956 35936
rect 6020 35872 6036 35936
rect 6100 35872 6108 35936
rect 5788 34848 6108 35872
rect 5788 34784 5796 34848
rect 5860 34784 5876 34848
rect 5940 34784 5956 34848
rect 6020 34784 6036 34848
rect 6100 34784 6108 34848
rect 5788 33760 6108 34784
rect 5788 33696 5796 33760
rect 5860 33696 5876 33760
rect 5940 33696 5956 33760
rect 6020 33696 6036 33760
rect 6100 33696 6108 33760
rect 5788 32672 6108 33696
rect 5788 32608 5796 32672
rect 5860 32608 5876 32672
rect 5940 32608 5956 32672
rect 6020 32608 6036 32672
rect 6100 32608 6108 32672
rect 5788 31584 6108 32608
rect 5788 31520 5796 31584
rect 5860 31520 5876 31584
rect 5940 31520 5956 31584
rect 6020 31520 6036 31584
rect 6100 31520 6108 31584
rect 5788 30496 6108 31520
rect 5788 30432 5796 30496
rect 5860 30432 5876 30496
rect 5940 30432 5956 30496
rect 6020 30432 6036 30496
rect 6100 30432 6108 30496
rect 5788 29408 6108 30432
rect 5788 29344 5796 29408
rect 5860 29344 5876 29408
rect 5940 29344 5956 29408
rect 6020 29344 6036 29408
rect 6100 29344 6108 29408
rect 5788 28320 6108 29344
rect 5788 28256 5796 28320
rect 5860 28256 5876 28320
rect 5940 28256 5956 28320
rect 6020 28256 6036 28320
rect 6100 28256 6108 28320
rect 5788 27232 6108 28256
rect 5788 27168 5796 27232
rect 5860 27168 5876 27232
rect 5940 27168 5956 27232
rect 6020 27168 6036 27232
rect 6100 27168 6108 27232
rect 5788 26144 6108 27168
rect 5788 26080 5796 26144
rect 5860 26080 5876 26144
rect 5940 26080 5956 26144
rect 6020 26080 6036 26144
rect 6100 26080 6108 26144
rect 5788 25056 6108 26080
rect 5788 24992 5796 25056
rect 5860 24992 5876 25056
rect 5940 24992 5956 25056
rect 6020 24992 6036 25056
rect 6100 24992 6108 25056
rect 5788 23968 6108 24992
rect 5788 23904 5796 23968
rect 5860 23904 5876 23968
rect 5940 23904 5956 23968
rect 6020 23904 6036 23968
rect 6100 23904 6108 23968
rect 5788 22880 6108 23904
rect 5788 22816 5796 22880
rect 5860 22816 5876 22880
rect 5940 22816 5956 22880
rect 6020 22816 6036 22880
rect 6100 22816 6108 22880
rect 5788 21792 6108 22816
rect 5788 21728 5796 21792
rect 5860 21728 5876 21792
rect 5940 21728 5956 21792
rect 6020 21728 6036 21792
rect 6100 21728 6108 21792
rect 5788 20704 6108 21728
rect 5788 20640 5796 20704
rect 5860 20640 5876 20704
rect 5940 20640 5956 20704
rect 6020 20640 6036 20704
rect 6100 20640 6108 20704
rect 5788 19616 6108 20640
rect 5788 19552 5796 19616
rect 5860 19552 5876 19616
rect 5940 19552 5956 19616
rect 6020 19552 6036 19616
rect 6100 19552 6108 19616
rect 5788 18528 6108 19552
rect 5788 18464 5796 18528
rect 5860 18464 5876 18528
rect 5940 18464 5956 18528
rect 6020 18464 6036 18528
rect 6100 18464 6108 18528
rect 5788 17440 6108 18464
rect 5788 17376 5796 17440
rect 5860 17376 5876 17440
rect 5940 17376 5956 17440
rect 6020 17376 6036 17440
rect 6100 17376 6108 17440
rect 5788 16352 6108 17376
rect 5788 16288 5796 16352
rect 5860 16288 5876 16352
rect 5940 16288 5956 16352
rect 6020 16288 6036 16352
rect 6100 16288 6108 16352
rect 5788 15264 6108 16288
rect 5788 15200 5796 15264
rect 5860 15200 5876 15264
rect 5940 15200 5956 15264
rect 6020 15200 6036 15264
rect 6100 15200 6108 15264
rect 5788 14176 6108 15200
rect 5788 14112 5796 14176
rect 5860 14112 5876 14176
rect 5940 14112 5956 14176
rect 6020 14112 6036 14176
rect 6100 14112 6108 14176
rect 5788 13088 6108 14112
rect 5788 13024 5796 13088
rect 5860 13024 5876 13088
rect 5940 13024 5956 13088
rect 6020 13024 6036 13088
rect 6100 13024 6108 13088
rect 5788 12000 6108 13024
rect 5788 11936 5796 12000
rect 5860 11936 5876 12000
rect 5940 11936 5956 12000
rect 6020 11936 6036 12000
rect 6100 11936 6108 12000
rect 5788 10912 6108 11936
rect 11467 11388 11533 11389
rect 11467 11324 11468 11388
rect 11532 11324 11533 11388
rect 11467 11323 11533 11324
rect 5788 10848 5796 10912
rect 5860 10848 5876 10912
rect 5940 10848 5956 10912
rect 6020 10848 6036 10912
rect 6100 10848 6108 10912
rect 5788 9824 6108 10848
rect 8155 10436 8221 10437
rect 8155 10372 8156 10436
rect 8220 10372 8221 10436
rect 8155 10371 8221 10372
rect 5788 9760 5796 9824
rect 5860 9760 5876 9824
rect 5940 9760 5956 9824
rect 6020 9760 6036 9824
rect 6100 9760 6108 9824
rect 5788 8736 6108 9760
rect 5788 8672 5796 8736
rect 5860 8672 5876 8736
rect 5940 8672 5956 8736
rect 6020 8672 6036 8736
rect 6100 8672 6108 8736
rect 5788 7648 6108 8672
rect 5788 7584 5796 7648
rect 5860 7584 5876 7648
rect 5940 7584 5956 7648
rect 6020 7584 6036 7648
rect 6100 7584 6108 7648
rect 5788 6560 6108 7584
rect 5788 6496 5796 6560
rect 5860 6496 5876 6560
rect 5940 6496 5956 6560
rect 6020 6496 6036 6560
rect 6100 6496 6108 6560
rect 5788 5472 6108 6496
rect 5788 5408 5796 5472
rect 5860 5408 5876 5472
rect 5940 5408 5956 5472
rect 6020 5408 6036 5472
rect 6100 5408 6108 5472
rect 5788 4384 6108 5408
rect 5788 4320 5796 4384
rect 5860 4320 5876 4384
rect 5940 4320 5956 4384
rect 6020 4320 6036 4384
rect 6100 4320 6108 4384
rect 5788 3296 6108 4320
rect 5788 3232 5796 3296
rect 5860 3232 5876 3296
rect 5940 3232 5956 3296
rect 6020 3232 6036 3296
rect 6100 3232 6108 3296
rect 5788 2208 6108 3232
rect 8158 3229 8218 10371
rect 10179 10028 10245 10029
rect 10179 9964 10180 10028
rect 10244 9964 10245 10028
rect 10179 9963 10245 9964
rect 9995 8396 10061 8397
rect 9995 8332 9996 8396
rect 10060 8332 10061 8396
rect 9995 8331 10061 8332
rect 8155 3228 8221 3229
rect 8155 3164 8156 3228
rect 8220 3164 8221 3228
rect 8155 3163 8221 3164
rect 9998 3093 10058 8331
rect 10182 4045 10242 9963
rect 10731 9892 10797 9893
rect 10731 9828 10732 9892
rect 10796 9828 10797 9892
rect 10731 9827 10797 9828
rect 10734 4725 10794 9827
rect 11470 4725 11530 11323
rect 11651 11252 11717 11253
rect 11651 11188 11652 11252
rect 11716 11188 11717 11252
rect 11651 11187 11717 11188
rect 10731 4724 10797 4725
rect 10731 4660 10732 4724
rect 10796 4660 10797 4724
rect 10731 4659 10797 4660
rect 11467 4724 11533 4725
rect 11467 4660 11468 4724
rect 11532 4660 11533 4724
rect 11467 4659 11533 4660
rect 10179 4044 10245 4045
rect 10179 3980 10180 4044
rect 10244 3980 10245 4044
rect 10179 3979 10245 3980
rect 11654 3773 11714 11187
rect 12203 11116 12269 11117
rect 12203 11052 12204 11116
rect 12268 11052 12269 11116
rect 12203 11051 12269 11052
rect 12206 4725 12266 11051
rect 13675 9484 13741 9485
rect 13675 9420 13676 9484
rect 13740 9420 13741 9484
rect 13675 9419 13741 9420
rect 13678 4725 13738 9419
rect 12203 4724 12269 4725
rect 12203 4660 12204 4724
rect 12268 4660 12269 4724
rect 12203 4659 12269 4660
rect 13675 4724 13741 4725
rect 13675 4660 13676 4724
rect 13740 4660 13741 4724
rect 13675 4659 13741 4660
rect 11651 3772 11717 3773
rect 11651 3708 11652 3772
rect 11716 3708 11717 3772
rect 11651 3707 11717 3708
rect 14230 3637 14290 11102
rect 14598 6357 14658 36483
rect 35848 36480 36168 37504
rect 35848 36416 35856 36480
rect 35920 36416 35936 36480
rect 36000 36416 36016 36480
rect 36080 36416 36096 36480
rect 36160 36416 36168 36480
rect 31523 36412 31589 36413
rect 31523 36348 31524 36412
rect 31588 36348 31589 36412
rect 31523 36347 31589 36348
rect 26739 29612 26805 29613
rect 26739 29548 26740 29612
rect 26804 29548 26805 29612
rect 26739 29547 26805 29548
rect 26742 12450 26802 29547
rect 26742 12390 27170 12450
rect 20667 11932 20733 11933
rect 20667 11868 20668 11932
rect 20732 11868 20733 11932
rect 20667 11867 20733 11868
rect 17539 11660 17605 11661
rect 17539 11596 17540 11660
rect 17604 11596 17605 11660
rect 17539 11595 17605 11596
rect 15699 11524 15765 11525
rect 15699 11460 15700 11524
rect 15764 11460 15765 11524
rect 15699 11459 15765 11460
rect 14963 7852 15029 7853
rect 14963 7788 14964 7852
rect 15028 7788 15029 7852
rect 14963 7787 15029 7788
rect 14595 6356 14661 6357
rect 14595 6292 14596 6356
rect 14660 6292 14661 6356
rect 14595 6291 14661 6292
rect 14779 5132 14845 5133
rect 14779 5068 14780 5132
rect 14844 5068 14845 5132
rect 14779 5067 14845 5068
rect 14227 3636 14293 3637
rect 14227 3572 14228 3636
rect 14292 3572 14293 3636
rect 14227 3571 14293 3572
rect 9995 3092 10061 3093
rect 9995 3028 9996 3092
rect 10060 3028 10061 3092
rect 9995 3027 10061 3028
rect 5788 2144 5796 2208
rect 5860 2144 5876 2208
rect 5940 2144 5956 2208
rect 6020 2144 6036 2208
rect 6100 2144 6108 2208
rect 5788 2128 6108 2144
rect 14782 237 14842 5067
rect 14966 3637 15026 7787
rect 15147 7036 15213 7037
rect 15147 6972 15148 7036
rect 15212 6972 15213 7036
rect 15147 6971 15213 6972
rect 14963 3636 15029 3637
rect 14963 3572 14964 3636
rect 15028 3572 15029 3636
rect 14963 3571 15029 3572
rect 15150 2685 15210 6971
rect 15702 5541 15762 11459
rect 15883 10980 15949 10981
rect 15883 10916 15884 10980
rect 15948 10916 15949 10980
rect 15883 10915 15949 10916
rect 15699 5540 15765 5541
rect 15699 5476 15700 5540
rect 15764 5476 15765 5540
rect 15699 5475 15765 5476
rect 15886 3909 15946 10915
rect 17171 9212 17237 9213
rect 17171 9148 17172 9212
rect 17236 9148 17237 9212
rect 17171 9147 17237 9148
rect 16803 9076 16869 9077
rect 16803 9012 16804 9076
rect 16868 9012 16869 9076
rect 16803 9011 16869 9012
rect 16806 4045 16866 9011
rect 16803 4044 16869 4045
rect 16803 3980 16804 4044
rect 16868 3980 16869 4044
rect 16803 3979 16869 3980
rect 15883 3908 15949 3909
rect 15883 3844 15884 3908
rect 15948 3844 15949 3908
rect 15883 3843 15949 3844
rect 17174 3365 17234 9147
rect 17542 4317 17602 11595
rect 19747 9756 19813 9757
rect 19747 9692 19748 9756
rect 19812 9692 19813 9756
rect 19747 9691 19813 9692
rect 20483 9756 20549 9757
rect 20483 9692 20484 9756
rect 20548 9692 20549 9756
rect 20483 9691 20549 9692
rect 19195 9212 19261 9213
rect 19195 9148 19196 9212
rect 19260 9148 19261 9212
rect 19195 9147 19261 9148
rect 18091 8804 18157 8805
rect 18091 8740 18092 8804
rect 18156 8740 18157 8804
rect 18091 8739 18157 8740
rect 17907 7580 17973 7581
rect 17907 7516 17908 7580
rect 17972 7516 17973 7580
rect 17907 7515 17973 7516
rect 17910 5405 17970 7515
rect 17907 5404 17973 5405
rect 17907 5340 17908 5404
rect 17972 5340 17973 5404
rect 17907 5339 17973 5340
rect 17539 4316 17605 4317
rect 17539 4252 17540 4316
rect 17604 4252 17605 4316
rect 17539 4251 17605 4252
rect 17171 3364 17237 3365
rect 17171 3300 17172 3364
rect 17236 3300 17237 3364
rect 17171 3299 17237 3300
rect 15147 2684 15213 2685
rect 15147 2620 15148 2684
rect 15212 2620 15213 2684
rect 15147 2619 15213 2620
rect 18094 2277 18154 8739
rect 18275 8260 18341 8261
rect 18275 8196 18276 8260
rect 18340 8196 18341 8260
rect 18275 8195 18341 8196
rect 18278 3773 18338 8195
rect 19198 5677 19258 9147
rect 19563 8396 19629 8397
rect 19563 8332 19564 8396
rect 19628 8332 19629 8396
rect 19563 8331 19629 8332
rect 19195 5676 19261 5677
rect 19195 5612 19196 5676
rect 19260 5612 19261 5676
rect 19195 5611 19261 5612
rect 18275 3772 18341 3773
rect 18275 3708 18276 3772
rect 18340 3708 18341 3772
rect 18275 3707 18341 3708
rect 18091 2276 18157 2277
rect 18091 2212 18092 2276
rect 18156 2212 18157 2276
rect 18091 2211 18157 2212
rect 18278 1869 18338 3707
rect 19566 2413 19626 8331
rect 19750 2549 19810 9691
rect 20115 8532 20181 8533
rect 20115 8468 20116 8532
rect 20180 8468 20181 8532
rect 20115 8467 20181 8468
rect 20118 7938 20178 8467
rect 20486 3773 20546 9691
rect 20670 4045 20730 11867
rect 23427 11252 23493 11253
rect 23427 11188 23428 11252
rect 23492 11188 23493 11252
rect 23427 11187 23493 11188
rect 21219 10300 21285 10301
rect 21219 10236 21220 10300
rect 21284 10236 21285 10300
rect 21219 10235 21285 10236
rect 20851 10028 20917 10029
rect 20851 9964 20852 10028
rect 20916 9964 20917 10028
rect 20851 9963 20917 9964
rect 20854 5677 20914 9963
rect 21222 6221 21282 10235
rect 21403 9756 21469 9757
rect 21403 9692 21404 9756
rect 21468 9692 21469 9756
rect 21403 9691 21469 9692
rect 21219 6220 21285 6221
rect 21219 6156 21220 6220
rect 21284 6156 21285 6220
rect 21219 6155 21285 6156
rect 20851 5676 20917 5677
rect 20851 5612 20852 5676
rect 20916 5612 20917 5676
rect 20851 5611 20917 5612
rect 21406 4045 21466 9691
rect 23059 8532 23125 8533
rect 23059 8468 23060 8532
rect 23124 8468 23125 8532
rect 23059 8467 23125 8468
rect 22507 8124 22573 8125
rect 22507 8060 22508 8124
rect 22572 8060 22573 8124
rect 22507 8059 22573 8060
rect 22510 7581 22570 8059
rect 22507 7580 22573 7581
rect 22507 7516 22508 7580
rect 22572 7516 22573 7580
rect 22507 7515 22573 7516
rect 22510 6901 22570 7515
rect 22507 6900 22573 6901
rect 22507 6836 22508 6900
rect 22572 6836 22573 6900
rect 22507 6835 22573 6836
rect 20667 4044 20733 4045
rect 20667 3980 20668 4044
rect 20732 3980 20733 4044
rect 20667 3979 20733 3980
rect 21403 4044 21469 4045
rect 21403 3980 21404 4044
rect 21468 3980 21469 4044
rect 21403 3979 21469 3980
rect 20483 3772 20549 3773
rect 20483 3708 20484 3772
rect 20548 3708 20549 3772
rect 20483 3707 20549 3708
rect 22510 2685 22570 6835
rect 23062 5677 23122 8467
rect 23059 5676 23125 5677
rect 23059 5612 23060 5676
rect 23124 5612 23125 5676
rect 23059 5611 23125 5612
rect 23430 5218 23490 11187
rect 24531 11116 24597 11117
rect 24531 11052 24532 11116
rect 24596 11052 24597 11116
rect 24531 11051 24597 11052
rect 24163 9756 24229 9757
rect 24163 9692 24164 9756
rect 24228 9692 24229 9756
rect 24163 9691 24229 9692
rect 24166 5677 24226 9691
rect 24347 9620 24413 9621
rect 24347 9556 24348 9620
rect 24412 9556 24413 9620
rect 24347 9555 24413 9556
rect 24350 8125 24410 9555
rect 24347 8124 24413 8125
rect 24347 8060 24348 8124
rect 24412 8060 24413 8124
rect 24347 8059 24413 8060
rect 24534 6493 24594 11051
rect 25819 10844 25885 10845
rect 25819 10780 25820 10844
rect 25884 10780 25885 10844
rect 25819 10779 25885 10780
rect 24899 8940 24965 8941
rect 24899 8876 24900 8940
rect 24964 8876 24965 8940
rect 24899 8875 24965 8876
rect 24531 6492 24597 6493
rect 24531 6428 24532 6492
rect 24596 6428 24597 6492
rect 24531 6427 24597 6428
rect 24163 5676 24229 5677
rect 24163 5612 24164 5676
rect 24228 5612 24229 5676
rect 24163 5611 24229 5612
rect 23430 4725 23490 4982
rect 23427 4724 23493 4725
rect 23427 4660 23428 4724
rect 23492 4660 23493 4724
rect 23427 4659 23493 4660
rect 24902 4181 24962 8875
rect 25083 7852 25149 7853
rect 25083 7788 25084 7852
rect 25148 7788 25149 7852
rect 25083 7787 25149 7788
rect 25086 5677 25146 7787
rect 25822 7445 25882 10779
rect 26003 10436 26069 10437
rect 26003 10372 26004 10436
rect 26068 10372 26069 10436
rect 26003 10371 26069 10372
rect 25819 7444 25885 7445
rect 25819 7380 25820 7444
rect 25884 7380 25885 7444
rect 25819 7379 25885 7380
rect 26006 7173 26066 10371
rect 26187 9756 26253 9757
rect 26187 9692 26188 9756
rect 26252 9692 26253 9756
rect 26187 9691 26253 9692
rect 26003 7172 26069 7173
rect 26003 7108 26004 7172
rect 26068 7108 26069 7172
rect 26003 7107 26069 7108
rect 25635 6764 25701 6765
rect 25635 6700 25636 6764
rect 25700 6700 25701 6764
rect 25635 6699 25701 6700
rect 25083 5676 25149 5677
rect 25083 5612 25084 5676
rect 25148 5612 25149 5676
rect 25083 5611 25149 5612
rect 24899 4180 24965 4181
rect 24899 4116 24900 4180
rect 24964 4116 24965 4180
rect 24899 4115 24965 4116
rect 22507 2684 22573 2685
rect 22507 2620 22508 2684
rect 22572 2620 22573 2684
rect 22507 2619 22573 2620
rect 19747 2548 19813 2549
rect 19747 2484 19748 2548
rect 19812 2484 19813 2548
rect 19747 2483 19813 2484
rect 19563 2412 19629 2413
rect 19563 2348 19564 2412
rect 19628 2348 19629 2412
rect 19563 2347 19629 2348
rect 24902 2141 24962 4115
rect 25638 3773 25698 6699
rect 26190 3909 26250 9691
rect 27110 9349 27170 12390
rect 30787 10164 30853 10165
rect 30787 10100 30788 10164
rect 30852 10100 30853 10164
rect 30787 10099 30853 10100
rect 28027 10028 28093 10029
rect 28027 9964 28028 10028
rect 28092 9964 28093 10028
rect 28027 9963 28093 9964
rect 27107 9348 27173 9349
rect 27107 9284 27108 9348
rect 27172 9284 27173 9348
rect 27107 9283 27173 9284
rect 26923 5948 26989 5949
rect 26923 5884 26924 5948
rect 26988 5884 26989 5948
rect 26923 5883 26989 5884
rect 26926 4453 26986 5883
rect 26923 4452 26989 4453
rect 26923 4388 26924 4452
rect 26988 4388 26989 4452
rect 26923 4387 26989 4388
rect 26187 3908 26253 3909
rect 26187 3844 26188 3908
rect 26252 3844 26253 3908
rect 26187 3843 26253 3844
rect 25635 3772 25701 3773
rect 25635 3708 25636 3772
rect 25700 3708 25701 3772
rect 25635 3707 25701 3708
rect 26926 3365 26986 4387
rect 26923 3364 26989 3365
rect 26923 3300 26924 3364
rect 26988 3300 26989 3364
rect 26923 3299 26989 3300
rect 27110 2957 27170 9283
rect 27291 9212 27357 9213
rect 27291 9148 27292 9212
rect 27356 9148 27357 9212
rect 27291 9147 27357 9148
rect 27294 6901 27354 9147
rect 27475 8940 27541 8941
rect 27475 8876 27476 8940
rect 27540 8876 27541 8940
rect 27475 8875 27541 8876
rect 27291 6900 27357 6901
rect 27291 6836 27292 6900
rect 27356 6836 27357 6900
rect 27291 6835 27357 6836
rect 27478 5813 27538 8875
rect 27659 8668 27725 8669
rect 27659 8604 27660 8668
rect 27724 8604 27725 8668
rect 27659 8603 27725 8604
rect 27475 5812 27541 5813
rect 27475 5748 27476 5812
rect 27540 5748 27541 5812
rect 27475 5747 27541 5748
rect 27662 5269 27722 8603
rect 27659 5268 27725 5269
rect 27659 5204 27660 5268
rect 27724 5204 27725 5268
rect 27659 5203 27725 5204
rect 28030 4589 28090 9963
rect 29131 9756 29197 9757
rect 29131 9692 29132 9756
rect 29196 9692 29197 9756
rect 29131 9691 29197 9692
rect 28211 8396 28277 8397
rect 28211 8332 28212 8396
rect 28276 8332 28277 8396
rect 28211 8331 28277 8332
rect 28214 7173 28274 8331
rect 28211 7172 28277 7173
rect 28211 7108 28212 7172
rect 28276 7108 28277 7172
rect 28211 7107 28277 7108
rect 29134 5677 29194 9691
rect 29315 9620 29381 9621
rect 29315 9556 29316 9620
rect 29380 9556 29381 9620
rect 29315 9555 29381 9556
rect 29683 9620 29749 9621
rect 29683 9556 29684 9620
rect 29748 9556 29749 9620
rect 29683 9555 29749 9556
rect 29318 6629 29378 9555
rect 29315 6628 29381 6629
rect 29315 6564 29316 6628
rect 29380 6564 29381 6628
rect 29315 6563 29381 6564
rect 29131 5676 29197 5677
rect 29131 5612 29132 5676
rect 29196 5612 29197 5676
rect 29131 5611 29197 5612
rect 28027 4588 28093 4589
rect 28027 4524 28028 4588
rect 28092 4524 28093 4588
rect 28027 4523 28093 4524
rect 28947 4588 29013 4589
rect 28947 4524 28948 4588
rect 29012 4524 29013 4588
rect 28947 4523 29013 4524
rect 27107 2956 27173 2957
rect 27107 2892 27108 2956
rect 27172 2892 27173 2956
rect 27107 2891 27173 2892
rect 24899 2140 24965 2141
rect 24899 2076 24900 2140
rect 24964 2076 24965 2140
rect 24899 2075 24965 2076
rect 18275 1868 18341 1869
rect 18275 1804 18276 1868
rect 18340 1804 18341 1868
rect 18275 1803 18341 1804
rect 14779 236 14845 237
rect 14779 172 14780 236
rect 14844 172 14845 236
rect 14779 171 14845 172
rect 28950 101 29010 4523
rect 29686 2277 29746 9555
rect 30603 8532 30669 8533
rect 30603 8468 30604 8532
rect 30668 8468 30669 8532
rect 30603 8467 30669 8468
rect 30606 5269 30666 8467
rect 30603 5268 30669 5269
rect 30603 5204 30604 5268
rect 30668 5204 30669 5268
rect 30603 5203 30669 5204
rect 29683 2276 29749 2277
rect 29683 2212 29684 2276
rect 29748 2212 29749 2276
rect 29683 2211 29749 2212
rect 30790 1597 30850 10099
rect 31155 9620 31221 9621
rect 31155 9556 31156 9620
rect 31220 9556 31221 9620
rect 31155 9555 31221 9556
rect 30971 9484 31037 9485
rect 30971 9420 30972 9484
rect 31036 9420 31037 9484
rect 30971 9419 31037 9420
rect 30974 4861 31034 9419
rect 31158 6493 31218 9555
rect 31526 7581 31586 36347
rect 35848 35392 36168 36416
rect 35848 35328 35856 35392
rect 35920 35328 35936 35392
rect 36000 35328 36016 35392
rect 36080 35328 36096 35392
rect 36160 35328 36168 35392
rect 35848 34304 36168 35328
rect 35848 34240 35856 34304
rect 35920 34240 35936 34304
rect 36000 34240 36016 34304
rect 36080 34240 36096 34304
rect 36160 34240 36168 34304
rect 35848 33216 36168 34240
rect 35848 33152 35856 33216
rect 35920 33152 35936 33216
rect 36000 33152 36016 33216
rect 36080 33152 36096 33216
rect 36160 33152 36168 33216
rect 33179 32468 33245 32469
rect 33179 32404 33180 32468
rect 33244 32404 33245 32468
rect 33179 32403 33245 32404
rect 32627 9620 32693 9621
rect 32627 9556 32628 9620
rect 32692 9556 32693 9620
rect 32627 9555 32693 9556
rect 32443 9484 32509 9485
rect 32443 9420 32444 9484
rect 32508 9420 32509 9484
rect 32443 9419 32509 9420
rect 31523 7580 31589 7581
rect 31523 7516 31524 7580
rect 31588 7516 31589 7580
rect 31523 7515 31589 7516
rect 31155 6492 31221 6493
rect 31155 6428 31156 6492
rect 31220 6428 31221 6492
rect 31155 6427 31221 6428
rect 31523 5812 31589 5813
rect 31523 5748 31524 5812
rect 31588 5748 31589 5812
rect 31523 5747 31589 5748
rect 30971 4860 31037 4861
rect 30971 4796 30972 4860
rect 31036 4796 31037 4860
rect 30971 4795 31037 4796
rect 30787 1596 30853 1597
rect 30787 1532 30788 1596
rect 30852 1532 30853 1596
rect 30787 1531 30853 1532
rect 31526 1325 31586 5747
rect 32446 5405 32506 9419
rect 32630 6765 32690 9555
rect 32995 8396 33061 8397
rect 32995 8332 32996 8396
rect 33060 8332 33061 8396
rect 32995 8331 33061 8332
rect 32811 7444 32877 7445
rect 32811 7380 32812 7444
rect 32876 7380 32877 7444
rect 32811 7379 32877 7380
rect 32627 6764 32693 6765
rect 32627 6700 32628 6764
rect 32692 6700 32693 6764
rect 32627 6699 32693 6700
rect 32443 5404 32509 5405
rect 32443 5340 32444 5404
rect 32508 5340 32509 5404
rect 32443 5339 32509 5340
rect 32814 3365 32874 7379
rect 32811 3364 32877 3365
rect 32811 3300 32812 3364
rect 32876 3300 32877 3364
rect 32811 3299 32877 3300
rect 32998 2957 33058 8331
rect 33182 8125 33242 32403
rect 35848 32128 36168 33152
rect 35848 32064 35856 32128
rect 35920 32064 35936 32128
rect 36000 32064 36016 32128
rect 36080 32064 36096 32128
rect 36160 32064 36168 32128
rect 35848 31040 36168 32064
rect 35848 30976 35856 31040
rect 35920 30976 35936 31040
rect 36000 30976 36016 31040
rect 36080 30976 36096 31040
rect 36160 30976 36168 31040
rect 35848 29952 36168 30976
rect 35848 29888 35856 29952
rect 35920 29888 35936 29952
rect 36000 29888 36016 29952
rect 36080 29888 36096 29952
rect 36160 29888 36168 29952
rect 35848 28864 36168 29888
rect 35848 28800 35856 28864
rect 35920 28800 35936 28864
rect 36000 28800 36016 28864
rect 36080 28800 36096 28864
rect 36160 28800 36168 28864
rect 35848 27776 36168 28800
rect 35848 27712 35856 27776
rect 35920 27712 35936 27776
rect 36000 27712 36016 27776
rect 36080 27712 36096 27776
rect 36160 27712 36168 27776
rect 35848 26688 36168 27712
rect 35848 26624 35856 26688
rect 35920 26624 35936 26688
rect 36000 26624 36016 26688
rect 36080 26624 36096 26688
rect 36160 26624 36168 26688
rect 35848 25600 36168 26624
rect 35848 25536 35856 25600
rect 35920 25536 35936 25600
rect 36000 25536 36016 25600
rect 36080 25536 36096 25600
rect 36160 25536 36168 25600
rect 35848 24512 36168 25536
rect 35848 24448 35856 24512
rect 35920 24448 35936 24512
rect 36000 24448 36016 24512
rect 36080 24448 36096 24512
rect 36160 24448 36168 24512
rect 35848 23424 36168 24448
rect 35848 23360 35856 23424
rect 35920 23360 35936 23424
rect 36000 23360 36016 23424
rect 36080 23360 36096 23424
rect 36160 23360 36168 23424
rect 35848 22336 36168 23360
rect 35848 22272 35856 22336
rect 35920 22272 35936 22336
rect 36000 22272 36016 22336
rect 36080 22272 36096 22336
rect 36160 22272 36168 22336
rect 35848 21248 36168 22272
rect 35848 21184 35856 21248
rect 35920 21184 35936 21248
rect 36000 21184 36016 21248
rect 36080 21184 36096 21248
rect 36160 21184 36168 21248
rect 35848 20160 36168 21184
rect 35848 20096 35856 20160
rect 35920 20096 35936 20160
rect 36000 20096 36016 20160
rect 36080 20096 36096 20160
rect 36160 20096 36168 20160
rect 35848 19072 36168 20096
rect 35848 19008 35856 19072
rect 35920 19008 35936 19072
rect 36000 19008 36016 19072
rect 36080 19008 36096 19072
rect 36160 19008 36168 19072
rect 35848 17984 36168 19008
rect 35848 17920 35856 17984
rect 35920 17920 35936 17984
rect 36000 17920 36016 17984
rect 36080 17920 36096 17984
rect 36160 17920 36168 17984
rect 35848 16896 36168 17920
rect 35848 16832 35856 16896
rect 35920 16832 35936 16896
rect 36000 16832 36016 16896
rect 36080 16832 36096 16896
rect 36160 16832 36168 16896
rect 35848 15808 36168 16832
rect 35848 15744 35856 15808
rect 35920 15744 35936 15808
rect 36000 15744 36016 15808
rect 36080 15744 36096 15808
rect 36160 15744 36168 15808
rect 35848 14720 36168 15744
rect 35848 14656 35856 14720
rect 35920 14656 35936 14720
rect 36000 14656 36016 14720
rect 36080 14656 36096 14720
rect 36160 14656 36168 14720
rect 35848 13632 36168 14656
rect 35848 13568 35856 13632
rect 35920 13568 35936 13632
rect 36000 13568 36016 13632
rect 36080 13568 36096 13632
rect 36160 13568 36168 13632
rect 35848 12544 36168 13568
rect 35848 12480 35856 12544
rect 35920 12480 35936 12544
rect 36000 12480 36016 12544
rect 36080 12480 36096 12544
rect 36160 12480 36168 12544
rect 35848 11456 36168 12480
rect 35848 11392 35856 11456
rect 35920 11392 35936 11456
rect 36000 11392 36016 11456
rect 36080 11392 36096 11456
rect 36160 11392 36168 11456
rect 35848 10368 36168 11392
rect 35848 10304 35856 10368
rect 35920 10304 35936 10368
rect 36000 10304 36016 10368
rect 36080 10304 36096 10368
rect 36160 10304 36168 10368
rect 34283 9756 34349 9757
rect 34283 9692 34284 9756
rect 34348 9692 34349 9756
rect 34283 9691 34349 9692
rect 33915 9212 33981 9213
rect 33915 9148 33916 9212
rect 33980 9148 33981 9212
rect 33915 9147 33981 9148
rect 33363 8532 33429 8533
rect 33363 8468 33364 8532
rect 33428 8468 33429 8532
rect 33363 8467 33429 8468
rect 33179 8124 33245 8125
rect 33179 8060 33180 8124
rect 33244 8060 33245 8124
rect 33179 8059 33245 8060
rect 33366 3229 33426 8467
rect 33918 7173 33978 9147
rect 33915 7172 33981 7173
rect 33915 7108 33916 7172
rect 33980 7108 33981 7172
rect 33915 7107 33981 7108
rect 33363 3228 33429 3229
rect 33363 3164 33364 3228
rect 33428 3164 33429 3228
rect 33363 3163 33429 3164
rect 32995 2956 33061 2957
rect 32995 2892 32996 2956
rect 33060 2892 33061 2956
rect 32995 2891 33061 2892
rect 34286 2141 34346 9691
rect 35848 9280 36168 10304
rect 35848 9216 35856 9280
rect 35920 9216 35936 9280
rect 36000 9216 36016 9280
rect 36080 9216 36096 9280
rect 36160 9216 36168 9280
rect 35203 8940 35269 8941
rect 35203 8876 35204 8940
rect 35268 8876 35269 8940
rect 35203 8875 35269 8876
rect 34835 8396 34901 8397
rect 34835 8332 34836 8396
rect 34900 8332 34901 8396
rect 34835 8331 34901 8332
rect 34838 5133 34898 8331
rect 34835 5132 34901 5133
rect 34835 5068 34836 5132
rect 34900 5068 34901 5132
rect 34835 5067 34901 5068
rect 35206 3365 35266 8875
rect 35571 8668 35637 8669
rect 35571 8604 35572 8668
rect 35636 8604 35637 8668
rect 35571 8603 35637 8604
rect 35387 7580 35453 7581
rect 35387 7516 35388 7580
rect 35452 7516 35453 7580
rect 35387 7515 35453 7516
rect 35390 5541 35450 7515
rect 35387 5540 35453 5541
rect 35387 5476 35388 5540
rect 35452 5476 35453 5540
rect 35387 5475 35453 5476
rect 35574 5133 35634 8603
rect 35848 8192 36168 9216
rect 36508 37024 36828 37584
rect 36508 36960 36516 37024
rect 36580 36960 36596 37024
rect 36660 36960 36676 37024
rect 36740 36960 36756 37024
rect 36820 36960 36828 37024
rect 36508 35936 36828 36960
rect 36508 35872 36516 35936
rect 36580 35872 36596 35936
rect 36660 35872 36676 35936
rect 36740 35872 36756 35936
rect 36820 35872 36828 35936
rect 36508 34848 36828 35872
rect 36508 34784 36516 34848
rect 36580 34784 36596 34848
rect 36660 34784 36676 34848
rect 36740 34784 36756 34848
rect 36820 34784 36828 34848
rect 36508 33760 36828 34784
rect 36508 33696 36516 33760
rect 36580 33696 36596 33760
rect 36660 33696 36676 33760
rect 36740 33696 36756 33760
rect 36820 33696 36828 33760
rect 36508 32672 36828 33696
rect 36508 32608 36516 32672
rect 36580 32608 36596 32672
rect 36660 32608 36676 32672
rect 36740 32608 36756 32672
rect 36820 32608 36828 32672
rect 36508 31584 36828 32608
rect 36508 31520 36516 31584
rect 36580 31520 36596 31584
rect 36660 31520 36676 31584
rect 36740 31520 36756 31584
rect 36820 31520 36828 31584
rect 36508 30496 36828 31520
rect 36508 30432 36516 30496
rect 36580 30432 36596 30496
rect 36660 30432 36676 30496
rect 36740 30432 36756 30496
rect 36820 30432 36828 30496
rect 36508 29408 36828 30432
rect 36508 29344 36516 29408
rect 36580 29344 36596 29408
rect 36660 29344 36676 29408
rect 36740 29344 36756 29408
rect 36820 29344 36828 29408
rect 36508 28320 36828 29344
rect 36508 28256 36516 28320
rect 36580 28256 36596 28320
rect 36660 28256 36676 28320
rect 36740 28256 36756 28320
rect 36820 28256 36828 28320
rect 36508 27232 36828 28256
rect 36508 27168 36516 27232
rect 36580 27168 36596 27232
rect 36660 27168 36676 27232
rect 36740 27168 36756 27232
rect 36820 27168 36828 27232
rect 36508 26144 36828 27168
rect 36508 26080 36516 26144
rect 36580 26080 36596 26144
rect 36660 26080 36676 26144
rect 36740 26080 36756 26144
rect 36820 26080 36828 26144
rect 36508 25056 36828 26080
rect 36508 24992 36516 25056
rect 36580 24992 36596 25056
rect 36660 24992 36676 25056
rect 36740 24992 36756 25056
rect 36820 24992 36828 25056
rect 36508 23968 36828 24992
rect 36508 23904 36516 23968
rect 36580 23904 36596 23968
rect 36660 23904 36676 23968
rect 36740 23904 36756 23968
rect 36820 23904 36828 23968
rect 36508 22880 36828 23904
rect 36508 22816 36516 22880
rect 36580 22816 36596 22880
rect 36660 22816 36676 22880
rect 36740 22816 36756 22880
rect 36820 22816 36828 22880
rect 36508 21792 36828 22816
rect 36508 21728 36516 21792
rect 36580 21728 36596 21792
rect 36660 21728 36676 21792
rect 36740 21728 36756 21792
rect 36820 21728 36828 21792
rect 36508 20704 36828 21728
rect 36508 20640 36516 20704
rect 36580 20640 36596 20704
rect 36660 20640 36676 20704
rect 36740 20640 36756 20704
rect 36820 20640 36828 20704
rect 36508 19616 36828 20640
rect 36508 19552 36516 19616
rect 36580 19552 36596 19616
rect 36660 19552 36676 19616
rect 36740 19552 36756 19616
rect 36820 19552 36828 19616
rect 36508 18528 36828 19552
rect 36508 18464 36516 18528
rect 36580 18464 36596 18528
rect 36660 18464 36676 18528
rect 36740 18464 36756 18528
rect 36820 18464 36828 18528
rect 36508 17440 36828 18464
rect 36508 17376 36516 17440
rect 36580 17376 36596 17440
rect 36660 17376 36676 17440
rect 36740 17376 36756 17440
rect 36820 17376 36828 17440
rect 36508 16352 36828 17376
rect 36508 16288 36516 16352
rect 36580 16288 36596 16352
rect 36660 16288 36676 16352
rect 36740 16288 36756 16352
rect 36820 16288 36828 16352
rect 36508 15264 36828 16288
rect 36508 15200 36516 15264
rect 36580 15200 36596 15264
rect 36660 15200 36676 15264
rect 36740 15200 36756 15264
rect 36820 15200 36828 15264
rect 36508 14176 36828 15200
rect 36508 14112 36516 14176
rect 36580 14112 36596 14176
rect 36660 14112 36676 14176
rect 36740 14112 36756 14176
rect 36820 14112 36828 14176
rect 36508 13088 36828 14112
rect 36508 13024 36516 13088
rect 36580 13024 36596 13088
rect 36660 13024 36676 13088
rect 36740 13024 36756 13088
rect 36820 13024 36828 13088
rect 36508 12000 36828 13024
rect 36508 11936 36516 12000
rect 36580 11936 36596 12000
rect 36660 11936 36676 12000
rect 36740 11936 36756 12000
rect 36820 11936 36828 12000
rect 36508 10912 36828 11936
rect 36508 10848 36516 10912
rect 36580 10848 36596 10912
rect 36660 10848 36676 10912
rect 36740 10848 36756 10912
rect 36820 10848 36828 10912
rect 36508 9824 36828 10848
rect 66568 37568 66888 37584
rect 66568 37504 66576 37568
rect 66640 37504 66656 37568
rect 66720 37504 66736 37568
rect 66800 37504 66816 37568
rect 66880 37504 66888 37568
rect 66568 36480 66888 37504
rect 66568 36416 66576 36480
rect 66640 36416 66656 36480
rect 66720 36416 66736 36480
rect 66800 36416 66816 36480
rect 66880 36416 66888 36480
rect 66568 35392 66888 36416
rect 66568 35328 66576 35392
rect 66640 35328 66656 35392
rect 66720 35328 66736 35392
rect 66800 35328 66816 35392
rect 66880 35328 66888 35392
rect 66568 34304 66888 35328
rect 66568 34240 66576 34304
rect 66640 34240 66656 34304
rect 66720 34240 66736 34304
rect 66800 34240 66816 34304
rect 66880 34240 66888 34304
rect 66568 33216 66888 34240
rect 66568 33152 66576 33216
rect 66640 33152 66656 33216
rect 66720 33152 66736 33216
rect 66800 33152 66816 33216
rect 66880 33152 66888 33216
rect 66568 32128 66888 33152
rect 66568 32064 66576 32128
rect 66640 32064 66656 32128
rect 66720 32064 66736 32128
rect 66800 32064 66816 32128
rect 66880 32064 66888 32128
rect 66568 31040 66888 32064
rect 66568 30976 66576 31040
rect 66640 30976 66656 31040
rect 66720 30976 66736 31040
rect 66800 30976 66816 31040
rect 66880 30976 66888 31040
rect 66568 29952 66888 30976
rect 66568 29888 66576 29952
rect 66640 29888 66656 29952
rect 66720 29888 66736 29952
rect 66800 29888 66816 29952
rect 66880 29888 66888 29952
rect 66568 28864 66888 29888
rect 66568 28800 66576 28864
rect 66640 28800 66656 28864
rect 66720 28800 66736 28864
rect 66800 28800 66816 28864
rect 66880 28800 66888 28864
rect 66568 27776 66888 28800
rect 66568 27712 66576 27776
rect 66640 27712 66656 27776
rect 66720 27712 66736 27776
rect 66800 27712 66816 27776
rect 66880 27712 66888 27776
rect 66568 26688 66888 27712
rect 66568 26624 66576 26688
rect 66640 26624 66656 26688
rect 66720 26624 66736 26688
rect 66800 26624 66816 26688
rect 66880 26624 66888 26688
rect 66568 25600 66888 26624
rect 66568 25536 66576 25600
rect 66640 25536 66656 25600
rect 66720 25536 66736 25600
rect 66800 25536 66816 25600
rect 66880 25536 66888 25600
rect 66568 24512 66888 25536
rect 66568 24448 66576 24512
rect 66640 24448 66656 24512
rect 66720 24448 66736 24512
rect 66800 24448 66816 24512
rect 66880 24448 66888 24512
rect 66568 23424 66888 24448
rect 66568 23360 66576 23424
rect 66640 23360 66656 23424
rect 66720 23360 66736 23424
rect 66800 23360 66816 23424
rect 66880 23360 66888 23424
rect 66568 22336 66888 23360
rect 66568 22272 66576 22336
rect 66640 22272 66656 22336
rect 66720 22272 66736 22336
rect 66800 22272 66816 22336
rect 66880 22272 66888 22336
rect 66568 21248 66888 22272
rect 66568 21184 66576 21248
rect 66640 21184 66656 21248
rect 66720 21184 66736 21248
rect 66800 21184 66816 21248
rect 66880 21184 66888 21248
rect 66568 20160 66888 21184
rect 66568 20096 66576 20160
rect 66640 20096 66656 20160
rect 66720 20096 66736 20160
rect 66800 20096 66816 20160
rect 66880 20096 66888 20160
rect 66568 19072 66888 20096
rect 66568 19008 66576 19072
rect 66640 19008 66656 19072
rect 66720 19008 66736 19072
rect 66800 19008 66816 19072
rect 66880 19008 66888 19072
rect 66568 17984 66888 19008
rect 66568 17920 66576 17984
rect 66640 17920 66656 17984
rect 66720 17920 66736 17984
rect 66800 17920 66816 17984
rect 66880 17920 66888 17984
rect 66568 16896 66888 17920
rect 66568 16832 66576 16896
rect 66640 16832 66656 16896
rect 66720 16832 66736 16896
rect 66800 16832 66816 16896
rect 66880 16832 66888 16896
rect 66568 15808 66888 16832
rect 66568 15744 66576 15808
rect 66640 15744 66656 15808
rect 66720 15744 66736 15808
rect 66800 15744 66816 15808
rect 66880 15744 66888 15808
rect 66568 14720 66888 15744
rect 66568 14656 66576 14720
rect 66640 14656 66656 14720
rect 66720 14656 66736 14720
rect 66800 14656 66816 14720
rect 66880 14656 66888 14720
rect 66568 13632 66888 14656
rect 66568 13568 66576 13632
rect 66640 13568 66656 13632
rect 66720 13568 66736 13632
rect 66800 13568 66816 13632
rect 66880 13568 66888 13632
rect 66568 12544 66888 13568
rect 66568 12480 66576 12544
rect 66640 12480 66656 12544
rect 66720 12480 66736 12544
rect 66800 12480 66816 12544
rect 66880 12480 66888 12544
rect 66568 11456 66888 12480
rect 66568 11392 66576 11456
rect 66640 11392 66656 11456
rect 66720 11392 66736 11456
rect 66800 11392 66816 11456
rect 66880 11392 66888 11456
rect 37411 10572 37477 10573
rect 37411 10508 37412 10572
rect 37476 10508 37477 10572
rect 37411 10507 37477 10508
rect 37227 10164 37293 10165
rect 37227 10100 37228 10164
rect 37292 10100 37293 10164
rect 37227 10099 37293 10100
rect 36508 9760 36516 9824
rect 36580 9760 36596 9824
rect 36660 9760 36676 9824
rect 36740 9760 36756 9824
rect 36820 9760 36828 9824
rect 36307 9076 36373 9077
rect 36307 9012 36308 9076
rect 36372 9012 36373 9076
rect 36307 9011 36373 9012
rect 35848 8128 35856 8192
rect 35920 8128 35936 8192
rect 36000 8128 36016 8192
rect 36080 8128 36096 8192
rect 36160 8128 36168 8192
rect 35848 7104 36168 8128
rect 35848 7040 35856 7104
rect 35920 7040 35936 7104
rect 36000 7040 36016 7104
rect 36080 7040 36096 7104
rect 36160 7040 36168 7104
rect 35848 6016 36168 7040
rect 35848 5952 35856 6016
rect 35920 5952 35936 6016
rect 36000 5952 36016 6016
rect 36080 5952 36096 6016
rect 36160 5952 36168 6016
rect 35571 5132 35637 5133
rect 35571 5068 35572 5132
rect 35636 5068 35637 5132
rect 35571 5067 35637 5068
rect 35574 4453 35634 5067
rect 35848 4928 36168 5952
rect 35848 4864 35856 4928
rect 35920 4864 35936 4928
rect 36000 4864 36016 4928
rect 36080 4864 36096 4928
rect 36160 4864 36168 4928
rect 35571 4452 35637 4453
rect 35571 4388 35572 4452
rect 35636 4388 35637 4452
rect 35571 4387 35637 4388
rect 35848 3840 36168 4864
rect 35848 3776 35856 3840
rect 35920 3776 35936 3840
rect 36000 3776 36016 3840
rect 36080 3776 36096 3840
rect 36160 3776 36168 3840
rect 35203 3364 35269 3365
rect 35203 3300 35204 3364
rect 35268 3300 35269 3364
rect 35203 3299 35269 3300
rect 35848 2752 36168 3776
rect 35848 2688 35856 2752
rect 35920 2688 35936 2752
rect 36000 2688 36016 2752
rect 36080 2688 36096 2752
rect 36160 2688 36168 2752
rect 34283 2140 34349 2141
rect 34283 2076 34284 2140
rect 34348 2076 34349 2140
rect 35848 2128 36168 2688
rect 36310 2413 36370 9011
rect 36508 8736 36828 9760
rect 36508 8672 36516 8736
rect 36580 8672 36596 8736
rect 36660 8672 36676 8736
rect 36740 8672 36756 8736
rect 36820 8672 36828 8736
rect 36508 7648 36828 8672
rect 36508 7584 36516 7648
rect 36580 7584 36596 7648
rect 36660 7584 36676 7648
rect 36740 7584 36756 7648
rect 36820 7584 36828 7648
rect 36508 6560 36828 7584
rect 36508 6496 36516 6560
rect 36580 6496 36596 6560
rect 36660 6496 36676 6560
rect 36740 6496 36756 6560
rect 36820 6496 36828 6560
rect 36508 5472 36828 6496
rect 36508 5408 36516 5472
rect 36580 5408 36596 5472
rect 36660 5408 36676 5472
rect 36740 5408 36756 5472
rect 36820 5408 36828 5472
rect 36508 4384 36828 5408
rect 36508 4320 36516 4384
rect 36580 4320 36596 4384
rect 36660 4320 36676 4384
rect 36740 4320 36756 4384
rect 36820 4320 36828 4384
rect 36508 3296 36828 4320
rect 36508 3232 36516 3296
rect 36580 3232 36596 3296
rect 36660 3232 36676 3296
rect 36740 3232 36756 3296
rect 36820 3232 36828 3296
rect 36307 2412 36373 2413
rect 36307 2348 36308 2412
rect 36372 2348 36373 2412
rect 36307 2347 36373 2348
rect 36508 2208 36828 3232
rect 37230 2549 37290 10099
rect 37414 3093 37474 10507
rect 66568 10368 66888 11392
rect 66568 10304 66576 10368
rect 66640 10304 66656 10368
rect 66720 10304 66736 10368
rect 66800 10304 66816 10368
rect 66880 10304 66888 10368
rect 66568 9280 66888 10304
rect 66568 9216 66576 9280
rect 66640 9216 66656 9280
rect 66720 9216 66736 9280
rect 66800 9216 66816 9280
rect 66880 9216 66888 9280
rect 66568 8192 66888 9216
rect 66568 8128 66576 8192
rect 66640 8128 66656 8192
rect 66720 8128 66736 8192
rect 66800 8128 66816 8192
rect 66880 8128 66888 8192
rect 66568 7104 66888 8128
rect 66568 7040 66576 7104
rect 66640 7040 66656 7104
rect 66720 7040 66736 7104
rect 66800 7040 66816 7104
rect 66880 7040 66888 7104
rect 66568 6016 66888 7040
rect 66568 5952 66576 6016
rect 66640 5952 66656 6016
rect 66720 5952 66736 6016
rect 66800 5952 66816 6016
rect 66880 5952 66888 6016
rect 66568 4928 66888 5952
rect 66568 4864 66576 4928
rect 66640 4864 66656 4928
rect 66720 4864 66736 4928
rect 66800 4864 66816 4928
rect 66880 4864 66888 4928
rect 66568 3840 66888 4864
rect 66568 3776 66576 3840
rect 66640 3776 66656 3840
rect 66720 3776 66736 3840
rect 66800 3776 66816 3840
rect 66880 3776 66888 3840
rect 37411 3092 37477 3093
rect 37411 3028 37412 3092
rect 37476 3028 37477 3092
rect 37411 3027 37477 3028
rect 66568 2752 66888 3776
rect 66568 2688 66576 2752
rect 66640 2688 66656 2752
rect 66720 2688 66736 2752
rect 66800 2688 66816 2752
rect 66880 2688 66888 2752
rect 37227 2548 37293 2549
rect 37227 2484 37228 2548
rect 37292 2484 37293 2548
rect 37227 2483 37293 2484
rect 36508 2144 36516 2208
rect 36580 2144 36596 2208
rect 36660 2144 36676 2208
rect 36740 2144 36756 2208
rect 36820 2144 36828 2208
rect 36508 2128 36828 2144
rect 66568 2128 66888 2688
rect 67228 37024 67548 37584
rect 67228 36960 67236 37024
rect 67300 36960 67316 37024
rect 67380 36960 67396 37024
rect 67460 36960 67476 37024
rect 67540 36960 67548 37024
rect 67228 35936 67548 36960
rect 67228 35872 67236 35936
rect 67300 35872 67316 35936
rect 67380 35872 67396 35936
rect 67460 35872 67476 35936
rect 67540 35872 67548 35936
rect 67228 34848 67548 35872
rect 67228 34784 67236 34848
rect 67300 34784 67316 34848
rect 67380 34784 67396 34848
rect 67460 34784 67476 34848
rect 67540 34784 67548 34848
rect 67228 33760 67548 34784
rect 67228 33696 67236 33760
rect 67300 33696 67316 33760
rect 67380 33696 67396 33760
rect 67460 33696 67476 33760
rect 67540 33696 67548 33760
rect 67228 32672 67548 33696
rect 67228 32608 67236 32672
rect 67300 32608 67316 32672
rect 67380 32608 67396 32672
rect 67460 32608 67476 32672
rect 67540 32608 67548 32672
rect 67228 31584 67548 32608
rect 67228 31520 67236 31584
rect 67300 31520 67316 31584
rect 67380 31520 67396 31584
rect 67460 31520 67476 31584
rect 67540 31520 67548 31584
rect 67228 30496 67548 31520
rect 67228 30432 67236 30496
rect 67300 30432 67316 30496
rect 67380 30432 67396 30496
rect 67460 30432 67476 30496
rect 67540 30432 67548 30496
rect 67228 29408 67548 30432
rect 67228 29344 67236 29408
rect 67300 29344 67316 29408
rect 67380 29344 67396 29408
rect 67460 29344 67476 29408
rect 67540 29344 67548 29408
rect 67228 28320 67548 29344
rect 67228 28256 67236 28320
rect 67300 28256 67316 28320
rect 67380 28256 67396 28320
rect 67460 28256 67476 28320
rect 67540 28256 67548 28320
rect 67228 27232 67548 28256
rect 67228 27168 67236 27232
rect 67300 27168 67316 27232
rect 67380 27168 67396 27232
rect 67460 27168 67476 27232
rect 67540 27168 67548 27232
rect 67228 26144 67548 27168
rect 67228 26080 67236 26144
rect 67300 26080 67316 26144
rect 67380 26080 67396 26144
rect 67460 26080 67476 26144
rect 67540 26080 67548 26144
rect 67228 25056 67548 26080
rect 67228 24992 67236 25056
rect 67300 24992 67316 25056
rect 67380 24992 67396 25056
rect 67460 24992 67476 25056
rect 67540 24992 67548 25056
rect 67228 23968 67548 24992
rect 67228 23904 67236 23968
rect 67300 23904 67316 23968
rect 67380 23904 67396 23968
rect 67460 23904 67476 23968
rect 67540 23904 67548 23968
rect 67228 22880 67548 23904
rect 67228 22816 67236 22880
rect 67300 22816 67316 22880
rect 67380 22816 67396 22880
rect 67460 22816 67476 22880
rect 67540 22816 67548 22880
rect 67228 21792 67548 22816
rect 67228 21728 67236 21792
rect 67300 21728 67316 21792
rect 67380 21728 67396 21792
rect 67460 21728 67476 21792
rect 67540 21728 67548 21792
rect 67228 20704 67548 21728
rect 67228 20640 67236 20704
rect 67300 20640 67316 20704
rect 67380 20640 67396 20704
rect 67460 20640 67476 20704
rect 67540 20640 67548 20704
rect 67228 19616 67548 20640
rect 67228 19552 67236 19616
rect 67300 19552 67316 19616
rect 67380 19552 67396 19616
rect 67460 19552 67476 19616
rect 67540 19552 67548 19616
rect 67228 18528 67548 19552
rect 67228 18464 67236 18528
rect 67300 18464 67316 18528
rect 67380 18464 67396 18528
rect 67460 18464 67476 18528
rect 67540 18464 67548 18528
rect 67228 17440 67548 18464
rect 67228 17376 67236 17440
rect 67300 17376 67316 17440
rect 67380 17376 67396 17440
rect 67460 17376 67476 17440
rect 67540 17376 67548 17440
rect 67228 16352 67548 17376
rect 67228 16288 67236 16352
rect 67300 16288 67316 16352
rect 67380 16288 67396 16352
rect 67460 16288 67476 16352
rect 67540 16288 67548 16352
rect 67228 15264 67548 16288
rect 67228 15200 67236 15264
rect 67300 15200 67316 15264
rect 67380 15200 67396 15264
rect 67460 15200 67476 15264
rect 67540 15200 67548 15264
rect 67228 14176 67548 15200
rect 67228 14112 67236 14176
rect 67300 14112 67316 14176
rect 67380 14112 67396 14176
rect 67460 14112 67476 14176
rect 67540 14112 67548 14176
rect 67228 13088 67548 14112
rect 67228 13024 67236 13088
rect 67300 13024 67316 13088
rect 67380 13024 67396 13088
rect 67460 13024 67476 13088
rect 67540 13024 67548 13088
rect 67228 12000 67548 13024
rect 67228 11936 67236 12000
rect 67300 11936 67316 12000
rect 67380 11936 67396 12000
rect 67460 11936 67476 12000
rect 67540 11936 67548 12000
rect 67228 10912 67548 11936
rect 67228 10848 67236 10912
rect 67300 10848 67316 10912
rect 67380 10848 67396 10912
rect 67460 10848 67476 10912
rect 67540 10848 67548 10912
rect 67228 9824 67548 10848
rect 67228 9760 67236 9824
rect 67300 9760 67316 9824
rect 67380 9760 67396 9824
rect 67460 9760 67476 9824
rect 67540 9760 67548 9824
rect 67228 8736 67548 9760
rect 67228 8672 67236 8736
rect 67300 8672 67316 8736
rect 67380 8672 67396 8736
rect 67460 8672 67476 8736
rect 67540 8672 67548 8736
rect 67228 7648 67548 8672
rect 67228 7584 67236 7648
rect 67300 7584 67316 7648
rect 67380 7584 67396 7648
rect 67460 7584 67476 7648
rect 67540 7584 67548 7648
rect 67228 6560 67548 7584
rect 67228 6496 67236 6560
rect 67300 6496 67316 6560
rect 67380 6496 67396 6560
rect 67460 6496 67476 6560
rect 67540 6496 67548 6560
rect 67228 5472 67548 6496
rect 67228 5408 67236 5472
rect 67300 5408 67316 5472
rect 67380 5408 67396 5472
rect 67460 5408 67476 5472
rect 67540 5408 67548 5472
rect 67228 4384 67548 5408
rect 67228 4320 67236 4384
rect 67300 4320 67316 4384
rect 67380 4320 67396 4384
rect 67460 4320 67476 4384
rect 67540 4320 67548 4384
rect 67228 3296 67548 4320
rect 67228 3232 67236 3296
rect 67300 3232 67316 3296
rect 67380 3232 67396 3296
rect 67460 3232 67476 3296
rect 67540 3232 67548 3296
rect 67228 2208 67548 3232
rect 67228 2144 67236 2208
rect 67300 2144 67316 2208
rect 67380 2144 67396 2208
rect 67460 2144 67476 2208
rect 67540 2144 67548 2208
rect 67228 2128 67548 2144
rect 34283 2075 34349 2076
rect 31523 1324 31589 1325
rect 31523 1260 31524 1324
rect 31588 1260 31589 1324
rect 31523 1259 31589 1260
rect 28947 100 29013 101
rect 28947 36 28948 100
rect 29012 36 29013 100
rect 28947 35 29013 36
<< via4 >>
rect 14142 11102 14378 11338
rect 20030 7702 20266 7938
rect 26102 11252 26338 11338
rect 26102 11188 26188 11252
rect 26188 11188 26252 11252
rect 26252 11188 26338 11252
rect 26102 11102 26338 11188
rect 23342 4982 23578 5218
rect 41374 7852 41610 7938
rect 41374 7788 41460 7852
rect 41460 7788 41524 7852
rect 41524 7788 41610 7852
rect 41374 7702 41610 7788
rect 40270 5132 40506 5218
rect 40270 5068 40356 5132
rect 40356 5068 40420 5132
rect 40420 5068 40506 5132
rect 40270 4982 40506 5068
<< metal5 >>
rect 14100 11338 26380 11380
rect 14100 11102 14142 11338
rect 14378 11102 26102 11338
rect 26338 11102 26380 11338
rect 14100 11060 26380 11102
rect 19988 7938 41652 7980
rect 19988 7702 20030 7938
rect 20266 7702 41374 7938
rect 41610 7702 41652 7938
rect 19988 7660 41652 7702
rect 23300 5218 40548 5260
rect 23300 4982 23342 5218
rect 23578 4982 40270 5218
rect 40506 4982 40548 5218
rect 23300 4940 40548 4982
use sky130_fd_sc_hd__inv_2  _099_
timestamp 25201
transform 1 0 21712 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 25201
transform 1 0 32568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 25201
transform -1 0 32936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 25201
transform -1 0 35880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 25201
transform 1 0 11592 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _104_
timestamp 25201
transform -1 0 41308 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _105_
timestamp 25201
transform 1 0 27876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _106_
timestamp 25201
transform -1 0 16744 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _107_
timestamp 25201
transform 1 0 20148 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _108_
timestamp 25201
transform -1 0 24104 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _109_
timestamp 25201
transform -1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _110_
timestamp 25201
transform 1 0 14996 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 25201
transform 1 0 20516 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _112_
timestamp 25201
transform -1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _113_
timestamp 25201
transform 1 0 17572 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _114_
timestamp 25201
transform 1 0 9936 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _115_
timestamp 25201
transform 1 0 7360 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _116_
timestamp 25201
transform -1 0 15640 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _117_
timestamp 25201
transform -1 0 22264 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _118_
timestamp 25201
transform 1 0 26772 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _119_
timestamp 25201
transform 1 0 28428 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _120_
timestamp 25201
transform -1 0 31004 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _121_
timestamp 25201
transform -1 0 32936 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _122_
timestamp 25201
transform -1 0 30912 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _123_
timestamp 25201
transform 1 0 31280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _124_
timestamp 25201
transform -1 0 35696 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _125_
timestamp 25201
transform -1 0 36156 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _126_
timestamp 25201
transform -1 0 43240 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _127_
timestamp 25201
transform -1 0 33304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _128_
timestamp 25201
transform -1 0 34684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _129_
timestamp 25201
transform -1 0 16008 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_2  _130_
timestamp 25201
transform -1 0 14536 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _131_
timestamp 25201
transform -1 0 22632 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _132_
timestamp 25201
transform 1 0 14996 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _133_
timestamp 25201
transform 1 0 20792 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _134_
timestamp 25201
transform -1 0 23184 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _135_
timestamp 25201
transform 1 0 17572 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _136_
timestamp 25201
transform 1 0 26404 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 25201
transform 1 0 38916 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _138_
timestamp 25201
transform 1 0 20240 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _139_
timestamp 25201
transform 1 0 24196 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _140_
timestamp 25201
transform -1 0 18216 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _141_
timestamp 25201
transform 1 0 21344 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _142_
timestamp 25201
transform 1 0 20792 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _143_
timestamp 25201
transform -1 0 24472 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _144_
timestamp 25201
transform -1 0 23644 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _145_
timestamp 25201
transform 1 0 22264 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _146_
timestamp 25201
transform 1 0 24472 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _147_
timestamp 25201
transform -1 0 22724 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _148_
timestamp 25201
transform -1 0 20792 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _149_
timestamp 25201
transform 1 0 20424 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _150_
timestamp 25201
transform 1 0 22724 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _151_
timestamp 25201
transform -1 0 26496 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _152_
timestamp 25201
transform -1 0 25484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _153_
timestamp 25201
transform -1 0 22264 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _154_
timestamp 25201
transform 1 0 24288 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _155_
timestamp 25201
transform 1 0 26772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _156_
timestamp 25201
transform 1 0 25300 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _157_
timestamp 25201
transform -1 0 25208 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _158_
timestamp 25201
transform -1 0 25668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _159_
timestamp 25201
transform 1 0 22172 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _160_
timestamp 25201
transform -1 0 28152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _161_
timestamp 25201
transform 1 0 26864 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _162_
timestamp 25201
transform -1 0 35144 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _163_
timestamp 25201
transform -1 0 27784 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _164_
timestamp 25201
transform 1 0 27140 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _165_
timestamp 25201
transform 1 0 25300 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _166_
timestamp 25201
transform 1 0 30452 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _167_
timestamp 25201
transform 1 0 23000 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _168_
timestamp 25201
transform 1 0 33028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _169_
timestamp 25201
transform 1 0 30452 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _170_
timestamp 25201
transform -1 0 29532 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _171_
timestamp 25201
transform 1 0 31096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _172_
timestamp 25201
transform 1 0 25300 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _173_
timestamp 25201
transform -1 0 32200 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _174_
timestamp 25201
transform 1 0 33764 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _175_
timestamp 25201
transform 1 0 32200 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _176_
timestamp 25201
transform -1 0 30360 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _177_
timestamp 25201
transform 1 0 33028 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _178_
timestamp 25201
transform 1 0 35604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _179_
timestamp 25201
transform 1 0 33028 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _180_
timestamp 25201
transform 1 0 34408 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _181_
timestamp 25201
transform 1 0 33856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _182_
timestamp 25201
transform -1 0 40664 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _183_
timestamp 25201
transform -1 0 38088 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _184_
timestamp 25201
transform -1 0 43240 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 25201
transform 1 0 37076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _186_
timestamp 25201
transform -1 0 35512 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _187_
timestamp 25201
transform 1 0 27140 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _188_
timestamp 25201
transform 1 0 35604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _189_
timestamp 25201
transform -1 0 36616 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _190_
timestamp 25201
transform 1 0 34224 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _191_
timestamp 25201
transform -1 0 34776 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _192_
timestamp 25201
transform -1 0 36064 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _193_
timestamp 25201
transform -1 0 28520 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _194_
timestamp 25201
transform -1 0 35880 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _195_
timestamp 25201
transform 1 0 38180 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _196_
timestamp 25201
transform 1 0 32200 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _197_
timestamp 25201
transform 1 0 34776 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _198_
timestamp 25201
transform 1 0 11224 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _199_
timestamp 25201
transform 1 0 12420 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _200_
timestamp 25201
transform 1 0 13800 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _201_
timestamp 25201
transform 1 0 17572 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _202_
timestamp 25201
transform 1 0 19044 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _203_
timestamp 25201
transform 1 0 20884 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _204_
timestamp 25201
transform 1 0 23368 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp 25201
transform 1 0 25668 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 25201
transform 1 0 27876 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _207_
timestamp 25201
transform 1 0 29900 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 25201
transform 1 0 31372 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 25201
transform 1 0 33028 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 25201
transform 1 0 34684 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _211_
timestamp 25201
transform 1 0 36340 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 25201
transform 1 0 40020 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 25201
transform -1 0 41676 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 25201
transform -1 0 44160 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _215_
timestamp 25201
transform -1 0 43240 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _216_
timestamp 25201
transform 1 0 14904 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _217_
timestamp 25201
transform 1 0 18952 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _218_
timestamp 25201
transform -1 0 22264 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _219_
timestamp 25201
transform 1 0 22080 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _220_
timestamp 25201
transform 1 0 23920 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _221_
timestamp 25201
transform 1 0 24196 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _222_
timestamp 25201
transform 1 0 25024 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _223_
timestamp 25201
transform 1 0 26680 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _224_
timestamp 25201
transform 1 0 29624 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _225_
timestamp 25201
transform 1 0 29716 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _226_
timestamp 25201
transform 1 0 30544 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _227_
timestamp 25201
transform 1 0 32108 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _228_
timestamp 25201
transform 1 0 34868 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _229_
timestamp 25201
transform 1 0 35972 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _230_
timestamp 25201
transform 1 0 37904 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _231_
timestamp 25201
transform 1 0 38180 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _232_
timestamp 25201
transform 1 0 33028 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _233_
timestamp 25201
transform 1 0 37444 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _234_
timestamp 25201
transform 1 0 10488 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _235_
timestamp 25201
transform 1 0 11960 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _236_
timestamp 25201
transform 1 0 13064 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _237_
timestamp 25201
transform 1 0 16376 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _238_
timestamp 25201
transform 1 0 18032 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _239_
timestamp 25201
transform 1 0 19872 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _240_
timestamp 25201
transform -1 0 24840 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _241_
timestamp 25201
transform 1 0 25300 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _242_
timestamp 25201
transform 1 0 26680 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _243_
timestamp 25201
transform -1 0 30360 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _244_
timestamp 25201
transform -1 0 32752 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _245_
timestamp 25201
transform 1 0 32292 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _246_
timestamp 25201
transform -1 0 35972 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _247_
timestamp 25201
transform 1 0 36156 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _248_
timestamp 25201
transform 1 0 38364 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _249_
timestamp 25201
transform -1 0 42044 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _250_
timestamp 25201
transform -1 0 43884 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _251_
timestamp 25201
transform 1 0 43332 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _258_
timestamp 25201
transform 1 0 48116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _259_
timestamp 25201
transform 1 0 51520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _260_
timestamp 25201
transform 1 0 53636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _261_
timestamp 25201
transform 1 0 57132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _262_
timestamp 25201
transform 1 0 60720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _263_
timestamp 25201
transform -1 0 64768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _264_
timestamp 25201
transform 1 0 66976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _265_
timestamp 25201
transform 1 0 69092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _266_
timestamp 25201
transform 1 0 70656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _267_
timestamp 25201
transform 1 0 74244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _268_
timestamp 25201
transform 1 0 58420 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _269_
timestamp 25201
transform 1 0 55384 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _270_
timestamp 25201
transform 1 0 51704 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _271_
timestamp 25201
transform 1 0 48024 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _272_
timestamp 25201
transform 1 0 44344 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _273_
timestamp 25201
transform 1 0 40664 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _274_
timestamp 25201
transform -1 0 37260 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _275_
timestamp 25201
transform -1 0 34040 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _276_
timestamp 25201
transform 1 0 29624 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _277_
timestamp 25201
transform 1 0 25944 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _278_
timestamp 25201
transform 1 0 22264 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _279_
timestamp 25201
transform -1 0 19320 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _280_
timestamp 25201
transform 1 0 14904 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _281_
timestamp 25201
transform -1 0 12144 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _282_
timestamp 25201
transform 1 0 7544 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_115
timestamp 25201
transform -1 0 50968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_116
timestamp 25201
transform -1 0 55752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_117
timestamp 25201
transform -1 0 59616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_118
timestamp 25201
transform -1 0 63480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_119
timestamp 25201
transform -1 0 73416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ahb_counter_120
timestamp 25201
transform -1 0 10120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 25201
transform 1 0 27048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 25201
transform -1 0 9016 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 25201
transform 1 0 23092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 25201
transform -1 0 27140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 25201
transform -1 0 29716 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 25201
transform -1 0 17756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 25201
transform -1 0 31096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 25201
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 25201
transform -1 0 26220 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 25201
transform -1 0 28152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 25201
transform 1 0 24472 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 25201
transform -1 0 32016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 25201
transform -1 0 31464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 25201
transform 1 0 36524 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 25201
transform -1 0 26404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 25201
transform -1 0 21896 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 25201
transform 1 0 28980 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 25201
transform -1 0 23920 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 25201
transform 1 0 23276 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 25201
transform 1 0 21712 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 25201
transform -1 0 22908 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 25201
transform -1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 25201
transform 1 0 22080 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 25201
transform 1 0 26496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 25201
transform 1 0 20148 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 25201
transform -1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 25201
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 25201
transform 1 0 30728 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 25201
transform -1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 25201
transform -1 0 33212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 25201
transform -1 0 16928 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 25201
transform 1 0 34868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 25201
transform 1 0 24288 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 25201
transform 1 0 25024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 25201
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 25201
transform -1 0 39100 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 25201
transform 1 0 33304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 25201
transform 1 0 30176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 25201
transform -1 0 20700 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_HCLK
timestamp 25201
transform 1 0 27876 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_HCLK
timestamp 25201
transform -1 0 19872 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_HCLK
timestamp 25201
transform 1 0 22724 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_HCLK
timestamp 25201
transform 1 0 37076 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_HCLK
timestamp 25201
transform 1 0 32568 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp 25201
transform 1 0 18032 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp 25201
transform -1 0 22540 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload2
timestamp 25201
transform -1 0 31096 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout96
timestamp 25201
transform -1 0 23368 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout97
timestamp 25201
transform 1 0 27416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout98
timestamp 25201
transform 1 0 22724 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout99
timestamp 25201
transform -1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout100
timestamp 25201
transform -1 0 38088 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout101
timestamp 25201
transform 1 0 17664 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout104
timestamp 25201
transform -1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout105
timestamp 25201
transform -1 0 33304 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout106
timestamp 25201
transform -1 0 11868 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout107
timestamp 25201
transform 1 0 33396 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout108
timestamp 25201
transform -1 0 10488 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout109
timestamp 25201
transform -1 0 28888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout110
timestamp 25201
transform 1 0 24656 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout111
timestamp 25201
transform 1 0 12512 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout112
timestamp 25201
transform 1 0 9752 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout113
timestamp 25201
transform -1 0 12972 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout114
timestamp 25201
transform 1 0 29900 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3
timestamp 25201
transform 1 0 2300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 25201
transform 1 0 9200 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 25201
transform 1 0 9844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 25201
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 25201
transform 1 0 14996 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 25201
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_273
timestamp 25201
transform 1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_281
timestamp 25201
transform 1 0 27876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_421
timestamp 25201
transform 1 0 40756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_431
timestamp 25201
transform 1 0 41676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_533
timestamp 25201
transform 1 0 51060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_555
timestamp 25201
transform 1 0 53084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 25201
transform 1 0 53452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_577
timestamp 25201
transform 1 0 55108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_584
timestamp 25201
transform 1 0 55752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_589
timestamp 25201
transform 1 0 56212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_597
timestamp 25201
transform 1 0 56948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_633
timestamp 25201
transform 1 0 60260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 25201
transform 1 0 60996 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_661
timestamp 25201
transform 1 0 62836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_668
timestamp 25201
transform 1 0 63480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_673
timestamp 25201
transform 1 0 63940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_681
timestamp 25201
transform 1 0 64676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_701
timestamp 25201
transform 1 0 66516 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_723
timestamp 25201
transform 1 0 68540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_727
timestamp 25201
transform 1 0 68908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_745
timestamp 25201
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_749
timestamp 25201
transform 1 0 70932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_755
timestamp 25201
transform 1 0 71484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_785
timestamp 25201
transform 1 0 74244 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_807
timestamp 25201
transform 1 0 76268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_811
timestamp 25201
transform 1 0 76636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_821
timestamp 25201
transform 1 0 77556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 25201
transform 1 0 2300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_11
timestamp 25201
transform 1 0 3036 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 25201
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 25201
transform 1 0 12420 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_171
timestamp 25201
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 25201
transform 1 0 32752 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_369
timestamp 25201
transform 1 0 35972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 25201
transform 1 0 37996 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 25201
transform 1 0 38180 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_438
timestamp 25201
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_505
timestamp 25201
transform 1 0 48484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_541
timestamp 25201
transform 1 0 51796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_564
timestamp 25201
transform 1 0 53912 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_589
timestamp 25201
transform 1 0 56212 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_597
timestamp 25201
transform 1 0 56948 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_610
timestamp 25201
transform 1 0 58144 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_617
timestamp 25201
transform 1 0 58788 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_626
timestamp 1636993656
transform 1 0 59616 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 25201
transform 1 0 63204 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 25201
transform 1 0 63756 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_673
timestamp 25201
transform 1 0 63940 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_709
timestamp 25201
transform 1 0 67252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_732
timestamp 25201
transform 1 0 69368 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_757
timestamp 25201
transform 1 0 71668 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_774
timestamp 25201
transform 1 0 73232 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_782
timestamp 25201
transform 1 0 73968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_820
timestamp 25201
transform 1 0 77464 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636993656
transform 1 0 2300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636993656
transform 1 0 3404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 25201
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 25201
transform 1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 25201
transform 1 0 5060 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp 25201
transform 1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 25201
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 25201
transform 1 0 14996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_192
timestamp 25201
transform 1 0 19688 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_325
timestamp 25201
transform 1 0 31924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_387
timestamp 25201
transform 1 0 37628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 25201
transform 1 0 45632 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 25201
transform 1 0 50324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 25201
transform 1 0 50876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_533
timestamp 25201
transform 1 0 51060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_539
timestamp 25201
transform 1 0 51612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_580
timestamp 25201
transform 1 0 55384 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636993656
transform 1 0 56212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_601
timestamp 25201
transform 1 0 57316 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_626
timestamp 1636993656
transform 1 0 59616 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_638
timestamp 25201
transform 1 0 60720 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_669
timestamp 25201
transform 1 0 63572 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_677
timestamp 25201
transform 1 0 64308 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_694
timestamp 25201
transform 1 0 65872 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_701
timestamp 25201
transform 1 0 66516 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_707
timestamp 25201
transform 1 0 67068 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_748
timestamp 25201
transform 1 0 70840 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_781
timestamp 25201
transform 1 0 73876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_787
timestamp 25201
transform 1 0 74428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_813
timestamp 25201
transform 1 0 76820 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636993656
transform 1 0 2300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636993656
transform 1 0 3404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636993656
transform 1 0 4508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_39
timestamp 25201
transform 1 0 5612 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 25201
transform 1 0 7268 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_140
timestamp 25201
transform 1 0 14904 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_158
timestamp 25201
transform 1 0 16560 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_240
timestamp 25201
transform 1 0 24104 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_364
timestamp 25201
transform 1 0 35512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_393
timestamp 25201
transform 1 0 38180 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_521
timestamp 1636993656
transform 1 0 49956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_533
timestamp 25201
transform 1 0 51060 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_541
timestamp 25201
transform 1 0 51796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_552
timestamp 25201
transform 1 0 52808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_561
timestamp 25201
transform 1 0 53636 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_570
timestamp 1636993656
transform 1 0 54464 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_582
timestamp 1636993656
transform 1 0 55568 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_594
timestamp 1636993656
transform 1 0 56672 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_606
timestamp 25201
transform 1 0 57776 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_614
timestamp 25201
transform 1 0 58512 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636993656
transform 1 0 58788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636993656
transform 1 0 59892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636993656
transform 1 0 60996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636993656
transform 1 0 62100 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 25201
transform 1 0 63204 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 25201
transform 1 0 63756 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636993656
transform 1 0 63940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_685
timestamp 25201
transform 1 0 65044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_689
timestamp 25201
transform 1 0 65412 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_698
timestamp 1636993656
transform 1 0 66240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_710
timestamp 25201
transform 1 0 67344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_720
timestamp 25201
transform 1 0 68264 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_729
timestamp 25201
transform 1 0 69092 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_738
timestamp 1636993656
transform 1 0 69920 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_750
timestamp 25201
transform 1 0 71024 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_762
timestamp 1636993656
transform 1 0 72128 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_774
timestamp 25201
transform 1 0 73232 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_782
timestamp 25201
transform 1 0 73968 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_785
timestamp 25201
transform 1 0 74244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_789
timestamp 25201
transform 1 0 74612 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636993656
transform 1 0 2300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636993656
transform 1 0 3404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 25201
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636993656
transform 1 0 4692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp 25201
transform 1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 25201
transform 1 0 9844 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 25201
transform 1 0 14996 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 25201
transform 1 0 19872 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 25201
transform 1 0 20148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_241
timestamp 25201
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 25201
transform 1 0 25116 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp 25201
transform 1 0 25300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_280
timestamp 25201
transform 1 0 27784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_290
timestamp 25201
transform 1 0 28704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 25201
transform 1 0 30452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_429
timestamp 25201
transform 1 0 41492 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_439
timestamp 25201
transform 1 0 42412 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 25201
transform 1 0 45724 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_517
timestamp 1636993656
transform 1 0 49588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_529
timestamp 25201
transform 1 0 50692 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636993656
transform 1 0 51060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636993656
transform 1 0 52164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1636993656
transform 1 0 53268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1636993656
transform 1 0 54372 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 25201
transform 1 0 55476 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 25201
transform 1 0 56028 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636993656
transform 1 0 56212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636993656
transform 1 0 57316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1636993656
transform 1 0 58420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1636993656
transform 1 0 59524 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 25201
transform 1 0 60628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 25201
transform 1 0 61180 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636993656
transform 1 0 61364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636993656
transform 1 0 62468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1636993656
transform 1 0 63572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1636993656
transform 1 0 64676 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 25201
transform 1 0 65780 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 25201
transform 1 0 66332 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636993656
transform 1 0 66516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636993656
transform 1 0 67620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1636993656
transform 1 0 68724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1636993656
transform 1 0 69828 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 25201
transform 1 0 70932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 25201
transform 1 0 71484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636993656
transform 1 0 71668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636993656
transform 1 0 72772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1636993656
transform 1 0 73876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1636993656
transform 1 0 74980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 25201
transform 1 0 76084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 25201
transform 1 0 76636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_813
timestamp 25201
transform 1 0 76820 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636993656
transform 1 0 2300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636993656
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636993656
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636993656
transform 1 0 5612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 25201
transform 1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 25201
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 25201
transform 1 0 7268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_116
timestamp 25201
transform 1 0 12696 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_308
timestamp 25201
transform 1 0 30360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 25201
transform 1 0 43056 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 25201
transform 1 0 47748 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 25201
transform 1 0 48300 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1636993656
transform 1 0 48484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1636993656
transform 1 0 49588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1636993656
transform 1 0 50692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1636993656
transform 1 0 51796 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 25201
transform 1 0 52900 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 25201
transform 1 0 53452 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1636993656
transform 1 0 53636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1636993656
transform 1 0 54740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1636993656
transform 1 0 55844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1636993656
transform 1 0 56948 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 25201
transform 1 0 58052 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 25201
transform 1 0 58604 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1636993656
transform 1 0 58788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1636993656
transform 1 0 59892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1636993656
transform 1 0 60996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1636993656
transform 1 0 62100 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 25201
transform 1 0 63204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 25201
transform 1 0 63756 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1636993656
transform 1 0 63940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1636993656
transform 1 0 65044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1636993656
transform 1 0 66148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1636993656
transform 1 0 67252 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 25201
transform 1 0 68356 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 25201
transform 1 0 68908 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1636993656
transform 1 0 69092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1636993656
transform 1 0 70196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1636993656
transform 1 0 71300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1636993656
transform 1 0 72404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 25201
transform 1 0 73508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 25201
transform 1 0 74060 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1636993656
transform 1 0 74244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1636993656
transform 1 0 75348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_809
timestamp 25201
transform 1 0 76452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_813
timestamp 25201
transform 1 0 76820 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636993656
transform 1 0 2300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636993656
transform 1 0 3404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 25201
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636993656
transform 1 0 4692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636993656
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_53
timestamp 25201
transform 1 0 6900 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_61
timestamp 25201
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 25201
transform 1 0 8648 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 25201
transform 1 0 9844 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 25201
transform 1 0 14996 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 25201
transform 1 0 45172 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 25201
transform 1 0 45724 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_485
timestamp 1636993656
transform 1 0 46644 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_497
timestamp 1636993656
transform 1 0 47748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_509
timestamp 1636993656
transform 1 0 48852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_521
timestamp 25201
transform 1 0 49956 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_529
timestamp 25201
transform 1 0 50692 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1636993656
transform 1 0 51060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1636993656
transform 1 0 52164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1636993656
transform 1 0 53268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1636993656
transform 1 0 54372 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 25201
transform 1 0 55476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 25201
transform 1 0 56028 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1636993656
transform 1 0 56212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1636993656
transform 1 0 57316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1636993656
transform 1 0 58420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1636993656
transform 1 0 59524 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 25201
transform 1 0 60628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 25201
transform 1 0 61180 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1636993656
transform 1 0 61364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1636993656
transform 1 0 62468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1636993656
transform 1 0 63572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1636993656
transform 1 0 64676 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 25201
transform 1 0 65780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 25201
transform 1 0 66332 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1636993656
transform 1 0 66516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1636993656
transform 1 0 67620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1636993656
transform 1 0 68724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1636993656
transform 1 0 69828 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 25201
transform 1 0 70932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 25201
transform 1 0 71484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1636993656
transform 1 0 71668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1636993656
transform 1 0 72772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1636993656
transform 1 0 73876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1636993656
transform 1 0 74980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 25201
transform 1 0 76084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 25201
transform 1 0 76636 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_813
timestamp 25201
transform 1 0 76820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_821
timestamp 25201
transform 1 0 77556 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636993656
transform 1 0 2300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636993656
transform 1 0 3404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636993656
transform 1 0 4508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636993656
transform 1 0 5612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 25201
transform 1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 25201
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636993656
transform 1 0 7268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_69
timestamp 25201
transform 1 0 8372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_75
timestamp 25201
transform 1 0 8924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_119
timestamp 25201
transform 1 0 12972 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 25201
transform 1 0 17572 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 25201
transform 1 0 22724 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_268
timestamp 25201
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 25201
transform 1 0 27692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 25201
transform 1 0 32844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_374
timestamp 25201
transform 1 0 36432 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_416
timestamp 25201
transform 1 0 40296 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_465
timestamp 1636993656
transform 1 0 44804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_477
timestamp 1636993656
transform 1 0 45908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_489
timestamp 1636993656
transform 1 0 47012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_501
timestamp 25201
transform 1 0 48116 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1636993656
transform 1 0 48484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1636993656
transform 1 0 49588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1636993656
transform 1 0 50692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1636993656
transform 1 0 51796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 25201
transform 1 0 52900 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 25201
transform 1 0 53452 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1636993656
transform 1 0 53636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1636993656
transform 1 0 54740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1636993656
transform 1 0 55844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1636993656
transform 1 0 56948 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 25201
transform 1 0 58052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 25201
transform 1 0 58604 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1636993656
transform 1 0 58788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1636993656
transform 1 0 59892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1636993656
transform 1 0 60996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1636993656
transform 1 0 62100 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 25201
transform 1 0 63204 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 25201
transform 1 0 63756 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1636993656
transform 1 0 63940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1636993656
transform 1 0 65044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1636993656
transform 1 0 66148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1636993656
transform 1 0 67252 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 25201
transform 1 0 68356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 25201
transform 1 0 68908 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1636993656
transform 1 0 69092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1636993656
transform 1 0 70196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1636993656
transform 1 0 71300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1636993656
transform 1 0 72404 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 25201
transform 1 0 73508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 25201
transform 1 0 74060 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1636993656
transform 1 0 74244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1636993656
transform 1 0 75348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1636993656
transform 1 0 76452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_821
timestamp 25201
transform 1 0 77556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636993656
transform 1 0 2300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636993656
transform 1 0 3404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 25201
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636993656
transform 1 0 4692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636993656
transform 1 0 5796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636993656
transform 1 0 6900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636993656
transform 1 0 8004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 25201
transform 1 0 9108 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 25201
transform 1 0 9660 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_88
timestamp 25201
transform 1 0 10120 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_96
timestamp 25201
transform 1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_107
timestamp 25201
transform 1 0 11868 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 25201
transform 1 0 19688 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_225
timestamp 25201
transform 1 0 22724 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_242
timestamp 25201
transform 1 0 24288 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_291
timestamp 25201
transform 1 0 28796 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 25201
transform 1 0 30452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_327
timestamp 25201
transform 1 0 32108 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_331
timestamp 25201
transform 1 0 32476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_384
timestamp 25201
transform 1 0 37352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_416
timestamp 25201
transform 1 0 40296 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1636993656
transform 1 0 42964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1636993656
transform 1 0 44068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 25201
transform 1 0 45172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 25201
transform 1 0 45724 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1636993656
transform 1 0 45908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1636993656
transform 1 0 47012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1636993656
transform 1 0 48116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1636993656
transform 1 0 49220 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 25201
transform 1 0 50324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 25201
transform 1 0 50876 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1636993656
transform 1 0 51060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1636993656
transform 1 0 52164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1636993656
transform 1 0 53268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1636993656
transform 1 0 54372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 25201
transform 1 0 55476 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 25201
transform 1 0 56028 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1636993656
transform 1 0 56212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1636993656
transform 1 0 57316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1636993656
transform 1 0 58420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1636993656
transform 1 0 59524 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 25201
transform 1 0 60628 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 25201
transform 1 0 61180 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1636993656
transform 1 0 61364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1636993656
transform 1 0 62468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1636993656
transform 1 0 63572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1636993656
transform 1 0 64676 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 25201
transform 1 0 65780 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 25201
transform 1 0 66332 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1636993656
transform 1 0 66516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1636993656
transform 1 0 67620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1636993656
transform 1 0 68724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1636993656
transform 1 0 69828 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 25201
transform 1 0 70932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 25201
transform 1 0 71484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1636993656
transform 1 0 71668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1636993656
transform 1 0 72772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1636993656
transform 1 0 73876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1636993656
transform 1 0 74980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 25201
transform 1 0 76084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 25201
transform 1 0 76636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_813
timestamp 25201
transform 1 0 76820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_821
timestamp 25201
transform 1 0 77556 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636993656
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636993656
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636993656
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636993656
transform 1 0 5612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 25201
transform 1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 25201
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636993656
transform 1 0 7268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636993656
transform 1 0 8372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636993656
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_93
timestamp 25201
transform 1 0 10580 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 25201
transform 1 0 11132 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 25201
transform 1 0 11960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 25201
transform 1 0 12420 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 25201
transform 1 0 22724 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_229
timestamp 25201
transform 1 0 23092 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_238
timestamp 25201
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_281
timestamp 25201
transform 1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_300
timestamp 25201
transform 1 0 29624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_417
timestamp 25201
transform 1 0 40388 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_443
timestamp 25201
transform 1 0 42780 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 25201
transform 1 0 43148 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1636993656
transform 1 0 43332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1636993656
transform 1 0 44436 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1636993656
transform 1 0 45540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1636993656
transform 1 0 46644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 25201
transform 1 0 47748 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 25201
transform 1 0 48300 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1636993656
transform 1 0 48484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1636993656
transform 1 0 49588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1636993656
transform 1 0 50692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1636993656
transform 1 0 51796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 25201
transform 1 0 52900 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 25201
transform 1 0 53452 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1636993656
transform 1 0 53636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1636993656
transform 1 0 54740 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1636993656
transform 1 0 55844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1636993656
transform 1 0 56948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 25201
transform 1 0 58052 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 25201
transform 1 0 58604 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1636993656
transform 1 0 58788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1636993656
transform 1 0 59892 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1636993656
transform 1 0 60996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1636993656
transform 1 0 62100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 25201
transform 1 0 63204 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 25201
transform 1 0 63756 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1636993656
transform 1 0 63940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1636993656
transform 1 0 65044 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1636993656
transform 1 0 66148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1636993656
transform 1 0 67252 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 25201
transform 1 0 68356 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 25201
transform 1 0 68908 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1636993656
transform 1 0 69092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1636993656
transform 1 0 70196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_753
timestamp 1636993656
transform 1 0 71300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_765
timestamp 1636993656
transform 1 0 72404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 25201
transform 1 0 73508 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 25201
transform 1 0 74060 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1636993656
transform 1 0 74244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1636993656
transform 1 0 75348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_809
timestamp 1636993656
transform 1 0 76452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_821
timestamp 25201
transform 1 0 77556 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636993656
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636993656
transform 1 0 3404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 25201
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636993656
transform 1 0 4692 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636993656
transform 1 0 5796 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636993656
transform 1 0 6900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1636993656
transform 1 0 8004 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 25201
transform 1 0 9108 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 25201
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636993656
transform 1 0 9844 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636993656
transform 1 0 10948 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636993656
transform 1 0 12052 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_121
timestamp 25201
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_129
timestamp 25201
transform 1 0 13892 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 25201
transform 1 0 14812 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_147
timestamp 25201
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_322
timestamp 25201
transform 1 0 31648 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_326
timestamp 25201
transform 1 0 32016 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_368
timestamp 25201
transform 1 0 35880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 25201
transform 1 0 40296 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_435
timestamp 1636993656
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_447
timestamp 1636993656
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_459
timestamp 1636993656
transform 1 0 44252 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_471
timestamp 25201
transform 1 0 45356 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 25201
transform 1 0 45724 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1636993656
transform 1 0 45908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1636993656
transform 1 0 47012 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1636993656
transform 1 0 48116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1636993656
transform 1 0 49220 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 25201
transform 1 0 50324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 25201
transform 1 0 50876 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1636993656
transform 1 0 51060 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1636993656
transform 1 0 52164 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1636993656
transform 1 0 53268 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1636993656
transform 1 0 54372 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 25201
transform 1 0 55476 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 25201
transform 1 0 56028 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1636993656
transform 1 0 56212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1636993656
transform 1 0 57316 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1636993656
transform 1 0 58420 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1636993656
transform 1 0 59524 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 25201
transform 1 0 60628 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 25201
transform 1 0 61180 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1636993656
transform 1 0 61364 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1636993656
transform 1 0 62468 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1636993656
transform 1 0 63572 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1636993656
transform 1 0 64676 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 25201
transform 1 0 65780 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 25201
transform 1 0 66332 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1636993656
transform 1 0 66516 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1636993656
transform 1 0 67620 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_725
timestamp 1636993656
transform 1 0 68724 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_737
timestamp 1636993656
transform 1 0 69828 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 25201
transform 1 0 70932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 25201
transform 1 0 71484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1636993656
transform 1 0 71668 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_769
timestamp 1636993656
transform 1 0 72772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_781
timestamp 1636993656
transform 1 0 73876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_793
timestamp 1636993656
transform 1 0 74980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 25201
transform 1 0 76084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 25201
transform 1 0 76636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_813
timestamp 25201
transform 1 0 76820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_821
timestamp 25201
transform 1 0 77556 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636993656
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636993656
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636993656
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636993656
transform 1 0 5612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 25201
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 25201
transform 1 0 7084 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636993656
transform 1 0 7268 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1636993656
transform 1 0 8372 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1636993656
transform 1 0 9476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1636993656
transform 1 0 10580 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 25201
transform 1 0 11684 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 25201
transform 1 0 12236 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1636993656
transform 1 0 12420 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1636993656
transform 1 0 13524 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1636993656
transform 1 0 14628 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_149
timestamp 25201
transform 1 0 15732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp 25201
transform 1 0 17572 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_229
timestamp 25201
transform 1 0 23092 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_345
timestamp 25201
transform 1 0 33764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_356
timestamp 25201
transform 1 0 34776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 25201
transform 1 0 37720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_403
timestamp 25201
transform 1 0 39100 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_420
timestamp 1636993656
transform 1 0 40664 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_432
timestamp 1636993656
transform 1 0 41768 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_444
timestamp 25201
transform 1 0 42872 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1636993656
transform 1 0 43332 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1636993656
transform 1 0 44436 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1636993656
transform 1 0 45540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1636993656
transform 1 0 46644 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 25201
transform 1 0 47748 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 25201
transform 1 0 48300 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1636993656
transform 1 0 48484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1636993656
transform 1 0 49588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1636993656
transform 1 0 50692 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1636993656
transform 1 0 51796 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 25201
transform 1 0 52900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 25201
transform 1 0 53452 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1636993656
transform 1 0 53636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1636993656
transform 1 0 54740 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1636993656
transform 1 0 55844 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1636993656
transform 1 0 56948 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 25201
transform 1 0 58052 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 25201
transform 1 0 58604 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1636993656
transform 1 0 58788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1636993656
transform 1 0 59892 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1636993656
transform 1 0 60996 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1636993656
transform 1 0 62100 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 25201
transform 1 0 63204 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 25201
transform 1 0 63756 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1636993656
transform 1 0 63940 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1636993656
transform 1 0 65044 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1636993656
transform 1 0 66148 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1636993656
transform 1 0 67252 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 25201
transform 1 0 68356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 25201
transform 1 0 68908 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_729
timestamp 1636993656
transform 1 0 69092 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_741
timestamp 1636993656
transform 1 0 70196 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1636993656
transform 1 0 71300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1636993656
transform 1 0 72404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 25201
transform 1 0 73508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 25201
transform 1 0 74060 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_785
timestamp 1636993656
transform 1 0 74244 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_797
timestamp 1636993656
transform 1 0 75348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_809
timestamp 1636993656
transform 1 0 76452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_821
timestamp 25201
transform 1 0 77556 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636993656
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636993656
transform 1 0 3404 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 25201
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636993656
transform 1 0 4692 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636993656
transform 1 0 5796 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636993656
transform 1 0 6900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1636993656
transform 1 0 8004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 25201
transform 1 0 9108 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 25201
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1636993656
transform 1 0 9844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_97
timestamp 25201
transform 1 0 10948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_103
timestamp 25201
transform 1 0 11500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_107
timestamp 1636993656
transform 1 0 11868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_119
timestamp 1636993656
transform 1 0 12972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_131
timestamp 25201
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 25201
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_141
timestamp 25201
transform 1 0 14996 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 25201
transform 1 0 15732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_159
timestamp 25201
transform 1 0 16652 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_163
timestamp 25201
transform 1 0 17020 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 25201
transform 1 0 20148 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_280
timestamp 25201
transform 1 0 27784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_290
timestamp 25201
transform 1 0 28704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_309
timestamp 25201
transform 1 0 30452 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_324
timestamp 25201
transform 1 0 31832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_336
timestamp 25201
transform 1 0 32936 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_394
timestamp 25201
transform 1 0 38272 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_398
timestamp 25201
transform 1 0 38640 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_415
timestamp 25201
transform 1 0 40204 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 25201
transform 1 0 40572 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1636993656
transform 1 0 40756 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1636993656
transform 1 0 41860 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1636993656
transform 1 0 42964 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1636993656
transform 1 0 44068 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 25201
transform 1 0 45172 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 25201
transform 1 0 45724 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1636993656
transform 1 0 45908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1636993656
transform 1 0 47012 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1636993656
transform 1 0 48116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1636993656
transform 1 0 49220 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 25201
transform 1 0 50324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 25201
transform 1 0 50876 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1636993656
transform 1 0 51060 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1636993656
transform 1 0 52164 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1636993656
transform 1 0 53268 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1636993656
transform 1 0 54372 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 25201
transform 1 0 55476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 25201
transform 1 0 56028 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1636993656
transform 1 0 56212 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1636993656
transform 1 0 57316 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1636993656
transform 1 0 58420 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1636993656
transform 1 0 59524 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 25201
transform 1 0 60628 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 25201
transform 1 0 61180 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1636993656
transform 1 0 61364 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1636993656
transform 1 0 62468 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1636993656
transform 1 0 63572 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1636993656
transform 1 0 64676 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 25201
transform 1 0 65780 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 25201
transform 1 0 66332 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1636993656
transform 1 0 66516 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1636993656
transform 1 0 67620 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_725
timestamp 1636993656
transform 1 0 68724 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_737
timestamp 1636993656
transform 1 0 69828 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 25201
transform 1 0 70932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 25201
transform 1 0 71484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1636993656
transform 1 0 71668 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1636993656
transform 1 0 72772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1636993656
transform 1 0 73876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_793
timestamp 1636993656
transform 1 0 74980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 25201
transform 1 0 76084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 25201
transform 1 0 76636 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_813
timestamp 25201
transform 1 0 76820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_821
timestamp 25201
transform 1 0 77556 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636993656
transform 1 0 2300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636993656
transform 1 0 3404 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636993656
transform 1 0 4508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636993656
transform 1 0 5612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 25201
transform 1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 25201
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636993656
transform 1 0 7268 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1636993656
transform 1 0 8372 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1636993656
transform 1 0 9476 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1636993656
transform 1 0 10580 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 25201
transform 1 0 11684 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 25201
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1636993656
transform 1 0 12420 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1636993656
transform 1 0 13524 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1636993656
transform 1 0 14628 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1636993656
transform 1 0 15732 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 25201
transform 1 0 16836 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 25201
transform 1 0 17388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 25201
transform 1 0 17572 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_177
timestamp 25201
transform 1 0 18308 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_204
timestamp 25201
transform 1 0 20792 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 25201
transform 1 0 22724 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 25201
transform 1 0 24380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_281
timestamp 25201
transform 1 0 27876 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 25201
transform 1 0 32568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_337
timestamp 25201
transform 1 0 33028 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_401
timestamp 1636993656
transform 1 0 38916 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_413
timestamp 1636993656
transform 1 0 40020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_425
timestamp 1636993656
transform 1 0 41124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_437
timestamp 25201
transform 1 0 42228 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_445
timestamp 25201
transform 1 0 42964 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1636993656
transform 1 0 43332 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1636993656
transform 1 0 44436 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1636993656
transform 1 0 45540 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1636993656
transform 1 0 46644 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 25201
transform 1 0 47748 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 25201
transform 1 0 48300 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1636993656
transform 1 0 48484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1636993656
transform 1 0 49588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1636993656
transform 1 0 50692 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1636993656
transform 1 0 51796 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 25201
transform 1 0 52900 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 25201
transform 1 0 53452 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1636993656
transform 1 0 53636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1636993656
transform 1 0 54740 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1636993656
transform 1 0 55844 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1636993656
transform 1 0 56948 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 25201
transform 1 0 58052 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 25201
transform 1 0 58604 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1636993656
transform 1 0 58788 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1636993656
transform 1 0 59892 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1636993656
transform 1 0 60996 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1636993656
transform 1 0 62100 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 25201
transform 1 0 63204 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 25201
transform 1 0 63756 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1636993656
transform 1 0 63940 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1636993656
transform 1 0 65044 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1636993656
transform 1 0 66148 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1636993656
transform 1 0 67252 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 25201
transform 1 0 68356 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 25201
transform 1 0 68908 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_729
timestamp 1636993656
transform 1 0 69092 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_741
timestamp 1636993656
transform 1 0 70196 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_753
timestamp 1636993656
transform 1 0 71300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_765
timestamp 1636993656
transform 1 0 72404 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 25201
transform 1 0 73508 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 25201
transform 1 0 74060 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_785
timestamp 1636993656
transform 1 0 74244 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_797
timestamp 1636993656
transform 1 0 75348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_809
timestamp 1636993656
transform 1 0 76452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_821
timestamp 25201
transform 1 0 77556 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636993656
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636993656
transform 1 0 3404 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 25201
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636993656
transform 1 0 4692 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636993656
transform 1 0 5796 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636993656
transform 1 0 6900 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1636993656
transform 1 0 8004 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 25201
transform 1 0 9108 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 25201
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636993656
transform 1 0 9844 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1636993656
transform 1 0 10948 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1636993656
transform 1 0 12052 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1636993656
transform 1 0 13156 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 25201
transform 1 0 14260 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 25201
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1636993656
transform 1 0 14996 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1636993656
transform 1 0 16100 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1636993656
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1636993656
transform 1 0 18308 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 25201
transform 1 0 19964 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 25201
transform 1 0 20148 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_203
timestamp 25201
transform 1 0 20700 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_220
timestamp 25201
transform 1 0 22264 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 25201
transform 1 0 25116 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_253
timestamp 25201
transform 1 0 25300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_274
timestamp 25201
transform 1 0 27232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_309
timestamp 25201
transform 1 0 30452 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_320
timestamp 25201
transform 1 0 31464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_334
timestamp 25201
transform 1 0 32752 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 25201
transform 1 0 35052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 25201
transform 1 0 35420 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_365
timestamp 25201
transform 1 0 35604 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_384
timestamp 1636993656
transform 1 0 37352 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_396
timestamp 1636993656
transform 1 0 38456 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_408
timestamp 1636993656
transform 1 0 39560 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1636993656
transform 1 0 40756 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1636993656
transform 1 0 41860 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1636993656
transform 1 0 42964 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1636993656
transform 1 0 44068 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 25201
transform 1 0 45172 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 25201
transform 1 0 45724 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1636993656
transform 1 0 45908 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1636993656
transform 1 0 47012 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1636993656
transform 1 0 48116 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1636993656
transform 1 0 49220 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 25201
transform 1 0 50324 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 25201
transform 1 0 50876 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1636993656
transform 1 0 51060 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1636993656
transform 1 0 52164 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1636993656
transform 1 0 53268 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1636993656
transform 1 0 54372 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 25201
transform 1 0 55476 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 25201
transform 1 0 56028 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1636993656
transform 1 0 56212 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1636993656
transform 1 0 57316 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1636993656
transform 1 0 58420 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1636993656
transform 1 0 59524 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 25201
transform 1 0 60628 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 25201
transform 1 0 61180 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1636993656
transform 1 0 61364 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1636993656
transform 1 0 62468 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1636993656
transform 1 0 63572 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1636993656
transform 1 0 64676 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 25201
transform 1 0 65780 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 25201
transform 1 0 66332 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1636993656
transform 1 0 66516 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1636993656
transform 1 0 67620 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_725
timestamp 1636993656
transform 1 0 68724 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_737
timestamp 1636993656
transform 1 0 69828 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 25201
transform 1 0 70932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 25201
transform 1 0 71484 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_757
timestamp 1636993656
transform 1 0 71668 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_769
timestamp 1636993656
transform 1 0 72772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_781
timestamp 1636993656
transform 1 0 73876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_793
timestamp 1636993656
transform 1 0 74980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 25201
transform 1 0 76084 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 25201
transform 1 0 76636 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_813
timestamp 25201
transform 1 0 76820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_821
timestamp 25201
transform 1 0 77556 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636993656
transform 1 0 2300 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636993656
transform 1 0 3404 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636993656
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636993656
transform 1 0 5612 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 25201
transform 1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 25201
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636993656
transform 1 0 7268 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1636993656
transform 1 0 8372 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1636993656
transform 1 0 9476 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1636993656
transform 1 0 10580 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 25201
transform 1 0 11684 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 25201
transform 1 0 12236 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1636993656
transform 1 0 12420 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1636993656
transform 1 0 13524 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1636993656
transform 1 0 14628 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1636993656
transform 1 0 15732 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 25201
transform 1 0 16836 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 25201
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1636993656
transform 1 0 17572 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1636993656
transform 1 0 18676 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_193
timestamp 25201
transform 1 0 19780 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_210
timestamp 25201
transform 1 0 21344 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 25201
transform 1 0 22540 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_254
timestamp 25201
transform 1 0 25392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_271
timestamp 25201
transform 1 0 26956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_284
timestamp 25201
transform 1 0 28152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_311
timestamp 25201
transform 1 0 30636 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_316
timestamp 25201
transform 1 0 31096 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_339
timestamp 25201
transform 1 0 33212 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_366
timestamp 1636993656
transform 1 0 35696 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_378
timestamp 1636993656
transform 1 0 36800 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 25201
transform 1 0 37904 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1636993656
transform 1 0 38180 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1636993656
transform 1 0 39284 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1636993656
transform 1 0 40388 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1636993656
transform 1 0 41492 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 25201
transform 1 0 42596 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 25201
transform 1 0 43148 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1636993656
transform 1 0 43332 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1636993656
transform 1 0 44436 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1636993656
transform 1 0 45540 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1636993656
transform 1 0 46644 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 25201
transform 1 0 47748 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 25201
transform 1 0 48300 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1636993656
transform 1 0 48484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1636993656
transform 1 0 49588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1636993656
transform 1 0 50692 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1636993656
transform 1 0 51796 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 25201
transform 1 0 52900 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 25201
transform 1 0 53452 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1636993656
transform 1 0 53636 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1636993656
transform 1 0 54740 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1636993656
transform 1 0 55844 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1636993656
transform 1 0 56948 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 25201
transform 1 0 58052 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 25201
transform 1 0 58604 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1636993656
transform 1 0 58788 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1636993656
transform 1 0 59892 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1636993656
transform 1 0 60996 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1636993656
transform 1 0 62100 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 25201
transform 1 0 63204 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 25201
transform 1 0 63756 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1636993656
transform 1 0 63940 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1636993656
transform 1 0 65044 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1636993656
transform 1 0 66148 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1636993656
transform 1 0 67252 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 25201
transform 1 0 68356 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 25201
transform 1 0 68908 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_729
timestamp 1636993656
transform 1 0 69092 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_741
timestamp 1636993656
transform 1 0 70196 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_753
timestamp 1636993656
transform 1 0 71300 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_765
timestamp 1636993656
transform 1 0 72404 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 25201
transform 1 0 73508 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 25201
transform 1 0 74060 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_785
timestamp 1636993656
transform 1 0 74244 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_797
timestamp 1636993656
transform 1 0 75348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_809
timestamp 1636993656
transform 1 0 76452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_821
timestamp 25201
transform 1 0 77556 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636993656
transform 1 0 2300 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636993656
transform 1 0 3404 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 25201
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636993656
transform 1 0 4692 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636993656
transform 1 0 5796 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636993656
transform 1 0 6900 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1636993656
transform 1 0 8004 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 25201
transform 1 0 9108 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 25201
transform 1 0 9660 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636993656
transform 1 0 9844 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1636993656
transform 1 0 10948 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1636993656
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1636993656
transform 1 0 13156 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 25201
transform 1 0 14260 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 25201
transform 1 0 14812 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636993656
transform 1 0 14996 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1636993656
transform 1 0 16100 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1636993656
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1636993656
transform 1 0 18308 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 25201
transform 1 0 19412 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 25201
transform 1 0 19964 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1636993656
transform 1 0 20148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 25201
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 25201
transform 1 0 21620 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_289
timestamp 25201
transform 1 0 28612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 25201
transform 1 0 30268 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_309
timestamp 25201
transform 1 0 30452 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_320
timestamp 25201
transform 1 0 31464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_330
timestamp 25201
transform 1 0 32384 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_336
timestamp 25201
transform 1 0 32936 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_359
timestamp 25201
transform 1 0 35052 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 25201
transform 1 0 35420 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1636993656
transform 1 0 35604 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1636993656
transform 1 0 36708 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1636993656
transform 1 0 37812 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1636993656
transform 1 0 38916 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 25201
transform 1 0 40020 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 25201
transform 1 0 40572 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1636993656
transform 1 0 40756 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1636993656
transform 1 0 41860 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1636993656
transform 1 0 42964 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1636993656
transform 1 0 44068 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 25201
transform 1 0 45172 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 25201
transform 1 0 45724 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1636993656
transform 1 0 45908 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1636993656
transform 1 0 47012 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1636993656
transform 1 0 48116 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1636993656
transform 1 0 49220 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 25201
transform 1 0 50324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 25201
transform 1 0 50876 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1636993656
transform 1 0 51060 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1636993656
transform 1 0 52164 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1636993656
transform 1 0 53268 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1636993656
transform 1 0 54372 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 25201
transform 1 0 55476 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 25201
transform 1 0 56028 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1636993656
transform 1 0 56212 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1636993656
transform 1 0 57316 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1636993656
transform 1 0 58420 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1636993656
transform 1 0 59524 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 25201
transform 1 0 60628 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 25201
transform 1 0 61180 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1636993656
transform 1 0 61364 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1636993656
transform 1 0 62468 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1636993656
transform 1 0 63572 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1636993656
transform 1 0 64676 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 25201
transform 1 0 65780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 25201
transform 1 0 66332 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1636993656
transform 1 0 66516 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1636993656
transform 1 0 67620 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_725
timestamp 1636993656
transform 1 0 68724 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_737
timestamp 1636993656
transform 1 0 69828 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 25201
transform 1 0 70932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 25201
transform 1 0 71484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_757
timestamp 1636993656
transform 1 0 71668 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_769
timestamp 1636993656
transform 1 0 72772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_781
timestamp 1636993656
transform 1 0 73876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_793
timestamp 1636993656
transform 1 0 74980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 25201
transform 1 0 76084 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 25201
transform 1 0 76636 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_813
timestamp 25201
transform 1 0 76820 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_821
timestamp 25201
transform 1 0 77556 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636993656
transform 1 0 2300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636993656
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1636993656
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1636993656
transform 1 0 5612 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 25201
transform 1 0 6716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 25201
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636993656
transform 1 0 7268 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636993656
transform 1 0 8372 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1636993656
transform 1 0 9476 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1636993656
transform 1 0 10580 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 25201
transform 1 0 11684 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 25201
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636993656
transform 1 0 12420 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1636993656
transform 1 0 13524 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1636993656
transform 1 0 14628 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1636993656
transform 1 0 15732 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 25201
transform 1 0 16836 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 25201
transform 1 0 17388 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636993656
transform 1 0 17572 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1636993656
transform 1 0 18676 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1636993656
transform 1 0 19780 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1636993656
transform 1 0 20884 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_217
timestamp 25201
transform 1 0 21988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 25201
transform 1 0 22540 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_227
timestamp 25201
transform 1 0 22908 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_238
timestamp 25201
transform 1 0 23920 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_254
timestamp 25201
transform 1 0 25392 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_260
timestamp 25201
transform 1 0 25944 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_266
timestamp 25201
transform 1 0 26496 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 25201
transform 1 0 27324 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 25201
transform 1 0 27692 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_281
timestamp 25201
transform 1 0 27876 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_301
timestamp 25201
transform 1 0 29716 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_315
timestamp 1636993656
transform 1 0 31004 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_327
timestamp 25201
transform 1 0 32108 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 25201
transform 1 0 32844 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_344
timestamp 1636993656
transform 1 0 33672 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_356
timestamp 1636993656
transform 1 0 34776 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_368
timestamp 1636993656
transform 1 0 35880 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_380
timestamp 1636993656
transform 1 0 36984 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1636993656
transform 1 0 38180 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1636993656
transform 1 0 39284 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1636993656
transform 1 0 40388 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1636993656
transform 1 0 41492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 25201
transform 1 0 42596 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 25201
transform 1 0 43148 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1636993656
transform 1 0 43332 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1636993656
transform 1 0 44436 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1636993656
transform 1 0 45540 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1636993656
transform 1 0 46644 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 25201
transform 1 0 47748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 25201
transform 1 0 48300 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1636993656
transform 1 0 48484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1636993656
transform 1 0 49588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1636993656
transform 1 0 50692 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1636993656
transform 1 0 51796 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 25201
transform 1 0 52900 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 25201
transform 1 0 53452 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1636993656
transform 1 0 53636 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1636993656
transform 1 0 54740 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1636993656
transform 1 0 55844 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1636993656
transform 1 0 56948 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 25201
transform 1 0 58052 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 25201
transform 1 0 58604 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1636993656
transform 1 0 58788 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1636993656
transform 1 0 59892 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1636993656
transform 1 0 60996 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1636993656
transform 1 0 62100 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 25201
transform 1 0 63204 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 25201
transform 1 0 63756 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1636993656
transform 1 0 63940 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1636993656
transform 1 0 65044 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1636993656
transform 1 0 66148 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1636993656
transform 1 0 67252 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 25201
transform 1 0 68356 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 25201
transform 1 0 68908 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_729
timestamp 1636993656
transform 1 0 69092 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_741
timestamp 1636993656
transform 1 0 70196 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_753
timestamp 1636993656
transform 1 0 71300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_765
timestamp 1636993656
transform 1 0 72404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 25201
transform 1 0 73508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 25201
transform 1 0 74060 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_785
timestamp 1636993656
transform 1 0 74244 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_797
timestamp 1636993656
transform 1 0 75348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_809
timestamp 1636993656
transform 1 0 76452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_821
timestamp 25201
transform 1 0 77556 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636993656
transform 1 0 2300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636993656
transform 1 0 3404 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 25201
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636993656
transform 1 0 4692 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636993656
transform 1 0 5796 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636993656
transform 1 0 6900 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1636993656
transform 1 0 8004 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 25201
transform 1 0 9108 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 25201
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636993656
transform 1 0 9844 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636993656
transform 1 0 10948 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1636993656
transform 1 0 12052 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1636993656
transform 1 0 13156 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 25201
transform 1 0 14260 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 25201
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636993656
transform 1 0 14996 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636993656
transform 1 0 16100 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1636993656
transform 1 0 17204 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1636993656
transform 1 0 18308 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 25201
transform 1 0 19412 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 25201
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1636993656
transform 1 0 20148 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1636993656
transform 1 0 21252 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1636993656
transform 1 0 22356 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1636993656
transform 1 0 23460 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 25201
transform 1 0 24564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 25201
transform 1 0 25116 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1636993656
transform 1 0 25300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1636993656
transform 1 0 26404 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1636993656
transform 1 0 27508 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1636993656
transform 1 0 28612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 25201
transform 1 0 29716 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 25201
transform 1 0 30268 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1636993656
transform 1 0 30452 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1636993656
transform 1 0 31556 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1636993656
transform 1 0 32660 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1636993656
transform 1 0 33764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 25201
transform 1 0 34868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 25201
transform 1 0 35420 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1636993656
transform 1 0 35604 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1636993656
transform 1 0 36708 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1636993656
transform 1 0 37812 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1636993656
transform 1 0 38916 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 25201
transform 1 0 40020 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 25201
transform 1 0 40572 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1636993656
transform 1 0 40756 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1636993656
transform 1 0 41860 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1636993656
transform 1 0 42964 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1636993656
transform 1 0 44068 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 25201
transform 1 0 45172 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 25201
transform 1 0 45724 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1636993656
transform 1 0 45908 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1636993656
transform 1 0 47012 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1636993656
transform 1 0 48116 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1636993656
transform 1 0 49220 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 25201
transform 1 0 50324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 25201
transform 1 0 50876 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1636993656
transform 1 0 51060 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1636993656
transform 1 0 52164 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1636993656
transform 1 0 53268 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1636993656
transform 1 0 54372 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 25201
transform 1 0 55476 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 25201
transform 1 0 56028 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1636993656
transform 1 0 56212 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1636993656
transform 1 0 57316 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1636993656
transform 1 0 58420 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1636993656
transform 1 0 59524 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 25201
transform 1 0 60628 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 25201
transform 1 0 61180 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1636993656
transform 1 0 61364 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1636993656
transform 1 0 62468 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1636993656
transform 1 0 63572 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1636993656
transform 1 0 64676 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 25201
transform 1 0 65780 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 25201
transform 1 0 66332 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1636993656
transform 1 0 66516 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1636993656
transform 1 0 67620 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_725
timestamp 1636993656
transform 1 0 68724 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_737
timestamp 1636993656
transform 1 0 69828 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 25201
transform 1 0 70932 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 25201
transform 1 0 71484 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_757
timestamp 1636993656
transform 1 0 71668 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_769
timestamp 1636993656
transform 1 0 72772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_781
timestamp 1636993656
transform 1 0 73876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_793
timestamp 1636993656
transform 1 0 74980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_805
timestamp 25201
transform 1 0 76084 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_811
timestamp 25201
transform 1 0 76636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_813
timestamp 25201
transform 1 0 76820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_821
timestamp 25201
transform 1 0 77556 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636993656
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636993656
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636993656
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1636993656
transform 1 0 5612 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 25201
transform 1 0 6716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 25201
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636993656
transform 1 0 7268 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1636993656
transform 1 0 8372 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1636993656
transform 1 0 9476 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1636993656
transform 1 0 10580 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 25201
transform 1 0 11684 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 25201
transform 1 0 12236 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636993656
transform 1 0 12420 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1636993656
transform 1 0 13524 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1636993656
transform 1 0 14628 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1636993656
transform 1 0 15732 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 25201
transform 1 0 16836 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 25201
transform 1 0 17388 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636993656
transform 1 0 17572 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1636993656
transform 1 0 18676 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1636993656
transform 1 0 19780 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1636993656
transform 1 0 20884 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 25201
transform 1 0 21988 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 25201
transform 1 0 22540 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636993656
transform 1 0 22724 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1636993656
transform 1 0 23828 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1636993656
transform 1 0 24932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1636993656
transform 1 0 26036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 25201
transform 1 0 27140 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 25201
transform 1 0 27692 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1636993656
transform 1 0 27876 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1636993656
transform 1 0 28980 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1636993656
transform 1 0 30084 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1636993656
transform 1 0 31188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 25201
transform 1 0 32292 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 25201
transform 1 0 32844 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1636993656
transform 1 0 33028 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1636993656
transform 1 0 34132 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1636993656
transform 1 0 35236 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1636993656
transform 1 0 36340 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 25201
transform 1 0 37444 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 25201
transform 1 0 37996 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1636993656
transform 1 0 38180 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1636993656
transform 1 0 39284 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1636993656
transform 1 0 40388 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1636993656
transform 1 0 41492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 25201
transform 1 0 42596 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 25201
transform 1 0 43148 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1636993656
transform 1 0 43332 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1636993656
transform 1 0 44436 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1636993656
transform 1 0 45540 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1636993656
transform 1 0 46644 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 25201
transform 1 0 47748 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 25201
transform 1 0 48300 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1636993656
transform 1 0 48484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1636993656
transform 1 0 49588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1636993656
transform 1 0 50692 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1636993656
transform 1 0 51796 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 25201
transform 1 0 52900 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 25201
transform 1 0 53452 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1636993656
transform 1 0 53636 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1636993656
transform 1 0 54740 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1636993656
transform 1 0 55844 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1636993656
transform 1 0 56948 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 25201
transform 1 0 58052 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 25201
transform 1 0 58604 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1636993656
transform 1 0 58788 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1636993656
transform 1 0 59892 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1636993656
transform 1 0 60996 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1636993656
transform 1 0 62100 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 25201
transform 1 0 63204 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 25201
transform 1 0 63756 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1636993656
transform 1 0 63940 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1636993656
transform 1 0 65044 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1636993656
transform 1 0 66148 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1636993656
transform 1 0 67252 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 25201
transform 1 0 68356 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 25201
transform 1 0 68908 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_729
timestamp 1636993656
transform 1 0 69092 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_741
timestamp 1636993656
transform 1 0 70196 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_753
timestamp 1636993656
transform 1 0 71300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_765
timestamp 1636993656
transform 1 0 72404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_777
timestamp 25201
transform 1 0 73508 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 25201
transform 1 0 74060 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_785
timestamp 1636993656
transform 1 0 74244 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_797
timestamp 1636993656
transform 1 0 75348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_809
timestamp 1636993656
transform 1 0 76452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_821
timestamp 25201
transform 1 0 77556 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636993656
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636993656
transform 1 0 3404 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 25201
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636993656
transform 1 0 4692 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636993656
transform 1 0 5796 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636993656
transform 1 0 6900 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1636993656
transform 1 0 8004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 25201
transform 1 0 9108 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 25201
transform 1 0 9660 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636993656
transform 1 0 9844 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1636993656
transform 1 0 10948 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1636993656
transform 1 0 12052 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1636993656
transform 1 0 13156 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 25201
transform 1 0 14260 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 25201
transform 1 0 14812 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1636993656
transform 1 0 14996 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1636993656
transform 1 0 16100 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1636993656
transform 1 0 17204 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1636993656
transform 1 0 18308 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 25201
transform 1 0 19412 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 25201
transform 1 0 19964 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1636993656
transform 1 0 20148 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1636993656
transform 1 0 21252 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1636993656
transform 1 0 22356 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1636993656
transform 1 0 23460 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 25201
transform 1 0 24564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 25201
transform 1 0 25116 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1636993656
transform 1 0 25300 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1636993656
transform 1 0 26404 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1636993656
transform 1 0 27508 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1636993656
transform 1 0 28612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 25201
transform 1 0 29716 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 25201
transform 1 0 30268 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1636993656
transform 1 0 30452 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1636993656
transform 1 0 31556 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1636993656
transform 1 0 32660 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1636993656
transform 1 0 33764 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 25201
transform 1 0 34868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 25201
transform 1 0 35420 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1636993656
transform 1 0 35604 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1636993656
transform 1 0 36708 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1636993656
transform 1 0 37812 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1636993656
transform 1 0 38916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 25201
transform 1 0 40020 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 25201
transform 1 0 40572 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1636993656
transform 1 0 40756 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1636993656
transform 1 0 41860 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1636993656
transform 1 0 42964 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1636993656
transform 1 0 44068 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 25201
transform 1 0 45172 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 25201
transform 1 0 45724 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1636993656
transform 1 0 45908 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1636993656
transform 1 0 47012 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1636993656
transform 1 0 48116 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1636993656
transform 1 0 49220 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 25201
transform 1 0 50324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 25201
transform 1 0 50876 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1636993656
transform 1 0 51060 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1636993656
transform 1 0 52164 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1636993656
transform 1 0 53268 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1636993656
transform 1 0 54372 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 25201
transform 1 0 55476 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 25201
transform 1 0 56028 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1636993656
transform 1 0 56212 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1636993656
transform 1 0 57316 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1636993656
transform 1 0 58420 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1636993656
transform 1 0 59524 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 25201
transform 1 0 60628 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 25201
transform 1 0 61180 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1636993656
transform 1 0 61364 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1636993656
transform 1 0 62468 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1636993656
transform 1 0 63572 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1636993656
transform 1 0 64676 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 25201
transform 1 0 65780 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 25201
transform 1 0 66332 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1636993656
transform 1 0 66516 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_713
timestamp 1636993656
transform 1 0 67620 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_725
timestamp 1636993656
transform 1 0 68724 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_737
timestamp 1636993656
transform 1 0 69828 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_749
timestamp 25201
transform 1 0 70932 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_755
timestamp 25201
transform 1 0 71484 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_757
timestamp 1636993656
transform 1 0 71668 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_769
timestamp 1636993656
transform 1 0 72772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_781
timestamp 1636993656
transform 1 0 73876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_793
timestamp 1636993656
transform 1 0 74980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_805
timestamp 25201
transform 1 0 76084 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_811
timestamp 25201
transform 1 0 76636 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_813
timestamp 25201
transform 1 0 76820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_821
timestamp 25201
transform 1 0 77556 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636993656
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636993656
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636993656
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1636993656
transform 1 0 5612 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 25201
transform 1 0 6716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 25201
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636993656
transform 1 0 7268 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1636993656
transform 1 0 8372 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1636993656
transform 1 0 9476 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1636993656
transform 1 0 10580 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 25201
transform 1 0 11684 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 25201
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1636993656
transform 1 0 12420 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1636993656
transform 1 0 13524 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1636993656
transform 1 0 14628 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1636993656
transform 1 0 15732 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 25201
transform 1 0 16836 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 25201
transform 1 0 17388 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1636993656
transform 1 0 17572 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1636993656
transform 1 0 18676 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1636993656
transform 1 0 19780 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1636993656
transform 1 0 20884 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 25201
transform 1 0 21988 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 25201
transform 1 0 22540 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1636993656
transform 1 0 22724 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1636993656
transform 1 0 23828 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1636993656
transform 1 0 24932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1636993656
transform 1 0 26036 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 25201
transform 1 0 27140 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 25201
transform 1 0 27692 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1636993656
transform 1 0 27876 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1636993656
transform 1 0 28980 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1636993656
transform 1 0 30084 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1636993656
transform 1 0 31188 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 25201
transform 1 0 32292 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 25201
transform 1 0 32844 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1636993656
transform 1 0 33028 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1636993656
transform 1 0 34132 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1636993656
transform 1 0 35236 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1636993656
transform 1 0 36340 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 25201
transform 1 0 37444 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 25201
transform 1 0 37996 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1636993656
transform 1 0 38180 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1636993656
transform 1 0 39284 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1636993656
transform 1 0 40388 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1636993656
transform 1 0 41492 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 25201
transform 1 0 42596 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 25201
transform 1 0 43148 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1636993656
transform 1 0 43332 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1636993656
transform 1 0 44436 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1636993656
transform 1 0 45540 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1636993656
transform 1 0 46644 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 25201
transform 1 0 47748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 25201
transform 1 0 48300 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1636993656
transform 1 0 48484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1636993656
transform 1 0 49588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1636993656
transform 1 0 50692 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1636993656
transform 1 0 51796 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 25201
transform 1 0 52900 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 25201
transform 1 0 53452 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1636993656
transform 1 0 53636 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1636993656
transform 1 0 54740 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1636993656
transform 1 0 55844 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1636993656
transform 1 0 56948 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 25201
transform 1 0 58052 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 25201
transform 1 0 58604 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1636993656
transform 1 0 58788 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1636993656
transform 1 0 59892 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1636993656
transform 1 0 60996 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1636993656
transform 1 0 62100 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 25201
transform 1 0 63204 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 25201
transform 1 0 63756 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1636993656
transform 1 0 63940 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1636993656
transform 1 0 65044 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_697
timestamp 1636993656
transform 1 0 66148 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_709
timestamp 1636993656
transform 1 0 67252 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 25201
transform 1 0 68356 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 25201
transform 1 0 68908 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_729
timestamp 1636993656
transform 1 0 69092 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_741
timestamp 1636993656
transform 1 0 70196 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_753
timestamp 1636993656
transform 1 0 71300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_765
timestamp 1636993656
transform 1 0 72404 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_777
timestamp 25201
transform 1 0 73508 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_783
timestamp 25201
transform 1 0 74060 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_785
timestamp 1636993656
transform 1 0 74244 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_797
timestamp 1636993656
transform 1 0 75348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_809
timestamp 1636993656
transform 1 0 76452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_821
timestamp 25201
transform 1 0 77556 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636993656
transform 1 0 2300 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636993656
transform 1 0 3404 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 25201
transform 1 0 4508 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636993656
transform 1 0 4692 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636993656
transform 1 0 5796 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636993656
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1636993656
transform 1 0 8004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 25201
transform 1 0 9108 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 25201
transform 1 0 9660 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636993656
transform 1 0 9844 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1636993656
transform 1 0 10948 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1636993656
transform 1 0 12052 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1636993656
transform 1 0 13156 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 25201
transform 1 0 14260 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 25201
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636993656
transform 1 0 14996 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1636993656
transform 1 0 16100 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1636993656
transform 1 0 17204 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1636993656
transform 1 0 18308 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 25201
transform 1 0 19412 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 25201
transform 1 0 19964 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1636993656
transform 1 0 20148 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1636993656
transform 1 0 21252 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1636993656
transform 1 0 22356 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1636993656
transform 1 0 23460 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 25201
transform 1 0 24564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 25201
transform 1 0 25116 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1636993656
transform 1 0 25300 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1636993656
transform 1 0 26404 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1636993656
transform 1 0 27508 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1636993656
transform 1 0 28612 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 25201
transform 1 0 29716 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 25201
transform 1 0 30268 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1636993656
transform 1 0 30452 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1636993656
transform 1 0 31556 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1636993656
transform 1 0 32660 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1636993656
transform 1 0 33764 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 25201
transform 1 0 34868 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 25201
transform 1 0 35420 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1636993656
transform 1 0 35604 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1636993656
transform 1 0 36708 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1636993656
transform 1 0 37812 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1636993656
transform 1 0 38916 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 25201
transform 1 0 40020 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 25201
transform 1 0 40572 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1636993656
transform 1 0 40756 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1636993656
transform 1 0 41860 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1636993656
transform 1 0 42964 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1636993656
transform 1 0 44068 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 25201
transform 1 0 45172 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 25201
transform 1 0 45724 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1636993656
transform 1 0 45908 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1636993656
transform 1 0 47012 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1636993656
transform 1 0 48116 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1636993656
transform 1 0 49220 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 25201
transform 1 0 50324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 25201
transform 1 0 50876 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1636993656
transform 1 0 51060 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1636993656
transform 1 0 52164 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1636993656
transform 1 0 53268 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1636993656
transform 1 0 54372 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 25201
transform 1 0 55476 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 25201
transform 1 0 56028 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1636993656
transform 1 0 56212 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1636993656
transform 1 0 57316 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1636993656
transform 1 0 58420 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_625
timestamp 1636993656
transform 1 0 59524 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 25201
transform 1 0 60628 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 25201
transform 1 0 61180 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1636993656
transform 1 0 61364 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1636993656
transform 1 0 62468 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1636993656
transform 1 0 63572 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_681
timestamp 1636993656
transform 1 0 64676 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 25201
transform 1 0 65780 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 25201
transform 1 0 66332 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_701
timestamp 1636993656
transform 1 0 66516 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_713
timestamp 1636993656
transform 1 0 67620 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_725
timestamp 1636993656
transform 1 0 68724 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_737
timestamp 1636993656
transform 1 0 69828 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_749
timestamp 25201
transform 1 0 70932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_755
timestamp 25201
transform 1 0 71484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_757
timestamp 1636993656
transform 1 0 71668 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_769
timestamp 1636993656
transform 1 0 72772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_781
timestamp 1636993656
transform 1 0 73876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_793
timestamp 1636993656
transform 1 0 74980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_805
timestamp 25201
transform 1 0 76084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_811
timestamp 25201
transform 1 0 76636 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_813
timestamp 25201
transform 1 0 76820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_821
timestamp 25201
transform 1 0 77556 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636993656
transform 1 0 2300 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636993656
transform 1 0 3404 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636993656
transform 1 0 4508 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636993656
transform 1 0 5612 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 25201
transform 1 0 6716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 25201
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636993656
transform 1 0 7268 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1636993656
transform 1 0 8372 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1636993656
transform 1 0 9476 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1636993656
transform 1 0 10580 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 25201
transform 1 0 11684 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 25201
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1636993656
transform 1 0 12420 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1636993656
transform 1 0 13524 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1636993656
transform 1 0 14628 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1636993656
transform 1 0 15732 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 25201
transform 1 0 16836 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 25201
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636993656
transform 1 0 17572 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1636993656
transform 1 0 18676 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1636993656
transform 1 0 19780 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1636993656
transform 1 0 20884 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 25201
transform 1 0 21988 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 25201
transform 1 0 22540 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1636993656
transform 1 0 22724 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1636993656
transform 1 0 23828 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1636993656
transform 1 0 24932 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1636993656
transform 1 0 26036 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 25201
transform 1 0 27140 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 25201
transform 1 0 27692 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1636993656
transform 1 0 27876 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1636993656
transform 1 0 28980 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1636993656
transform 1 0 30084 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1636993656
transform 1 0 31188 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 25201
transform 1 0 32292 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 25201
transform 1 0 32844 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1636993656
transform 1 0 33028 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1636993656
transform 1 0 34132 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1636993656
transform 1 0 35236 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1636993656
transform 1 0 36340 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 25201
transform 1 0 37444 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 25201
transform 1 0 37996 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1636993656
transform 1 0 38180 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1636993656
transform 1 0 39284 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1636993656
transform 1 0 40388 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1636993656
transform 1 0 41492 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 25201
transform 1 0 42596 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 25201
transform 1 0 43148 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1636993656
transform 1 0 43332 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1636993656
transform 1 0 44436 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1636993656
transform 1 0 45540 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1636993656
transform 1 0 46644 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 25201
transform 1 0 47748 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 25201
transform 1 0 48300 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1636993656
transform 1 0 48484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1636993656
transform 1 0 49588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1636993656
transform 1 0 50692 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1636993656
transform 1 0 51796 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 25201
transform 1 0 52900 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 25201
transform 1 0 53452 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1636993656
transform 1 0 53636 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1636993656
transform 1 0 54740 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1636993656
transform 1 0 55844 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1636993656
transform 1 0 56948 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 25201
transform 1 0 58052 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 25201
transform 1 0 58604 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1636993656
transform 1 0 58788 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1636993656
transform 1 0 59892 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1636993656
transform 1 0 60996 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1636993656
transform 1 0 62100 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 25201
transform 1 0 63204 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 25201
transform 1 0 63756 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_673
timestamp 1636993656
transform 1 0 63940 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_685
timestamp 1636993656
transform 1 0 65044 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_697
timestamp 1636993656
transform 1 0 66148 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_709
timestamp 1636993656
transform 1 0 67252 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 25201
transform 1 0 68356 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 25201
transform 1 0 68908 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_729
timestamp 1636993656
transform 1 0 69092 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_741
timestamp 1636993656
transform 1 0 70196 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_753
timestamp 1636993656
transform 1 0 71300 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_765
timestamp 1636993656
transform 1 0 72404 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_777
timestamp 25201
transform 1 0 73508 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_783
timestamp 25201
transform 1 0 74060 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_785
timestamp 1636993656
transform 1 0 74244 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_797
timestamp 1636993656
transform 1 0 75348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_809
timestamp 1636993656
transform 1 0 76452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_821
timestamp 25201
transform 1 0 77556 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636993656
transform 1 0 2300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636993656
transform 1 0 3404 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 25201
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636993656
transform 1 0 4692 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636993656
transform 1 0 5796 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636993656
transform 1 0 6900 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1636993656
transform 1 0 8004 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 25201
transform 1 0 9108 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 25201
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1636993656
transform 1 0 9844 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1636993656
transform 1 0 10948 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1636993656
transform 1 0 12052 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1636993656
transform 1 0 13156 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 25201
transform 1 0 14260 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 25201
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1636993656
transform 1 0 14996 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1636993656
transform 1 0 16100 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1636993656
transform 1 0 17204 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1636993656
transform 1 0 18308 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 25201
transform 1 0 19412 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 25201
transform 1 0 19964 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1636993656
transform 1 0 20148 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1636993656
transform 1 0 21252 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1636993656
transform 1 0 22356 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1636993656
transform 1 0 23460 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 25201
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 25201
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1636993656
transform 1 0 25300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1636993656
transform 1 0 26404 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1636993656
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1636993656
transform 1 0 28612 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 25201
transform 1 0 29716 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 25201
transform 1 0 30268 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1636993656
transform 1 0 30452 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1636993656
transform 1 0 31556 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1636993656
transform 1 0 32660 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1636993656
transform 1 0 33764 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 25201
transform 1 0 34868 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 25201
transform 1 0 35420 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1636993656
transform 1 0 35604 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1636993656
transform 1 0 36708 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1636993656
transform 1 0 37812 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1636993656
transform 1 0 38916 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 25201
transform 1 0 40020 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 25201
transform 1 0 40572 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1636993656
transform 1 0 40756 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1636993656
transform 1 0 41860 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1636993656
transform 1 0 42964 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1636993656
transform 1 0 44068 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 25201
transform 1 0 45172 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 25201
transform 1 0 45724 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1636993656
transform 1 0 45908 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1636993656
transform 1 0 47012 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1636993656
transform 1 0 48116 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1636993656
transform 1 0 49220 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 25201
transform 1 0 50324 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 25201
transform 1 0 50876 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1636993656
transform 1 0 51060 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1636993656
transform 1 0 52164 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1636993656
transform 1 0 53268 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1636993656
transform 1 0 54372 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 25201
transform 1 0 55476 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 25201
transform 1 0 56028 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1636993656
transform 1 0 56212 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1636993656
transform 1 0 57316 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1636993656
transform 1 0 58420 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1636993656
transform 1 0 59524 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 25201
transform 1 0 60628 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 25201
transform 1 0 61180 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1636993656
transform 1 0 61364 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1636993656
transform 1 0 62468 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1636993656
transform 1 0 63572 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_681
timestamp 1636993656
transform 1 0 64676 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 25201
transform 1 0 65780 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 25201
transform 1 0 66332 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_701
timestamp 1636993656
transform 1 0 66516 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_713
timestamp 1636993656
transform 1 0 67620 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_725
timestamp 1636993656
transform 1 0 68724 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_737
timestamp 1636993656
transform 1 0 69828 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_749
timestamp 25201
transform 1 0 70932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_755
timestamp 25201
transform 1 0 71484 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_757
timestamp 1636993656
transform 1 0 71668 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_769
timestamp 1636993656
transform 1 0 72772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_781
timestamp 1636993656
transform 1 0 73876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_793
timestamp 1636993656
transform 1 0 74980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_805
timestamp 25201
transform 1 0 76084 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_811
timestamp 25201
transform 1 0 76636 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_813
timestamp 25201
transform 1 0 76820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_821
timestamp 25201
transform 1 0 77556 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636993656
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636993656
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1636993656
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1636993656
transform 1 0 5612 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 25201
transform 1 0 6716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 25201
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636993656
transform 1 0 7268 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1636993656
transform 1 0 8372 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1636993656
transform 1 0 9476 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1636993656
transform 1 0 10580 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 25201
transform 1 0 11684 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 25201
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1636993656
transform 1 0 12420 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1636993656
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1636993656
transform 1 0 14628 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1636993656
transform 1 0 15732 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 25201
transform 1 0 16836 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 25201
transform 1 0 17388 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1636993656
transform 1 0 17572 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1636993656
transform 1 0 18676 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1636993656
transform 1 0 19780 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1636993656
transform 1 0 20884 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 25201
transform 1 0 21988 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 25201
transform 1 0 22540 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636993656
transform 1 0 22724 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1636993656
transform 1 0 23828 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1636993656
transform 1 0 24932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1636993656
transform 1 0 26036 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 25201
transform 1 0 27140 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 25201
transform 1 0 27692 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1636993656
transform 1 0 27876 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1636993656
transform 1 0 28980 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1636993656
transform 1 0 30084 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1636993656
transform 1 0 31188 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 25201
transform 1 0 32292 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 25201
transform 1 0 32844 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1636993656
transform 1 0 33028 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1636993656
transform 1 0 34132 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1636993656
transform 1 0 35236 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1636993656
transform 1 0 36340 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 25201
transform 1 0 37444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 25201
transform 1 0 37996 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1636993656
transform 1 0 38180 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1636993656
transform 1 0 39284 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1636993656
transform 1 0 40388 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1636993656
transform 1 0 41492 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 25201
transform 1 0 42596 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 25201
transform 1 0 43148 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1636993656
transform 1 0 43332 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1636993656
transform 1 0 44436 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1636993656
transform 1 0 45540 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1636993656
transform 1 0 46644 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 25201
transform 1 0 47748 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 25201
transform 1 0 48300 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1636993656
transform 1 0 48484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1636993656
transform 1 0 49588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1636993656
transform 1 0 50692 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1636993656
transform 1 0 51796 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 25201
transform 1 0 52900 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 25201
transform 1 0 53452 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1636993656
transform 1 0 53636 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1636993656
transform 1 0 54740 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1636993656
transform 1 0 55844 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1636993656
transform 1 0 56948 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 25201
transform 1 0 58052 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 25201
transform 1 0 58604 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1636993656
transform 1 0 58788 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1636993656
transform 1 0 59892 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1636993656
transform 1 0 60996 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1636993656
transform 1 0 62100 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 25201
transform 1 0 63204 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 25201
transform 1 0 63756 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1636993656
transform 1 0 63940 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1636993656
transform 1 0 65044 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1636993656
transform 1 0 66148 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_709
timestamp 1636993656
transform 1 0 67252 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 25201
transform 1 0 68356 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 25201
transform 1 0 68908 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_729
timestamp 1636993656
transform 1 0 69092 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_741
timestamp 1636993656
transform 1 0 70196 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_753
timestamp 1636993656
transform 1 0 71300 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_765
timestamp 1636993656
transform 1 0 72404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_777
timestamp 25201
transform 1 0 73508 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_783
timestamp 25201
transform 1 0 74060 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_785
timestamp 1636993656
transform 1 0 74244 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_797
timestamp 1636993656
transform 1 0 75348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_809
timestamp 1636993656
transform 1 0 76452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_821
timestamp 25201
transform 1 0 77556 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636993656
transform 1 0 2300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636993656
transform 1 0 3404 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 25201
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636993656
transform 1 0 4692 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636993656
transform 1 0 5796 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636993656
transform 1 0 6900 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1636993656
transform 1 0 8004 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 25201
transform 1 0 9108 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 25201
transform 1 0 9660 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636993656
transform 1 0 9844 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1636993656
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1636993656
transform 1 0 12052 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1636993656
transform 1 0 13156 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 25201
transform 1 0 14260 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 25201
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636993656
transform 1 0 14996 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1636993656
transform 1 0 16100 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1636993656
transform 1 0 17204 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1636993656
transform 1 0 18308 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 25201
transform 1 0 19412 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 25201
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636993656
transform 1 0 20148 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1636993656
transform 1 0 21252 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1636993656
transform 1 0 22356 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1636993656
transform 1 0 23460 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 25201
transform 1 0 24564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 25201
transform 1 0 25116 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1636993656
transform 1 0 25300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1636993656
transform 1 0 26404 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1636993656
transform 1 0 27508 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1636993656
transform 1 0 28612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 25201
transform 1 0 29716 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 25201
transform 1 0 30268 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1636993656
transform 1 0 30452 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1636993656
transform 1 0 31556 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1636993656
transform 1 0 32660 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1636993656
transform 1 0 33764 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 25201
transform 1 0 34868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 25201
transform 1 0 35420 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1636993656
transform 1 0 35604 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1636993656
transform 1 0 36708 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1636993656
transform 1 0 37812 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1636993656
transform 1 0 38916 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 25201
transform 1 0 40020 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 25201
transform 1 0 40572 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1636993656
transform 1 0 40756 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1636993656
transform 1 0 41860 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1636993656
transform 1 0 42964 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1636993656
transform 1 0 44068 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 25201
transform 1 0 45172 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 25201
transform 1 0 45724 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1636993656
transform 1 0 45908 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1636993656
transform 1 0 47012 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1636993656
transform 1 0 48116 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1636993656
transform 1 0 49220 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 25201
transform 1 0 50324 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 25201
transform 1 0 50876 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1636993656
transform 1 0 51060 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1636993656
transform 1 0 52164 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1636993656
transform 1 0 53268 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1636993656
transform 1 0 54372 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 25201
transform 1 0 55476 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 25201
transform 1 0 56028 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1636993656
transform 1 0 56212 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1636993656
transform 1 0 57316 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1636993656
transform 1 0 58420 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1636993656
transform 1 0 59524 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 25201
transform 1 0 60628 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 25201
transform 1 0 61180 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1636993656
transform 1 0 61364 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1636993656
transform 1 0 62468 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1636993656
transform 1 0 63572 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1636993656
transform 1 0 64676 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 25201
transform 1 0 65780 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 25201
transform 1 0 66332 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1636993656
transform 1 0 66516 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_713
timestamp 1636993656
transform 1 0 67620 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_725
timestamp 1636993656
transform 1 0 68724 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_737
timestamp 1636993656
transform 1 0 69828 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_749
timestamp 25201
transform 1 0 70932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_755
timestamp 25201
transform 1 0 71484 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_757
timestamp 1636993656
transform 1 0 71668 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_769
timestamp 1636993656
transform 1 0 72772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_781
timestamp 1636993656
transform 1 0 73876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_793
timestamp 1636993656
transform 1 0 74980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_805
timestamp 25201
transform 1 0 76084 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_811
timestamp 25201
transform 1 0 76636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_813
timestamp 25201
transform 1 0 76820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_821
timestamp 25201
transform 1 0 77556 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636993656
transform 1 0 2300 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636993656
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636993656
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636993656
transform 1 0 5612 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 25201
transform 1 0 6716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 25201
transform 1 0 7084 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636993656
transform 1 0 7268 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1636993656
transform 1 0 8372 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1636993656
transform 1 0 9476 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1636993656
transform 1 0 10580 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 25201
transform 1 0 11684 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 25201
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1636993656
transform 1 0 12420 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1636993656
transform 1 0 13524 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1636993656
transform 1 0 14628 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1636993656
transform 1 0 15732 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 25201
transform 1 0 16836 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 25201
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1636993656
transform 1 0 17572 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1636993656
transform 1 0 18676 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1636993656
transform 1 0 19780 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1636993656
transform 1 0 20884 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 25201
transform 1 0 21988 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 25201
transform 1 0 22540 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1636993656
transform 1 0 22724 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1636993656
transform 1 0 23828 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1636993656
transform 1 0 24932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1636993656
transform 1 0 26036 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 25201
transform 1 0 27140 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 25201
transform 1 0 27692 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1636993656
transform 1 0 27876 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1636993656
transform 1 0 28980 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1636993656
transform 1 0 30084 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1636993656
transform 1 0 31188 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 25201
transform 1 0 32292 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 25201
transform 1 0 32844 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1636993656
transform 1 0 33028 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1636993656
transform 1 0 34132 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1636993656
transform 1 0 35236 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1636993656
transform 1 0 36340 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 25201
transform 1 0 37444 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 25201
transform 1 0 37996 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1636993656
transform 1 0 38180 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1636993656
transform 1 0 39284 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1636993656
transform 1 0 40388 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1636993656
transform 1 0 41492 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 25201
transform 1 0 42596 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 25201
transform 1 0 43148 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1636993656
transform 1 0 43332 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1636993656
transform 1 0 44436 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1636993656
transform 1 0 45540 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1636993656
transform 1 0 46644 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 25201
transform 1 0 47748 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 25201
transform 1 0 48300 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1636993656
transform 1 0 48484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1636993656
transform 1 0 49588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1636993656
transform 1 0 50692 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1636993656
transform 1 0 51796 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 25201
transform 1 0 52900 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 25201
transform 1 0 53452 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1636993656
transform 1 0 53636 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1636993656
transform 1 0 54740 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1636993656
transform 1 0 55844 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1636993656
transform 1 0 56948 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 25201
transform 1 0 58052 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 25201
transform 1 0 58604 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1636993656
transform 1 0 58788 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1636993656
transform 1 0 59892 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1636993656
transform 1 0 60996 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1636993656
transform 1 0 62100 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 25201
transform 1 0 63204 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 25201
transform 1 0 63756 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_673
timestamp 1636993656
transform 1 0 63940 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_685
timestamp 1636993656
transform 1 0 65044 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1636993656
transform 1 0 66148 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_709
timestamp 1636993656
transform 1 0 67252 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 25201
transform 1 0 68356 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 25201
transform 1 0 68908 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_729
timestamp 1636993656
transform 1 0 69092 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_741
timestamp 1636993656
transform 1 0 70196 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_753
timestamp 1636993656
transform 1 0 71300 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_765
timestamp 1636993656
transform 1 0 72404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_777
timestamp 25201
transform 1 0 73508 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_783
timestamp 25201
transform 1 0 74060 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_785
timestamp 1636993656
transform 1 0 74244 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_797
timestamp 1636993656
transform 1 0 75348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_809
timestamp 1636993656
transform 1 0 76452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_821
timestamp 25201
transform 1 0 77556 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636993656
transform 1 0 2300 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636993656
transform 1 0 3404 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 25201
transform 1 0 4508 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636993656
transform 1 0 4692 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636993656
transform 1 0 5796 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636993656
transform 1 0 6900 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1636993656
transform 1 0 8004 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 25201
transform 1 0 9108 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 25201
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1636993656
transform 1 0 9844 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1636993656
transform 1 0 10948 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1636993656
transform 1 0 12052 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1636993656
transform 1 0 13156 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 25201
transform 1 0 14260 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 25201
transform 1 0 14812 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1636993656
transform 1 0 14996 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1636993656
transform 1 0 16100 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1636993656
transform 1 0 17204 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1636993656
transform 1 0 18308 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 25201
transform 1 0 19412 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 25201
transform 1 0 19964 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1636993656
transform 1 0 20148 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1636993656
transform 1 0 21252 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1636993656
transform 1 0 22356 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1636993656
transform 1 0 23460 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 25201
transform 1 0 24564 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 25201
transform 1 0 25116 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1636993656
transform 1 0 25300 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1636993656
transform 1 0 26404 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1636993656
transform 1 0 27508 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1636993656
transform 1 0 28612 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 25201
transform 1 0 29716 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 25201
transform 1 0 30268 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1636993656
transform 1 0 30452 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1636993656
transform 1 0 31556 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1636993656
transform 1 0 32660 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1636993656
transform 1 0 33764 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 25201
transform 1 0 34868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 25201
transform 1 0 35420 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1636993656
transform 1 0 35604 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1636993656
transform 1 0 36708 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1636993656
transform 1 0 37812 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1636993656
transform 1 0 38916 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 25201
transform 1 0 40020 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 25201
transform 1 0 40572 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1636993656
transform 1 0 40756 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1636993656
transform 1 0 41860 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1636993656
transform 1 0 42964 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1636993656
transform 1 0 44068 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 25201
transform 1 0 45172 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 25201
transform 1 0 45724 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1636993656
transform 1 0 45908 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1636993656
transform 1 0 47012 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1636993656
transform 1 0 48116 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1636993656
transform 1 0 49220 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 25201
transform 1 0 50324 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 25201
transform 1 0 50876 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1636993656
transform 1 0 51060 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1636993656
transform 1 0 52164 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1636993656
transform 1 0 53268 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1636993656
transform 1 0 54372 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 25201
transform 1 0 55476 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 25201
transform 1 0 56028 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1636993656
transform 1 0 56212 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1636993656
transform 1 0 57316 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1636993656
transform 1 0 58420 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_625
timestamp 1636993656
transform 1 0 59524 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 25201
transform 1 0 60628 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 25201
transform 1 0 61180 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1636993656
transform 1 0 61364 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1636993656
transform 1 0 62468 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_669
timestamp 1636993656
transform 1 0 63572 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_681
timestamp 1636993656
transform 1 0 64676 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 25201
transform 1 0 65780 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 25201
transform 1 0 66332 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1636993656
transform 1 0 66516 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1636993656
transform 1 0 67620 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_725
timestamp 1636993656
transform 1 0 68724 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_737
timestamp 1636993656
transform 1 0 69828 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_749
timestamp 25201
transform 1 0 70932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_755
timestamp 25201
transform 1 0 71484 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_757
timestamp 1636993656
transform 1 0 71668 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_769
timestamp 1636993656
transform 1 0 72772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_781
timestamp 1636993656
transform 1 0 73876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_793
timestamp 1636993656
transform 1 0 74980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_805
timestamp 25201
transform 1 0 76084 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_811
timestamp 25201
transform 1 0 76636 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_813
timestamp 25201
transform 1 0 76820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_821
timestamp 25201
transform 1 0 77556 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636993656
transform 1 0 2300 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636993656
transform 1 0 3404 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636993656
transform 1 0 4508 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636993656
transform 1 0 5612 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 25201
transform 1 0 6716 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 25201
transform 1 0 7084 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636993656
transform 1 0 7268 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1636993656
transform 1 0 8372 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1636993656
transform 1 0 9476 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1636993656
transform 1 0 10580 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 25201
transform 1 0 11684 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 25201
transform 1 0 12236 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1636993656
transform 1 0 12420 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1636993656
transform 1 0 13524 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1636993656
transform 1 0 14628 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1636993656
transform 1 0 15732 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 25201
transform 1 0 16836 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 25201
transform 1 0 17388 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1636993656
transform 1 0 17572 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1636993656
transform 1 0 18676 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1636993656
transform 1 0 19780 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1636993656
transform 1 0 20884 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 25201
transform 1 0 21988 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 25201
transform 1 0 22540 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1636993656
transform 1 0 22724 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1636993656
transform 1 0 23828 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1636993656
transform 1 0 24932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1636993656
transform 1 0 26036 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 25201
transform 1 0 27140 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 25201
transform 1 0 27692 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1636993656
transform 1 0 27876 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1636993656
transform 1 0 28980 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1636993656
transform 1 0 30084 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1636993656
transform 1 0 31188 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 25201
transform 1 0 32292 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 25201
transform 1 0 32844 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1636993656
transform 1 0 33028 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1636993656
transform 1 0 34132 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1636993656
transform 1 0 35236 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1636993656
transform 1 0 36340 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 25201
transform 1 0 37444 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 25201
transform 1 0 37996 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1636993656
transform 1 0 38180 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1636993656
transform 1 0 39284 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1636993656
transform 1 0 40388 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1636993656
transform 1 0 41492 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 25201
transform 1 0 42596 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 25201
transform 1 0 43148 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1636993656
transform 1 0 43332 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1636993656
transform 1 0 44436 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1636993656
transform 1 0 45540 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1636993656
transform 1 0 46644 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 25201
transform 1 0 47748 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 25201
transform 1 0 48300 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1636993656
transform 1 0 48484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1636993656
transform 1 0 49588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1636993656
transform 1 0 50692 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1636993656
transform 1 0 51796 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 25201
transform 1 0 52900 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 25201
transform 1 0 53452 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1636993656
transform 1 0 53636 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1636993656
transform 1 0 54740 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1636993656
transform 1 0 55844 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1636993656
transform 1 0 56948 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 25201
transform 1 0 58052 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 25201
transform 1 0 58604 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1636993656
transform 1 0 58788 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1636993656
transform 1 0 59892 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1636993656
transform 1 0 60996 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1636993656
transform 1 0 62100 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 25201
transform 1 0 63204 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 25201
transform 1 0 63756 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1636993656
transform 1 0 63940 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1636993656
transform 1 0 65044 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1636993656
transform 1 0 66148 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1636993656
transform 1 0 67252 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 25201
transform 1 0 68356 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 25201
transform 1 0 68908 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_729
timestamp 1636993656
transform 1 0 69092 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_741
timestamp 1636993656
transform 1 0 70196 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_753
timestamp 1636993656
transform 1 0 71300 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_765
timestamp 1636993656
transform 1 0 72404 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_777
timestamp 25201
transform 1 0 73508 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_783
timestamp 25201
transform 1 0 74060 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_785
timestamp 1636993656
transform 1 0 74244 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_797
timestamp 1636993656
transform 1 0 75348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_809
timestamp 1636993656
transform 1 0 76452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_821
timestamp 25201
transform 1 0 77556 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636993656
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636993656
transform 1 0 3404 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 25201
transform 1 0 4508 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636993656
transform 1 0 4692 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636993656
transform 1 0 5796 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636993656
transform 1 0 6900 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1636993656
transform 1 0 8004 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 25201
transform 1 0 9108 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 25201
transform 1 0 9660 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1636993656
transform 1 0 9844 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1636993656
transform 1 0 10948 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1636993656
transform 1 0 12052 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1636993656
transform 1 0 13156 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 25201
transform 1 0 14260 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 25201
transform 1 0 14812 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1636993656
transform 1 0 14996 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1636993656
transform 1 0 16100 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1636993656
transform 1 0 17204 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1636993656
transform 1 0 18308 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 25201
transform 1 0 19412 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 25201
transform 1 0 19964 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1636993656
transform 1 0 20148 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1636993656
transform 1 0 21252 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1636993656
transform 1 0 22356 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1636993656
transform 1 0 23460 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 25201
transform 1 0 24564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 25201
transform 1 0 25116 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1636993656
transform 1 0 25300 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1636993656
transform 1 0 26404 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1636993656
transform 1 0 27508 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1636993656
transform 1 0 28612 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 25201
transform 1 0 29716 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 25201
transform 1 0 30268 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1636993656
transform 1 0 30452 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1636993656
transform 1 0 31556 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1636993656
transform 1 0 32660 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1636993656
transform 1 0 33764 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 25201
transform 1 0 34868 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 25201
transform 1 0 35420 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1636993656
transform 1 0 35604 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1636993656
transform 1 0 36708 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1636993656
transform 1 0 37812 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1636993656
transform 1 0 38916 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 25201
transform 1 0 40020 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 25201
transform 1 0 40572 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1636993656
transform 1 0 40756 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1636993656
transform 1 0 41860 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1636993656
transform 1 0 42964 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1636993656
transform 1 0 44068 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 25201
transform 1 0 45172 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 25201
transform 1 0 45724 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1636993656
transform 1 0 45908 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1636993656
transform 1 0 47012 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1636993656
transform 1 0 48116 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1636993656
transform 1 0 49220 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 25201
transform 1 0 50324 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 25201
transform 1 0 50876 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1636993656
transform 1 0 51060 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1636993656
transform 1 0 52164 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1636993656
transform 1 0 53268 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1636993656
transform 1 0 54372 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 25201
transform 1 0 55476 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 25201
transform 1 0 56028 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1636993656
transform 1 0 56212 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1636993656
transform 1 0 57316 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1636993656
transform 1 0 58420 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1636993656
transform 1 0 59524 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 25201
transform 1 0 60628 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 25201
transform 1 0 61180 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1636993656
transform 1 0 61364 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1636993656
transform 1 0 62468 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1636993656
transform 1 0 63572 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1636993656
transform 1 0 64676 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 25201
transform 1 0 65780 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 25201
transform 1 0 66332 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1636993656
transform 1 0 66516 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1636993656
transform 1 0 67620 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_725
timestamp 1636993656
transform 1 0 68724 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_737
timestamp 1636993656
transform 1 0 69828 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_749
timestamp 25201
transform 1 0 70932 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_755
timestamp 25201
transform 1 0 71484 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_757
timestamp 1636993656
transform 1 0 71668 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_769
timestamp 1636993656
transform 1 0 72772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_781
timestamp 1636993656
transform 1 0 73876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_793
timestamp 1636993656
transform 1 0 74980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_805
timestamp 25201
transform 1 0 76084 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_811
timestamp 25201
transform 1 0 76636 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_813
timestamp 25201
transform 1 0 76820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_821
timestamp 25201
transform 1 0 77556 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636993656
transform 1 0 2300 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636993656
transform 1 0 3404 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636993656
transform 1 0 4508 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1636993656
transform 1 0 5612 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 25201
transform 1 0 6716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 25201
transform 1 0 7084 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636993656
transform 1 0 7268 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1636993656
transform 1 0 8372 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1636993656
transform 1 0 9476 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1636993656
transform 1 0 10580 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 25201
transform 1 0 11684 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 25201
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1636993656
transform 1 0 12420 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1636993656
transform 1 0 13524 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1636993656
transform 1 0 14628 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1636993656
transform 1 0 15732 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 25201
transform 1 0 16836 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 25201
transform 1 0 17388 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1636993656
transform 1 0 17572 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1636993656
transform 1 0 18676 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1636993656
transform 1 0 19780 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1636993656
transform 1 0 20884 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 25201
transform 1 0 21988 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 25201
transform 1 0 22540 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1636993656
transform 1 0 22724 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1636993656
transform 1 0 23828 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1636993656
transform 1 0 24932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1636993656
transform 1 0 26036 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 25201
transform 1 0 27140 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 25201
transform 1 0 27692 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1636993656
transform 1 0 27876 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1636993656
transform 1 0 28980 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1636993656
transform 1 0 30084 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1636993656
transform 1 0 31188 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 25201
transform 1 0 32292 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 25201
transform 1 0 32844 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1636993656
transform 1 0 33028 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1636993656
transform 1 0 34132 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1636993656
transform 1 0 35236 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1636993656
transform 1 0 36340 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 25201
transform 1 0 37444 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 25201
transform 1 0 37996 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1636993656
transform 1 0 38180 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1636993656
transform 1 0 39284 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1636993656
transform 1 0 40388 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1636993656
transform 1 0 41492 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 25201
transform 1 0 42596 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 25201
transform 1 0 43148 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1636993656
transform 1 0 43332 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1636993656
transform 1 0 44436 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1636993656
transform 1 0 45540 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1636993656
transform 1 0 46644 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 25201
transform 1 0 47748 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 25201
transform 1 0 48300 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1636993656
transform 1 0 48484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1636993656
transform 1 0 49588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1636993656
transform 1 0 50692 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1636993656
transform 1 0 51796 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 25201
transform 1 0 52900 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 25201
transform 1 0 53452 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1636993656
transform 1 0 53636 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1636993656
transform 1 0 54740 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1636993656
transform 1 0 55844 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1636993656
transform 1 0 56948 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 25201
transform 1 0 58052 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 25201
transform 1 0 58604 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1636993656
transform 1 0 58788 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1636993656
transform 1 0 59892 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1636993656
transform 1 0 60996 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1636993656
transform 1 0 62100 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 25201
transform 1 0 63204 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 25201
transform 1 0 63756 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1636993656
transform 1 0 63940 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1636993656
transform 1 0 65044 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1636993656
transform 1 0 66148 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1636993656
transform 1 0 67252 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 25201
transform 1 0 68356 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 25201
transform 1 0 68908 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_729
timestamp 1636993656
transform 1 0 69092 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_741
timestamp 1636993656
transform 1 0 70196 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_753
timestamp 1636993656
transform 1 0 71300 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_765
timestamp 1636993656
transform 1 0 72404 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_777
timestamp 25201
transform 1 0 73508 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_783
timestamp 25201
transform 1 0 74060 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_785
timestamp 1636993656
transform 1 0 74244 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_797
timestamp 1636993656
transform 1 0 75348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_809
timestamp 1636993656
transform 1 0 76452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_821
timestamp 25201
transform 1 0 77556 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636993656
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636993656
transform 1 0 3404 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 25201
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636993656
transform 1 0 4692 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636993656
transform 1 0 5796 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636993656
transform 1 0 6900 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1636993656
transform 1 0 8004 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 25201
transform 1 0 9108 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 25201
transform 1 0 9660 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1636993656
transform 1 0 9844 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1636993656
transform 1 0 10948 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1636993656
transform 1 0 12052 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1636993656
transform 1 0 13156 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 25201
transform 1 0 14260 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 25201
transform 1 0 14812 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1636993656
transform 1 0 14996 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1636993656
transform 1 0 16100 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1636993656
transform 1 0 17204 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1636993656
transform 1 0 18308 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 25201
transform 1 0 19412 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 25201
transform 1 0 19964 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1636993656
transform 1 0 20148 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1636993656
transform 1 0 21252 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1636993656
transform 1 0 22356 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1636993656
transform 1 0 23460 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 25201
transform 1 0 24564 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 25201
transform 1 0 25116 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1636993656
transform 1 0 25300 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1636993656
transform 1 0 26404 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1636993656
transform 1 0 27508 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1636993656
transform 1 0 28612 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 25201
transform 1 0 29716 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 25201
transform 1 0 30268 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1636993656
transform 1 0 30452 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1636993656
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1636993656
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1636993656
transform 1 0 33764 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 25201
transform 1 0 34868 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 25201
transform 1 0 35420 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1636993656
transform 1 0 35604 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1636993656
transform 1 0 36708 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1636993656
transform 1 0 37812 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1636993656
transform 1 0 38916 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 25201
transform 1 0 40020 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 25201
transform 1 0 40572 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1636993656
transform 1 0 40756 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1636993656
transform 1 0 41860 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1636993656
transform 1 0 42964 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1636993656
transform 1 0 44068 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 25201
transform 1 0 45172 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 25201
transform 1 0 45724 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1636993656
transform 1 0 45908 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1636993656
transform 1 0 47012 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1636993656
transform 1 0 48116 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1636993656
transform 1 0 49220 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 25201
transform 1 0 50324 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 25201
transform 1 0 50876 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1636993656
transform 1 0 51060 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1636993656
transform 1 0 52164 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1636993656
transform 1 0 53268 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1636993656
transform 1 0 54372 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 25201
transform 1 0 55476 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 25201
transform 1 0 56028 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1636993656
transform 1 0 56212 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1636993656
transform 1 0 57316 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1636993656
transform 1 0 58420 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1636993656
transform 1 0 59524 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 25201
transform 1 0 60628 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 25201
transform 1 0 61180 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1636993656
transform 1 0 61364 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1636993656
transform 1 0 62468 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1636993656
transform 1 0 63572 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1636993656
transform 1 0 64676 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 25201
transform 1 0 65780 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 25201
transform 1 0 66332 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1636993656
transform 1 0 66516 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1636993656
transform 1 0 67620 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_725
timestamp 1636993656
transform 1 0 68724 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_737
timestamp 1636993656
transform 1 0 69828 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_749
timestamp 25201
transform 1 0 70932 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_755
timestamp 25201
transform 1 0 71484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_757
timestamp 1636993656
transform 1 0 71668 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_769
timestamp 1636993656
transform 1 0 72772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_781
timestamp 1636993656
transform 1 0 73876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_793
timestamp 1636993656
transform 1 0 74980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_805
timestamp 25201
transform 1 0 76084 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_811
timestamp 25201
transform 1 0 76636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_813
timestamp 25201
transform 1 0 76820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_821
timestamp 25201
transform 1 0 77556 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636993656
transform 1 0 2300 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636993656
transform 1 0 3404 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636993656
transform 1 0 4508 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1636993656
transform 1 0 5612 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 25201
transform 1 0 6716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 25201
transform 1 0 7084 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636993656
transform 1 0 7268 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1636993656
transform 1 0 8372 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1636993656
transform 1 0 9476 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1636993656
transform 1 0 10580 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 25201
transform 1 0 11684 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 25201
transform 1 0 12236 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1636993656
transform 1 0 12420 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1636993656
transform 1 0 13524 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1636993656
transform 1 0 14628 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1636993656
transform 1 0 15732 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 25201
transform 1 0 16836 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 25201
transform 1 0 17388 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1636993656
transform 1 0 17572 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1636993656
transform 1 0 18676 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1636993656
transform 1 0 19780 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1636993656
transform 1 0 20884 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 25201
transform 1 0 21988 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 25201
transform 1 0 22540 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1636993656
transform 1 0 22724 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1636993656
transform 1 0 23828 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1636993656
transform 1 0 24932 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1636993656
transform 1 0 26036 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 25201
transform 1 0 27140 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 25201
transform 1 0 27692 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1636993656
transform 1 0 27876 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1636993656
transform 1 0 28980 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1636993656
transform 1 0 30084 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1636993656
transform 1 0 31188 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 25201
transform 1 0 32292 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 25201
transform 1 0 32844 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1636993656
transform 1 0 33028 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1636993656
transform 1 0 34132 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1636993656
transform 1 0 35236 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1636993656
transform 1 0 36340 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 25201
transform 1 0 37444 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 25201
transform 1 0 37996 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1636993656
transform 1 0 38180 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1636993656
transform 1 0 39284 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1636993656
transform 1 0 40388 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1636993656
transform 1 0 41492 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 25201
transform 1 0 42596 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 25201
transform 1 0 43148 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1636993656
transform 1 0 43332 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1636993656
transform 1 0 44436 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1636993656
transform 1 0 45540 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1636993656
transform 1 0 46644 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 25201
transform 1 0 47748 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 25201
transform 1 0 48300 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1636993656
transform 1 0 48484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1636993656
transform 1 0 49588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1636993656
transform 1 0 50692 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1636993656
transform 1 0 51796 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 25201
transform 1 0 52900 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 25201
transform 1 0 53452 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1636993656
transform 1 0 53636 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1636993656
transform 1 0 54740 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1636993656
transform 1 0 55844 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1636993656
transform 1 0 56948 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 25201
transform 1 0 58052 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 25201
transform 1 0 58604 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1636993656
transform 1 0 58788 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1636993656
transform 1 0 59892 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1636993656
transform 1 0 60996 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1636993656
transform 1 0 62100 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 25201
transform 1 0 63204 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 25201
transform 1 0 63756 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1636993656
transform 1 0 63940 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1636993656
transform 1 0 65044 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1636993656
transform 1 0 66148 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1636993656
transform 1 0 67252 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 25201
transform 1 0 68356 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 25201
transform 1 0 68908 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_729
timestamp 1636993656
transform 1 0 69092 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_741
timestamp 1636993656
transform 1 0 70196 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_753
timestamp 1636993656
transform 1 0 71300 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_765
timestamp 1636993656
transform 1 0 72404 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_777
timestamp 25201
transform 1 0 73508 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_783
timestamp 25201
transform 1 0 74060 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_785
timestamp 1636993656
transform 1 0 74244 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_797
timestamp 1636993656
transform 1 0 75348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_809
timestamp 1636993656
transform 1 0 76452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_821
timestamp 25201
transform 1 0 77556 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636993656
transform 1 0 2300 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636993656
transform 1 0 3404 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 25201
transform 1 0 4508 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636993656
transform 1 0 4692 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1636993656
transform 1 0 5796 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1636993656
transform 1 0 6900 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1636993656
transform 1 0 8004 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 25201
transform 1 0 9108 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 25201
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1636993656
transform 1 0 9844 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1636993656
transform 1 0 10948 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1636993656
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1636993656
transform 1 0 13156 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 25201
transform 1 0 14260 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 25201
transform 1 0 14812 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1636993656
transform 1 0 14996 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1636993656
transform 1 0 16100 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1636993656
transform 1 0 17204 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1636993656
transform 1 0 18308 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 25201
transform 1 0 19412 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 25201
transform 1 0 19964 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1636993656
transform 1 0 20148 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1636993656
transform 1 0 21252 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1636993656
transform 1 0 22356 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1636993656
transform 1 0 23460 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 25201
transform 1 0 24564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 25201
transform 1 0 25116 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1636993656
transform 1 0 25300 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1636993656
transform 1 0 26404 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1636993656
transform 1 0 27508 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1636993656
transform 1 0 28612 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 25201
transform 1 0 29716 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 25201
transform 1 0 30268 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1636993656
transform 1 0 30452 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1636993656
transform 1 0 31556 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1636993656
transform 1 0 32660 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1636993656
transform 1 0 33764 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 25201
transform 1 0 34868 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 25201
transform 1 0 35420 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1636993656
transform 1 0 35604 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1636993656
transform 1 0 36708 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1636993656
transform 1 0 37812 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1636993656
transform 1 0 38916 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 25201
transform 1 0 40020 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 25201
transform 1 0 40572 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1636993656
transform 1 0 40756 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1636993656
transform 1 0 41860 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1636993656
transform 1 0 42964 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1636993656
transform 1 0 44068 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 25201
transform 1 0 45172 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 25201
transform 1 0 45724 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1636993656
transform 1 0 45908 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1636993656
transform 1 0 47012 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1636993656
transform 1 0 48116 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1636993656
transform 1 0 49220 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 25201
transform 1 0 50324 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 25201
transform 1 0 50876 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1636993656
transform 1 0 51060 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1636993656
transform 1 0 52164 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1636993656
transform 1 0 53268 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1636993656
transform 1 0 54372 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 25201
transform 1 0 55476 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 25201
transform 1 0 56028 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1636993656
transform 1 0 56212 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1636993656
transform 1 0 57316 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1636993656
transform 1 0 58420 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1636993656
transform 1 0 59524 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 25201
transform 1 0 60628 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 25201
transform 1 0 61180 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1636993656
transform 1 0 61364 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1636993656
transform 1 0 62468 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1636993656
transform 1 0 63572 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1636993656
transform 1 0 64676 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 25201
transform 1 0 65780 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 25201
transform 1 0 66332 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1636993656
transform 1 0 66516 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1636993656
transform 1 0 67620 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_725
timestamp 1636993656
transform 1 0 68724 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_737
timestamp 1636993656
transform 1 0 69828 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_749
timestamp 25201
transform 1 0 70932 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_755
timestamp 25201
transform 1 0 71484 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_757
timestamp 1636993656
transform 1 0 71668 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_769
timestamp 1636993656
transform 1 0 72772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_781
timestamp 1636993656
transform 1 0 73876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_793
timestamp 1636993656
transform 1 0 74980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_805
timestamp 25201
transform 1 0 76084 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_811
timestamp 25201
transform 1 0 76636 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_813
timestamp 25201
transform 1 0 76820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_821
timestamp 25201
transform 1 0 77556 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636993656
transform 1 0 2300 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636993656
transform 1 0 3404 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1636993656
transform 1 0 4508 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1636993656
transform 1 0 5612 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 25201
transform 1 0 6716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 25201
transform 1 0 7084 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636993656
transform 1 0 7268 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1636993656
transform 1 0 8372 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1636993656
transform 1 0 9476 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1636993656
transform 1 0 10580 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 25201
transform 1 0 11684 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 25201
transform 1 0 12236 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1636993656
transform 1 0 12420 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1636993656
transform 1 0 13524 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1636993656
transform 1 0 14628 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1636993656
transform 1 0 15732 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 25201
transform 1 0 16836 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 25201
transform 1 0 17388 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1636993656
transform 1 0 17572 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1636993656
transform 1 0 18676 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1636993656
transform 1 0 19780 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1636993656
transform 1 0 20884 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 25201
transform 1 0 21988 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 25201
transform 1 0 22540 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1636993656
transform 1 0 22724 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1636993656
transform 1 0 23828 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1636993656
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1636993656
transform 1 0 26036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 25201
transform 1 0 27140 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 25201
transform 1 0 27692 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1636993656
transform 1 0 27876 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1636993656
transform 1 0 28980 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1636993656
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1636993656
transform 1 0 31188 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 25201
transform 1 0 32292 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 25201
transform 1 0 32844 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1636993656
transform 1 0 33028 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1636993656
transform 1 0 34132 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1636993656
transform 1 0 35236 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1636993656
transform 1 0 36340 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 25201
transform 1 0 37444 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 25201
transform 1 0 37996 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1636993656
transform 1 0 38180 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1636993656
transform 1 0 39284 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1636993656
transform 1 0 40388 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1636993656
transform 1 0 41492 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 25201
transform 1 0 42596 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 25201
transform 1 0 43148 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1636993656
transform 1 0 43332 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1636993656
transform 1 0 44436 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1636993656
transform 1 0 45540 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1636993656
transform 1 0 46644 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 25201
transform 1 0 47748 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 25201
transform 1 0 48300 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1636993656
transform 1 0 48484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1636993656
transform 1 0 49588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1636993656
transform 1 0 50692 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1636993656
transform 1 0 51796 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 25201
transform 1 0 52900 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 25201
transform 1 0 53452 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1636993656
transform 1 0 53636 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1636993656
transform 1 0 54740 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1636993656
transform 1 0 55844 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1636993656
transform 1 0 56948 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 25201
transform 1 0 58052 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 25201
transform 1 0 58604 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1636993656
transform 1 0 58788 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1636993656
transform 1 0 59892 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1636993656
transform 1 0 60996 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1636993656
transform 1 0 62100 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 25201
transform 1 0 63204 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 25201
transform 1 0 63756 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1636993656
transform 1 0 63940 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1636993656
transform 1 0 65044 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1636993656
transform 1 0 66148 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1636993656
transform 1 0 67252 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 25201
transform 1 0 68356 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 25201
transform 1 0 68908 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_729
timestamp 1636993656
transform 1 0 69092 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_741
timestamp 1636993656
transform 1 0 70196 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_753
timestamp 1636993656
transform 1 0 71300 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_765
timestamp 1636993656
transform 1 0 72404 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_777
timestamp 25201
transform 1 0 73508 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_783
timestamp 25201
transform 1 0 74060 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_785
timestamp 1636993656
transform 1 0 74244 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_797
timestamp 1636993656
transform 1 0 75348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_809
timestamp 1636993656
transform 1 0 76452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_821
timestamp 25201
transform 1 0 77556 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636993656
transform 1 0 2300 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636993656
transform 1 0 3404 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 25201
transform 1 0 4508 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636993656
transform 1 0 4692 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1636993656
transform 1 0 5796 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1636993656
transform 1 0 6900 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1636993656
transform 1 0 8004 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 25201
transform 1 0 9108 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 25201
transform 1 0 9660 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1636993656
transform 1 0 9844 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1636993656
transform 1 0 10948 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1636993656
transform 1 0 12052 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1636993656
transform 1 0 13156 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 25201
transform 1 0 14260 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 25201
transform 1 0 14812 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1636993656
transform 1 0 14996 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1636993656
transform 1 0 16100 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1636993656
transform 1 0 17204 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1636993656
transform 1 0 18308 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 25201
transform 1 0 19412 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 25201
transform 1 0 19964 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1636993656
transform 1 0 20148 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1636993656
transform 1 0 21252 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1636993656
transform 1 0 22356 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1636993656
transform 1 0 23460 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 25201
transform 1 0 24564 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 25201
transform 1 0 25116 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1636993656
transform 1 0 25300 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1636993656
transform 1 0 26404 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1636993656
transform 1 0 27508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1636993656
transform 1 0 28612 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 25201
transform 1 0 29716 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 25201
transform 1 0 30268 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1636993656
transform 1 0 30452 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1636993656
transform 1 0 31556 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1636993656
transform 1 0 32660 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1636993656
transform 1 0 33764 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 25201
transform 1 0 34868 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 25201
transform 1 0 35420 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1636993656
transform 1 0 35604 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1636993656
transform 1 0 36708 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1636993656
transform 1 0 37812 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1636993656
transform 1 0 38916 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 25201
transform 1 0 40020 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 25201
transform 1 0 40572 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1636993656
transform 1 0 40756 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1636993656
transform 1 0 41860 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1636993656
transform 1 0 42964 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1636993656
transform 1 0 44068 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 25201
transform 1 0 45172 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 25201
transform 1 0 45724 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1636993656
transform 1 0 45908 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1636993656
transform 1 0 47012 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1636993656
transform 1 0 48116 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1636993656
transform 1 0 49220 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 25201
transform 1 0 50324 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 25201
transform 1 0 50876 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1636993656
transform 1 0 51060 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1636993656
transform 1 0 52164 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1636993656
transform 1 0 53268 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1636993656
transform 1 0 54372 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 25201
transform 1 0 55476 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 25201
transform 1 0 56028 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1636993656
transform 1 0 56212 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1636993656
transform 1 0 57316 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1636993656
transform 1 0 58420 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1636993656
transform 1 0 59524 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 25201
transform 1 0 60628 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 25201
transform 1 0 61180 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1636993656
transform 1 0 61364 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1636993656
transform 1 0 62468 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1636993656
transform 1 0 63572 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1636993656
transform 1 0 64676 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 25201
transform 1 0 65780 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 25201
transform 1 0 66332 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1636993656
transform 1 0 66516 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1636993656
transform 1 0 67620 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_725
timestamp 1636993656
transform 1 0 68724 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_737
timestamp 1636993656
transform 1 0 69828 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_749
timestamp 25201
transform 1 0 70932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_755
timestamp 25201
transform 1 0 71484 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_757
timestamp 1636993656
transform 1 0 71668 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_769
timestamp 1636993656
transform 1 0 72772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_781
timestamp 1636993656
transform 1 0 73876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_793
timestamp 1636993656
transform 1 0 74980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_805
timestamp 25201
transform 1 0 76084 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_811
timestamp 25201
transform 1 0 76636 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_813
timestamp 25201
transform 1 0 76820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_821
timestamp 25201
transform 1 0 77556 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1636993656
transform 1 0 2300 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1636993656
transform 1 0 3404 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1636993656
transform 1 0 4508 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1636993656
transform 1 0 5612 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 25201
transform 1 0 6716 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 25201
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636993656
transform 1 0 7268 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1636993656
transform 1 0 8372 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1636993656
transform 1 0 9476 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1636993656
transform 1 0 10580 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 25201
transform 1 0 11684 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 25201
transform 1 0 12236 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1636993656
transform 1 0 12420 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1636993656
transform 1 0 13524 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1636993656
transform 1 0 14628 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1636993656
transform 1 0 15732 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 25201
transform 1 0 16836 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 25201
transform 1 0 17388 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1636993656
transform 1 0 17572 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1636993656
transform 1 0 18676 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1636993656
transform 1 0 19780 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1636993656
transform 1 0 20884 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 25201
transform 1 0 21988 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 25201
transform 1 0 22540 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1636993656
transform 1 0 22724 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1636993656
transform 1 0 23828 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1636993656
transform 1 0 24932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1636993656
transform 1 0 26036 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 25201
transform 1 0 27140 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 25201
transform 1 0 27692 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1636993656
transform 1 0 27876 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1636993656
transform 1 0 28980 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1636993656
transform 1 0 30084 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1636993656
transform 1 0 31188 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 25201
transform 1 0 32292 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 25201
transform 1 0 32844 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1636993656
transform 1 0 33028 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1636993656
transform 1 0 34132 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1636993656
transform 1 0 35236 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1636993656
transform 1 0 36340 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 25201
transform 1 0 37444 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 25201
transform 1 0 37996 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1636993656
transform 1 0 38180 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1636993656
transform 1 0 39284 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1636993656
transform 1 0 40388 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1636993656
transform 1 0 41492 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 25201
transform 1 0 42596 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 25201
transform 1 0 43148 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1636993656
transform 1 0 43332 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1636993656
transform 1 0 44436 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1636993656
transform 1 0 45540 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1636993656
transform 1 0 46644 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 25201
transform 1 0 47748 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 25201
transform 1 0 48300 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1636993656
transform 1 0 48484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1636993656
transform 1 0 49588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1636993656
transform 1 0 50692 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1636993656
transform 1 0 51796 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 25201
transform 1 0 52900 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 25201
transform 1 0 53452 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1636993656
transform 1 0 53636 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1636993656
transform 1 0 54740 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1636993656
transform 1 0 55844 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1636993656
transform 1 0 56948 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 25201
transform 1 0 58052 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 25201
transform 1 0 58604 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1636993656
transform 1 0 58788 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1636993656
transform 1 0 59892 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1636993656
transform 1 0 60996 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1636993656
transform 1 0 62100 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 25201
transform 1 0 63204 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 25201
transform 1 0 63756 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1636993656
transform 1 0 63940 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1636993656
transform 1 0 65044 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1636993656
transform 1 0 66148 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1636993656
transform 1 0 67252 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 25201
transform 1 0 68356 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 25201
transform 1 0 68908 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_729
timestamp 1636993656
transform 1 0 69092 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_741
timestamp 1636993656
transform 1 0 70196 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_753
timestamp 1636993656
transform 1 0 71300 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_765
timestamp 1636993656
transform 1 0 72404 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_777
timestamp 25201
transform 1 0 73508 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_783
timestamp 25201
transform 1 0 74060 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_785
timestamp 1636993656
transform 1 0 74244 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_797
timestamp 1636993656
transform 1 0 75348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_809
timestamp 1636993656
transform 1 0 76452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_821
timestamp 25201
transform 1 0 77556 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636993656
transform 1 0 2300 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636993656
transform 1 0 3404 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 25201
transform 1 0 4508 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636993656
transform 1 0 4692 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636993656
transform 1 0 5796 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636993656
transform 1 0 6900 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1636993656
transform 1 0 8004 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 25201
transform 1 0 9108 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 25201
transform 1 0 9660 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1636993656
transform 1 0 9844 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1636993656
transform 1 0 10948 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1636993656
transform 1 0 12052 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1636993656
transform 1 0 13156 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 25201
transform 1 0 14260 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 25201
transform 1 0 14812 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1636993656
transform 1 0 14996 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1636993656
transform 1 0 16100 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1636993656
transform 1 0 17204 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1636993656
transform 1 0 18308 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 25201
transform 1 0 19412 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 25201
transform 1 0 19964 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1636993656
transform 1 0 20148 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1636993656
transform 1 0 21252 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1636993656
transform 1 0 22356 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1636993656
transform 1 0 23460 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 25201
transform 1 0 24564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 25201
transform 1 0 25116 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1636993656
transform 1 0 25300 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1636993656
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1636993656
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1636993656
transform 1 0 28612 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 25201
transform 1 0 29716 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 25201
transform 1 0 30268 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1636993656
transform 1 0 30452 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1636993656
transform 1 0 31556 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1636993656
transform 1 0 32660 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1636993656
transform 1 0 33764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 25201
transform 1 0 34868 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 25201
transform 1 0 35420 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1636993656
transform 1 0 35604 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1636993656
transform 1 0 36708 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1636993656
transform 1 0 37812 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1636993656
transform 1 0 38916 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 25201
transform 1 0 40020 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 25201
transform 1 0 40572 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1636993656
transform 1 0 40756 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1636993656
transform 1 0 41860 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1636993656
transform 1 0 42964 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1636993656
transform 1 0 44068 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 25201
transform 1 0 45172 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 25201
transform 1 0 45724 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1636993656
transform 1 0 45908 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1636993656
transform 1 0 47012 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1636993656
transform 1 0 48116 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1636993656
transform 1 0 49220 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 25201
transform 1 0 50324 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 25201
transform 1 0 50876 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1636993656
transform 1 0 51060 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1636993656
transform 1 0 52164 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1636993656
transform 1 0 53268 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1636993656
transform 1 0 54372 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 25201
transform 1 0 55476 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 25201
transform 1 0 56028 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1636993656
transform 1 0 56212 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1636993656
transform 1 0 57316 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1636993656
transform 1 0 58420 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1636993656
transform 1 0 59524 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 25201
transform 1 0 60628 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 25201
transform 1 0 61180 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1636993656
transform 1 0 61364 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1636993656
transform 1 0 62468 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1636993656
transform 1 0 63572 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1636993656
transform 1 0 64676 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 25201
transform 1 0 65780 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 25201
transform 1 0 66332 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1636993656
transform 1 0 66516 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1636993656
transform 1 0 67620 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_725
timestamp 1636993656
transform 1 0 68724 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_737
timestamp 1636993656
transform 1 0 69828 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_749
timestamp 25201
transform 1 0 70932 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_755
timestamp 25201
transform 1 0 71484 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_757
timestamp 1636993656
transform 1 0 71668 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_769
timestamp 1636993656
transform 1 0 72772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_781
timestamp 1636993656
transform 1 0 73876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_793
timestamp 1636993656
transform 1 0 74980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_805
timestamp 25201
transform 1 0 76084 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_811
timestamp 25201
transform 1 0 76636 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_813
timestamp 25201
transform 1 0 76820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_821
timestamp 25201
transform 1 0 77556 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636993656
transform 1 0 2300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636993656
transform 1 0 3404 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636993656
transform 1 0 4508 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1636993656
transform 1 0 5612 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 25201
transform 1 0 6716 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 25201
transform 1 0 7084 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636993656
transform 1 0 7268 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1636993656
transform 1 0 8372 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1636993656
transform 1 0 9476 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1636993656
transform 1 0 10580 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 25201
transform 1 0 11684 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 25201
transform 1 0 12236 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1636993656
transform 1 0 12420 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1636993656
transform 1 0 13524 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1636993656
transform 1 0 14628 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1636993656
transform 1 0 15732 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 25201
transform 1 0 16836 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 25201
transform 1 0 17388 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1636993656
transform 1 0 17572 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1636993656
transform 1 0 18676 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1636993656
transform 1 0 19780 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1636993656
transform 1 0 20884 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 25201
transform 1 0 21988 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 25201
transform 1 0 22540 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1636993656
transform 1 0 22724 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1636993656
transform 1 0 23828 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1636993656
transform 1 0 24932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1636993656
transform 1 0 26036 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 25201
transform 1 0 27140 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 25201
transform 1 0 27692 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1636993656
transform 1 0 27876 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1636993656
transform 1 0 28980 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1636993656
transform 1 0 30084 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1636993656
transform 1 0 31188 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 25201
transform 1 0 32292 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 25201
transform 1 0 32844 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1636993656
transform 1 0 33028 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1636993656
transform 1 0 34132 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1636993656
transform 1 0 35236 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1636993656
transform 1 0 36340 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 25201
transform 1 0 37444 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 25201
transform 1 0 37996 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1636993656
transform 1 0 38180 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1636993656
transform 1 0 39284 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1636993656
transform 1 0 40388 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1636993656
transform 1 0 41492 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 25201
transform 1 0 42596 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 25201
transform 1 0 43148 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1636993656
transform 1 0 43332 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1636993656
transform 1 0 44436 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1636993656
transform 1 0 45540 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1636993656
transform 1 0 46644 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 25201
transform 1 0 47748 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 25201
transform 1 0 48300 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1636993656
transform 1 0 48484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1636993656
transform 1 0 49588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1636993656
transform 1 0 50692 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1636993656
transform 1 0 51796 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 25201
transform 1 0 52900 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 25201
transform 1 0 53452 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1636993656
transform 1 0 53636 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1636993656
transform 1 0 54740 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1636993656
transform 1 0 55844 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1636993656
transform 1 0 56948 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 25201
transform 1 0 58052 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 25201
transform 1 0 58604 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1636993656
transform 1 0 58788 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1636993656
transform 1 0 59892 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1636993656
transform 1 0 60996 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1636993656
transform 1 0 62100 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 25201
transform 1 0 63204 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 25201
transform 1 0 63756 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1636993656
transform 1 0 63940 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1636993656
transform 1 0 65044 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1636993656
transform 1 0 66148 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1636993656
transform 1 0 67252 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 25201
transform 1 0 68356 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 25201
transform 1 0 68908 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_729
timestamp 1636993656
transform 1 0 69092 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_741
timestamp 1636993656
transform 1 0 70196 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_753
timestamp 1636993656
transform 1 0 71300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_765
timestamp 1636993656
transform 1 0 72404 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_777
timestamp 25201
transform 1 0 73508 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_783
timestamp 25201
transform 1 0 74060 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_785
timestamp 1636993656
transform 1 0 74244 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_797
timestamp 1636993656
transform 1 0 75348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_809
timestamp 1636993656
transform 1 0 76452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_821
timestamp 25201
transform 1 0 77556 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636993656
transform 1 0 2300 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636993656
transform 1 0 3404 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 25201
transform 1 0 4508 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636993656
transform 1 0 4692 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636993656
transform 1 0 5796 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1636993656
transform 1 0 6900 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1636993656
transform 1 0 8004 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 25201
transform 1 0 9108 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 25201
transform 1 0 9660 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1636993656
transform 1 0 9844 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1636993656
transform 1 0 10948 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1636993656
transform 1 0 12052 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1636993656
transform 1 0 13156 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 25201
transform 1 0 14260 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 25201
transform 1 0 14812 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1636993656
transform 1 0 14996 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1636993656
transform 1 0 16100 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1636993656
transform 1 0 17204 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1636993656
transform 1 0 18308 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 25201
transform 1 0 19412 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 25201
transform 1 0 19964 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1636993656
transform 1 0 20148 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1636993656
transform 1 0 21252 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1636993656
transform 1 0 22356 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1636993656
transform 1 0 23460 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 25201
transform 1 0 24564 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 25201
transform 1 0 25116 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1636993656
transform 1 0 25300 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1636993656
transform 1 0 26404 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1636993656
transform 1 0 27508 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1636993656
transform 1 0 28612 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 25201
transform 1 0 29716 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 25201
transform 1 0 30268 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1636993656
transform 1 0 30452 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1636993656
transform 1 0 31556 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1636993656
transform 1 0 32660 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1636993656
transform 1 0 33764 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 25201
transform 1 0 34868 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 25201
transform 1 0 35420 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1636993656
transform 1 0 35604 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1636993656
transform 1 0 36708 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1636993656
transform 1 0 37812 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1636993656
transform 1 0 38916 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 25201
transform 1 0 40020 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 25201
transform 1 0 40572 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1636993656
transform 1 0 40756 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1636993656
transform 1 0 41860 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1636993656
transform 1 0 42964 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1636993656
transform 1 0 44068 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 25201
transform 1 0 45172 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 25201
transform 1 0 45724 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1636993656
transform 1 0 45908 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1636993656
transform 1 0 47012 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1636993656
transform 1 0 48116 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1636993656
transform 1 0 49220 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 25201
transform 1 0 50324 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 25201
transform 1 0 50876 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1636993656
transform 1 0 51060 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1636993656
transform 1 0 52164 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1636993656
transform 1 0 53268 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1636993656
transform 1 0 54372 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 25201
transform 1 0 55476 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 25201
transform 1 0 56028 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1636993656
transform 1 0 56212 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1636993656
transform 1 0 57316 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1636993656
transform 1 0 58420 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1636993656
transform 1 0 59524 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 25201
transform 1 0 60628 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 25201
transform 1 0 61180 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1636993656
transform 1 0 61364 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1636993656
transform 1 0 62468 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1636993656
transform 1 0 63572 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1636993656
transform 1 0 64676 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 25201
transform 1 0 65780 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 25201
transform 1 0 66332 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1636993656
transform 1 0 66516 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1636993656
transform 1 0 67620 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_725
timestamp 1636993656
transform 1 0 68724 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_737
timestamp 1636993656
transform 1 0 69828 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_749
timestamp 25201
transform 1 0 70932 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_755
timestamp 25201
transform 1 0 71484 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_757
timestamp 1636993656
transform 1 0 71668 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_769
timestamp 1636993656
transform 1 0 72772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_781
timestamp 1636993656
transform 1 0 73876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_793
timestamp 1636993656
transform 1 0 74980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_805
timestamp 25201
transform 1 0 76084 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_811
timestamp 25201
transform 1 0 76636 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_813
timestamp 25201
transform 1 0 76820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_821
timestamp 25201
transform 1 0 77556 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636993656
transform 1 0 2300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636993656
transform 1 0 3404 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1636993656
transform 1 0 4508 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1636993656
transform 1 0 5612 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 25201
transform 1 0 6716 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 25201
transform 1 0 7084 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636993656
transform 1 0 7268 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1636993656
transform 1 0 8372 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1636993656
transform 1 0 9476 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1636993656
transform 1 0 10580 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 25201
transform 1 0 11684 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 25201
transform 1 0 12236 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1636993656
transform 1 0 12420 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1636993656
transform 1 0 13524 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1636993656
transform 1 0 14628 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1636993656
transform 1 0 15732 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 25201
transform 1 0 16836 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 25201
transform 1 0 17388 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1636993656
transform 1 0 17572 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1636993656
transform 1 0 18676 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1636993656
transform 1 0 19780 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1636993656
transform 1 0 20884 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 25201
transform 1 0 21988 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 25201
transform 1 0 22540 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1636993656
transform 1 0 22724 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1636993656
transform 1 0 23828 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1636993656
transform 1 0 24932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1636993656
transform 1 0 26036 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 25201
transform 1 0 27140 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 25201
transform 1 0 27692 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1636993656
transform 1 0 27876 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1636993656
transform 1 0 28980 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1636993656
transform 1 0 30084 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1636993656
transform 1 0 31188 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 25201
transform 1 0 32292 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 25201
transform 1 0 32844 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1636993656
transform 1 0 33028 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1636993656
transform 1 0 34132 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1636993656
transform 1 0 35236 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1636993656
transform 1 0 36340 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 25201
transform 1 0 37444 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 25201
transform 1 0 37996 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1636993656
transform 1 0 38180 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1636993656
transform 1 0 39284 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1636993656
transform 1 0 40388 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1636993656
transform 1 0 41492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 25201
transform 1 0 42596 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 25201
transform 1 0 43148 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1636993656
transform 1 0 43332 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1636993656
transform 1 0 44436 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1636993656
transform 1 0 45540 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1636993656
transform 1 0 46644 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 25201
transform 1 0 47748 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 25201
transform 1 0 48300 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1636993656
transform 1 0 48484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1636993656
transform 1 0 49588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1636993656
transform 1 0 50692 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1636993656
transform 1 0 51796 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 25201
transform 1 0 52900 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 25201
transform 1 0 53452 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1636993656
transform 1 0 53636 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1636993656
transform 1 0 54740 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1636993656
transform 1 0 55844 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1636993656
transform 1 0 56948 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 25201
transform 1 0 58052 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 25201
transform 1 0 58604 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1636993656
transform 1 0 58788 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1636993656
transform 1 0 59892 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1636993656
transform 1 0 60996 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1636993656
transform 1 0 62100 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 25201
transform 1 0 63204 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 25201
transform 1 0 63756 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1636993656
transform 1 0 63940 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1636993656
transform 1 0 65044 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1636993656
transform 1 0 66148 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1636993656
transform 1 0 67252 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 25201
transform 1 0 68356 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 25201
transform 1 0 68908 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_729
timestamp 1636993656
transform 1 0 69092 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_741
timestamp 1636993656
transform 1 0 70196 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_753
timestamp 1636993656
transform 1 0 71300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_765
timestamp 1636993656
transform 1 0 72404 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_777
timestamp 25201
transform 1 0 73508 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_783
timestamp 25201
transform 1 0 74060 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_785
timestamp 1636993656
transform 1 0 74244 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_797
timestamp 1636993656
transform 1 0 75348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_809
timestamp 1636993656
transform 1 0 76452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_821
timestamp 25201
transform 1 0 77556 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636993656
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636993656
transform 1 0 3404 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 25201
transform 1 0 4508 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636993656
transform 1 0 4692 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636993656
transform 1 0 5796 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636993656
transform 1 0 6900 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1636993656
transform 1 0 8004 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 25201
transform 1 0 9108 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 25201
transform 1 0 9660 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1636993656
transform 1 0 9844 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1636993656
transform 1 0 10948 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1636993656
transform 1 0 12052 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1636993656
transform 1 0 13156 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 25201
transform 1 0 14260 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 25201
transform 1 0 14812 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1636993656
transform 1 0 14996 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1636993656
transform 1 0 16100 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1636993656
transform 1 0 17204 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1636993656
transform 1 0 18308 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 25201
transform 1 0 19412 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 25201
transform 1 0 19964 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1636993656
transform 1 0 20148 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1636993656
transform 1 0 21252 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1636993656
transform 1 0 22356 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1636993656
transform 1 0 23460 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 25201
transform 1 0 24564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 25201
transform 1 0 25116 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1636993656
transform 1 0 25300 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1636993656
transform 1 0 26404 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1636993656
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1636993656
transform 1 0 28612 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 25201
transform 1 0 29716 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 25201
transform 1 0 30268 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1636993656
transform 1 0 30452 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1636993656
transform 1 0 31556 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1636993656
transform 1 0 32660 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1636993656
transform 1 0 33764 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 25201
transform 1 0 34868 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 25201
transform 1 0 35420 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1636993656
transform 1 0 35604 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1636993656
transform 1 0 36708 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1636993656
transform 1 0 37812 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1636993656
transform 1 0 38916 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 25201
transform 1 0 40020 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 25201
transform 1 0 40572 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1636993656
transform 1 0 40756 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1636993656
transform 1 0 41860 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1636993656
transform 1 0 42964 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1636993656
transform 1 0 44068 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 25201
transform 1 0 45172 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 25201
transform 1 0 45724 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1636993656
transform 1 0 45908 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1636993656
transform 1 0 47012 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1636993656
transform 1 0 48116 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1636993656
transform 1 0 49220 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 25201
transform 1 0 50324 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 25201
transform 1 0 50876 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1636993656
transform 1 0 51060 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1636993656
transform 1 0 52164 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1636993656
transform 1 0 53268 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1636993656
transform 1 0 54372 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 25201
transform 1 0 55476 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 25201
transform 1 0 56028 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1636993656
transform 1 0 56212 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1636993656
transform 1 0 57316 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1636993656
transform 1 0 58420 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1636993656
transform 1 0 59524 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 25201
transform 1 0 60628 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 25201
transform 1 0 61180 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1636993656
transform 1 0 61364 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1636993656
transform 1 0 62468 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1636993656
transform 1 0 63572 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_681
timestamp 1636993656
transform 1 0 64676 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 25201
transform 1 0 65780 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 25201
transform 1 0 66332 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1636993656
transform 1 0 66516 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1636993656
transform 1 0 67620 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_725
timestamp 1636993656
transform 1 0 68724 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_737
timestamp 1636993656
transform 1 0 69828 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_749
timestamp 25201
transform 1 0 70932 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_755
timestamp 25201
transform 1 0 71484 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_757
timestamp 1636993656
transform 1 0 71668 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_769
timestamp 1636993656
transform 1 0 72772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_781
timestamp 1636993656
transform 1 0 73876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_793
timestamp 1636993656
transform 1 0 74980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_805
timestamp 25201
transform 1 0 76084 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_811
timestamp 25201
transform 1 0 76636 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_813
timestamp 25201
transform 1 0 76820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_821
timestamp 25201
transform 1 0 77556 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636993656
transform 1 0 2300 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636993656
transform 1 0 3404 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636993656
transform 1 0 4508 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636993656
transform 1 0 5612 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 25201
transform 1 0 6716 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 25201
transform 1 0 7084 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636993656
transform 1 0 7268 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1636993656
transform 1 0 8372 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1636993656
transform 1 0 9476 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1636993656
transform 1 0 10580 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 25201
transform 1 0 11684 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 25201
transform 1 0 12236 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1636993656
transform 1 0 12420 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1636993656
transform 1 0 13524 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1636993656
transform 1 0 14628 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1636993656
transform 1 0 15732 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 25201
transform 1 0 16836 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 25201
transform 1 0 17388 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1636993656
transform 1 0 17572 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1636993656
transform 1 0 18676 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1636993656
transform 1 0 19780 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1636993656
transform 1 0 20884 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 25201
transform 1 0 21988 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 25201
transform 1 0 22540 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1636993656
transform 1 0 22724 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1636993656
transform 1 0 23828 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1636993656
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1636993656
transform 1 0 26036 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 25201
transform 1 0 27140 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 25201
transform 1 0 27692 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1636993656
transform 1 0 27876 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1636993656
transform 1 0 28980 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1636993656
transform 1 0 30084 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1636993656
transform 1 0 31188 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 25201
transform 1 0 32292 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 25201
transform 1 0 32844 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1636993656
transform 1 0 33028 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1636993656
transform 1 0 34132 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1636993656
transform 1 0 35236 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1636993656
transform 1 0 36340 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 25201
transform 1 0 37444 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 25201
transform 1 0 37996 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1636993656
transform 1 0 38180 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1636993656
transform 1 0 39284 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1636993656
transform 1 0 40388 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1636993656
transform 1 0 41492 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 25201
transform 1 0 42596 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 25201
transform 1 0 43148 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1636993656
transform 1 0 43332 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1636993656
transform 1 0 44436 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1636993656
transform 1 0 45540 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1636993656
transform 1 0 46644 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 25201
transform 1 0 47748 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 25201
transform 1 0 48300 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1636993656
transform 1 0 48484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1636993656
transform 1 0 49588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1636993656
transform 1 0 50692 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1636993656
transform 1 0 51796 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 25201
transform 1 0 52900 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 25201
transform 1 0 53452 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1636993656
transform 1 0 53636 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1636993656
transform 1 0 54740 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1636993656
transform 1 0 55844 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1636993656
transform 1 0 56948 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 25201
transform 1 0 58052 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 25201
transform 1 0 58604 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1636993656
transform 1 0 58788 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1636993656
transform 1 0 59892 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1636993656
transform 1 0 60996 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1636993656
transform 1 0 62100 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 25201
transform 1 0 63204 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 25201
transform 1 0 63756 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1636993656
transform 1 0 63940 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1636993656
transform 1 0 65044 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1636993656
transform 1 0 66148 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1636993656
transform 1 0 67252 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 25201
transform 1 0 68356 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 25201
transform 1 0 68908 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_729
timestamp 1636993656
transform 1 0 69092 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_741
timestamp 1636993656
transform 1 0 70196 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_753
timestamp 1636993656
transform 1 0 71300 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_765
timestamp 1636993656
transform 1 0 72404 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_777
timestamp 25201
transform 1 0 73508 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_783
timestamp 25201
transform 1 0 74060 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_785
timestamp 1636993656
transform 1 0 74244 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_797
timestamp 1636993656
transform 1 0 75348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_809
timestamp 1636993656
transform 1 0 76452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_821
timestamp 25201
transform 1 0 77556 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636993656
transform 1 0 2300 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636993656
transform 1 0 3404 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 25201
transform 1 0 4508 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636993656
transform 1 0 4692 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636993656
transform 1 0 5796 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636993656
transform 1 0 6900 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1636993656
transform 1 0 8004 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 25201
transform 1 0 9108 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 25201
transform 1 0 9660 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1636993656
transform 1 0 9844 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1636993656
transform 1 0 10948 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1636993656
transform 1 0 12052 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1636993656
transform 1 0 13156 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 25201
transform 1 0 14260 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 25201
transform 1 0 14812 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1636993656
transform 1 0 14996 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1636993656
transform 1 0 16100 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1636993656
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1636993656
transform 1 0 18308 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 25201
transform 1 0 19412 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 25201
transform 1 0 19964 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1636993656
transform 1 0 20148 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1636993656
transform 1 0 21252 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1636993656
transform 1 0 22356 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1636993656
transform 1 0 23460 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 25201
transform 1 0 24564 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 25201
transform 1 0 25116 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1636993656
transform 1 0 25300 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1636993656
transform 1 0 26404 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1636993656
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1636993656
transform 1 0 28612 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 25201
transform 1 0 29716 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 25201
transform 1 0 30268 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1636993656
transform 1 0 30452 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1636993656
transform 1 0 31556 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1636993656
transform 1 0 32660 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1636993656
transform 1 0 33764 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 25201
transform 1 0 34868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 25201
transform 1 0 35420 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1636993656
transform 1 0 35604 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1636993656
transform 1 0 36708 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1636993656
transform 1 0 37812 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1636993656
transform 1 0 38916 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 25201
transform 1 0 40020 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 25201
transform 1 0 40572 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1636993656
transform 1 0 40756 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1636993656
transform 1 0 41860 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1636993656
transform 1 0 42964 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1636993656
transform 1 0 44068 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 25201
transform 1 0 45172 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 25201
transform 1 0 45724 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1636993656
transform 1 0 45908 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1636993656
transform 1 0 47012 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1636993656
transform 1 0 48116 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1636993656
transform 1 0 49220 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 25201
transform 1 0 50324 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 25201
transform 1 0 50876 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1636993656
transform 1 0 51060 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1636993656
transform 1 0 52164 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1636993656
transform 1 0 53268 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1636993656
transform 1 0 54372 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 25201
transform 1 0 55476 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 25201
transform 1 0 56028 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1636993656
transform 1 0 56212 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1636993656
transform 1 0 57316 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1636993656
transform 1 0 58420 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1636993656
transform 1 0 59524 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 25201
transform 1 0 60628 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 25201
transform 1 0 61180 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1636993656
transform 1 0 61364 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1636993656
transform 1 0 62468 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1636993656
transform 1 0 63572 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1636993656
transform 1 0 64676 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 25201
transform 1 0 65780 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 25201
transform 1 0 66332 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1636993656
transform 1 0 66516 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1636993656
transform 1 0 67620 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_725
timestamp 1636993656
transform 1 0 68724 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_737
timestamp 1636993656
transform 1 0 69828 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_749
timestamp 25201
transform 1 0 70932 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_755
timestamp 25201
transform 1 0 71484 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_757
timestamp 1636993656
transform 1 0 71668 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_769
timestamp 1636993656
transform 1 0 72772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_781
timestamp 1636993656
transform 1 0 73876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_793
timestamp 1636993656
transform 1 0 74980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_805
timestamp 25201
transform 1 0 76084 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_811
timestamp 25201
transform 1 0 76636 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_813
timestamp 25201
transform 1 0 76820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_821
timestamp 25201
transform 1 0 77556 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636993656
transform 1 0 2300 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636993656
transform 1 0 3404 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636993656
transform 1 0 4508 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636993656
transform 1 0 5612 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 25201
transform 1 0 6716 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 25201
transform 1 0 7084 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636993656
transform 1 0 7268 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1636993656
transform 1 0 8372 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1636993656
transform 1 0 9476 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1636993656
transform 1 0 10580 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 25201
transform 1 0 11684 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 25201
transform 1 0 12236 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1636993656
transform 1 0 12420 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1636993656
transform 1 0 13524 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1636993656
transform 1 0 14628 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1636993656
transform 1 0 15732 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 25201
transform 1 0 16836 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 25201
transform 1 0 17388 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636993656
transform 1 0 17572 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1636993656
transform 1 0 18676 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1636993656
transform 1 0 19780 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1636993656
transform 1 0 20884 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 25201
transform 1 0 21988 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 25201
transform 1 0 22540 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1636993656
transform 1 0 22724 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1636993656
transform 1 0 23828 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1636993656
transform 1 0 24932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1636993656
transform 1 0 26036 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 25201
transform 1 0 27140 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 25201
transform 1 0 27692 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1636993656
transform 1 0 27876 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1636993656
transform 1 0 28980 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1636993656
transform 1 0 30084 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1636993656
transform 1 0 31188 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 25201
transform 1 0 32292 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 25201
transform 1 0 32844 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1636993656
transform 1 0 33028 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1636993656
transform 1 0 34132 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1636993656
transform 1 0 35236 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1636993656
transform 1 0 36340 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 25201
transform 1 0 37444 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 25201
transform 1 0 37996 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1636993656
transform 1 0 38180 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1636993656
transform 1 0 39284 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1636993656
transform 1 0 40388 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1636993656
transform 1 0 41492 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 25201
transform 1 0 42596 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 25201
transform 1 0 43148 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1636993656
transform 1 0 43332 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1636993656
transform 1 0 44436 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1636993656
transform 1 0 45540 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1636993656
transform 1 0 46644 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 25201
transform 1 0 47748 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 25201
transform 1 0 48300 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1636993656
transform 1 0 48484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1636993656
transform 1 0 49588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1636993656
transform 1 0 50692 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1636993656
transform 1 0 51796 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 25201
transform 1 0 52900 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 25201
transform 1 0 53452 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1636993656
transform 1 0 53636 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1636993656
transform 1 0 54740 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1636993656
transform 1 0 55844 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1636993656
transform 1 0 56948 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 25201
transform 1 0 58052 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 25201
transform 1 0 58604 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_617
timestamp 1636993656
transform 1 0 58788 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_629
timestamp 1636993656
transform 1 0 59892 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_641
timestamp 1636993656
transform 1 0 60996 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_653
timestamp 1636993656
transform 1 0 62100 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 25201
transform 1 0 63204 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 25201
transform 1 0 63756 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1636993656
transform 1 0 63940 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_685
timestamp 1636993656
transform 1 0 65044 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_697
timestamp 1636993656
transform 1 0 66148 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_709
timestamp 1636993656
transform 1 0 67252 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 25201
transform 1 0 68356 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 25201
transform 1 0 68908 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_729
timestamp 1636993656
transform 1 0 69092 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_741
timestamp 1636993656
transform 1 0 70196 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_753
timestamp 1636993656
transform 1 0 71300 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_765
timestamp 1636993656
transform 1 0 72404 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_777
timestamp 25201
transform 1 0 73508 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_783
timestamp 25201
transform 1 0 74060 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_785
timestamp 1636993656
transform 1 0 74244 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_797
timestamp 1636993656
transform 1 0 75348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_809
timestamp 1636993656
transform 1 0 76452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_821
timestamp 25201
transform 1 0 77556 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636993656
transform 1 0 2300 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636993656
transform 1 0 3404 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 25201
transform 1 0 4508 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636993656
transform 1 0 4692 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636993656
transform 1 0 5796 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1636993656
transform 1 0 6900 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1636993656
transform 1 0 8004 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 25201
transform 1 0 9108 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 25201
transform 1 0 9660 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1636993656
transform 1 0 9844 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1636993656
transform 1 0 10948 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1636993656
transform 1 0 12052 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1636993656
transform 1 0 13156 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 25201
transform 1 0 14260 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 25201
transform 1 0 14812 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1636993656
transform 1 0 14996 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1636993656
transform 1 0 16100 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1636993656
transform 1 0 17204 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1636993656
transform 1 0 18308 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 25201
transform 1 0 19412 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 25201
transform 1 0 19964 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1636993656
transform 1 0 20148 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1636993656
transform 1 0 21252 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1636993656
transform 1 0 22356 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1636993656
transform 1 0 23460 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 25201
transform 1 0 24564 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 25201
transform 1 0 25116 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1636993656
transform 1 0 25300 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1636993656
transform 1 0 26404 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1636993656
transform 1 0 27508 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1636993656
transform 1 0 28612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 25201
transform 1 0 29716 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 25201
transform 1 0 30268 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1636993656
transform 1 0 30452 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1636993656
transform 1 0 31556 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1636993656
transform 1 0 32660 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1636993656
transform 1 0 33764 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 25201
transform 1 0 34868 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 25201
transform 1 0 35420 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1636993656
transform 1 0 35604 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1636993656
transform 1 0 36708 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1636993656
transform 1 0 37812 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1636993656
transform 1 0 38916 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 25201
transform 1 0 40020 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 25201
transform 1 0 40572 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1636993656
transform 1 0 40756 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1636993656
transform 1 0 41860 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1636993656
transform 1 0 42964 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1636993656
transform 1 0 44068 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 25201
transform 1 0 45172 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 25201
transform 1 0 45724 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1636993656
transform 1 0 45908 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1636993656
transform 1 0 47012 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1636993656
transform 1 0 48116 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1636993656
transform 1 0 49220 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 25201
transform 1 0 50324 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 25201
transform 1 0 50876 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1636993656
transform 1 0 51060 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1636993656
transform 1 0 52164 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1636993656
transform 1 0 53268 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1636993656
transform 1 0 54372 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 25201
transform 1 0 55476 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 25201
transform 1 0 56028 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1636993656
transform 1 0 56212 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1636993656
transform 1 0 57316 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1636993656
transform 1 0 58420 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_625
timestamp 1636993656
transform 1 0 59524 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 25201
transform 1 0 60628 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 25201
transform 1 0 61180 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_645
timestamp 1636993656
transform 1 0 61364 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_657
timestamp 1636993656
transform 1 0 62468 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_669
timestamp 1636993656
transform 1 0 63572 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_681
timestamp 1636993656
transform 1 0 64676 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 25201
transform 1 0 65780 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 25201
transform 1 0 66332 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_701
timestamp 1636993656
transform 1 0 66516 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_713
timestamp 1636993656
transform 1 0 67620 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_725
timestamp 1636993656
transform 1 0 68724 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_737
timestamp 1636993656
transform 1 0 69828 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_749
timestamp 25201
transform 1 0 70932 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_755
timestamp 25201
transform 1 0 71484 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_757
timestamp 1636993656
transform 1 0 71668 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_769
timestamp 1636993656
transform 1 0 72772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_781
timestamp 1636993656
transform 1 0 73876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_793
timestamp 1636993656
transform 1 0 74980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_805
timestamp 25201
transform 1 0 76084 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_811
timestamp 25201
transform 1 0 76636 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_813
timestamp 25201
transform 1 0 76820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_821
timestamp 25201
transform 1 0 77556 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636993656
transform 1 0 2300 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636993656
transform 1 0 3404 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1636993656
transform 1 0 4508 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1636993656
transform 1 0 5612 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 25201
transform 1 0 6716 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 25201
transform 1 0 7084 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636993656
transform 1 0 7268 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1636993656
transform 1 0 8372 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1636993656
transform 1 0 9476 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1636993656
transform 1 0 10580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 25201
transform 1 0 11684 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 25201
transform 1 0 12236 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1636993656
transform 1 0 12420 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1636993656
transform 1 0 13524 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1636993656
transform 1 0 14628 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1636993656
transform 1 0 15732 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 25201
transform 1 0 16836 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 25201
transform 1 0 17388 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1636993656
transform 1 0 17572 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1636993656
transform 1 0 18676 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1636993656
transform 1 0 19780 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1636993656
transform 1 0 20884 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 25201
transform 1 0 21988 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 25201
transform 1 0 22540 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1636993656
transform 1 0 22724 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1636993656
transform 1 0 23828 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1636993656
transform 1 0 24932 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1636993656
transform 1 0 26036 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 25201
transform 1 0 27140 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 25201
transform 1 0 27692 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1636993656
transform 1 0 27876 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1636993656
transform 1 0 28980 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1636993656
transform 1 0 30084 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1636993656
transform 1 0 31188 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 25201
transform 1 0 32292 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 25201
transform 1 0 32844 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1636993656
transform 1 0 33028 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1636993656
transform 1 0 34132 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1636993656
transform 1 0 35236 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1636993656
transform 1 0 36340 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 25201
transform 1 0 37444 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 25201
transform 1 0 37996 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1636993656
transform 1 0 38180 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1636993656
transform 1 0 39284 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1636993656
transform 1 0 40388 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1636993656
transform 1 0 41492 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 25201
transform 1 0 42596 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 25201
transform 1 0 43148 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1636993656
transform 1 0 43332 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1636993656
transform 1 0 44436 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1636993656
transform 1 0 45540 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1636993656
transform 1 0 46644 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 25201
transform 1 0 47748 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 25201
transform 1 0 48300 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1636993656
transform 1 0 48484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1636993656
transform 1 0 49588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1636993656
transform 1 0 50692 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1636993656
transform 1 0 51796 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 25201
transform 1 0 52900 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 25201
transform 1 0 53452 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1636993656
transform 1 0 53636 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1636993656
transform 1 0 54740 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1636993656
transform 1 0 55844 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1636993656
transform 1 0 56948 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 25201
transform 1 0 58052 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 25201
transform 1 0 58604 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_617
timestamp 1636993656
transform 1 0 58788 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_629
timestamp 1636993656
transform 1 0 59892 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_641
timestamp 1636993656
transform 1 0 60996 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_653
timestamp 1636993656
transform 1 0 62100 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 25201
transform 1 0 63204 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 25201
transform 1 0 63756 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_673
timestamp 1636993656
transform 1 0 63940 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_685
timestamp 1636993656
transform 1 0 65044 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_697
timestamp 1636993656
transform 1 0 66148 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_709
timestamp 1636993656
transform 1 0 67252 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 25201
transform 1 0 68356 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 25201
transform 1 0 68908 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_729
timestamp 1636993656
transform 1 0 69092 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_741
timestamp 1636993656
transform 1 0 70196 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_753
timestamp 1636993656
transform 1 0 71300 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_765
timestamp 1636993656
transform 1 0 72404 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_777
timestamp 25201
transform 1 0 73508 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_783
timestamp 25201
transform 1 0 74060 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_785
timestamp 1636993656
transform 1 0 74244 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_797
timestamp 1636993656
transform 1 0 75348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_809
timestamp 1636993656
transform 1 0 76452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_821
timestamp 25201
transform 1 0 77556 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636993656
transform 1 0 2300 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636993656
transform 1 0 3404 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 25201
transform 1 0 4508 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636993656
transform 1 0 4692 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636993656
transform 1 0 5796 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1636993656
transform 1 0 6900 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1636993656
transform 1 0 8004 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 25201
transform 1 0 9108 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 25201
transform 1 0 9660 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1636993656
transform 1 0 9844 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1636993656
transform 1 0 10948 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1636993656
transform 1 0 12052 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1636993656
transform 1 0 13156 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 25201
transform 1 0 14260 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 25201
transform 1 0 14812 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1636993656
transform 1 0 14996 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1636993656
transform 1 0 16100 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1636993656
transform 1 0 17204 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1636993656
transform 1 0 18308 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 25201
transform 1 0 19412 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 25201
transform 1 0 19964 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1636993656
transform 1 0 20148 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1636993656
transform 1 0 21252 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1636993656
transform 1 0 22356 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1636993656
transform 1 0 23460 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 25201
transform 1 0 24564 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 25201
transform 1 0 25116 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1636993656
transform 1 0 25300 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1636993656
transform 1 0 26404 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1636993656
transform 1 0 27508 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1636993656
transform 1 0 28612 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 25201
transform 1 0 29716 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 25201
transform 1 0 30268 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1636993656
transform 1 0 30452 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1636993656
transform 1 0 31556 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1636993656
transform 1 0 32660 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1636993656
transform 1 0 33764 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 25201
transform 1 0 34868 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 25201
transform 1 0 35420 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1636993656
transform 1 0 35604 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1636993656
transform 1 0 36708 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1636993656
transform 1 0 37812 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1636993656
transform 1 0 38916 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 25201
transform 1 0 40020 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 25201
transform 1 0 40572 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1636993656
transform 1 0 40756 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1636993656
transform 1 0 41860 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1636993656
transform 1 0 42964 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1636993656
transform 1 0 44068 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 25201
transform 1 0 45172 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 25201
transform 1 0 45724 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1636993656
transform 1 0 45908 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1636993656
transform 1 0 47012 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1636993656
transform 1 0 48116 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1636993656
transform 1 0 49220 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 25201
transform 1 0 50324 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 25201
transform 1 0 50876 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1636993656
transform 1 0 51060 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1636993656
transform 1 0 52164 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1636993656
transform 1 0 53268 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1636993656
transform 1 0 54372 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 25201
transform 1 0 55476 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 25201
transform 1 0 56028 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1636993656
transform 1 0 56212 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1636993656
transform 1 0 57316 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1636993656
transform 1 0 58420 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_625
timestamp 1636993656
transform 1 0 59524 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 25201
transform 1 0 60628 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 25201
transform 1 0 61180 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_645
timestamp 1636993656
transform 1 0 61364 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_657
timestamp 1636993656
transform 1 0 62468 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_669
timestamp 1636993656
transform 1 0 63572 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_681
timestamp 1636993656
transform 1 0 64676 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 25201
transform 1 0 65780 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 25201
transform 1 0 66332 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_701
timestamp 1636993656
transform 1 0 66516 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_713
timestamp 1636993656
transform 1 0 67620 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_725
timestamp 1636993656
transform 1 0 68724 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_737
timestamp 1636993656
transform 1 0 69828 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_749
timestamp 25201
transform 1 0 70932 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_755
timestamp 25201
transform 1 0 71484 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_757
timestamp 1636993656
transform 1 0 71668 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_769
timestamp 1636993656
transform 1 0 72772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_781
timestamp 1636993656
transform 1 0 73876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_793
timestamp 1636993656
transform 1 0 74980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_805
timestamp 25201
transform 1 0 76084 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_811
timestamp 25201
transform 1 0 76636 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_813
timestamp 25201
transform 1 0 76820 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_821
timestamp 25201
transform 1 0 77556 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636993656
transform 1 0 2300 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1636993656
transform 1 0 3404 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1636993656
transform 1 0 4508 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1636993656
transform 1 0 5612 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 25201
transform 1 0 6716 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 25201
transform 1 0 7084 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1636993656
transform 1 0 7268 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1636993656
transform 1 0 8372 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1636993656
transform 1 0 9476 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1636993656
transform 1 0 10580 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 25201
transform 1 0 11684 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 25201
transform 1 0 12236 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1636993656
transform 1 0 12420 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1636993656
transform 1 0 13524 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1636993656
transform 1 0 14628 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1636993656
transform 1 0 15732 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 25201
transform 1 0 16836 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 25201
transform 1 0 17388 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1636993656
transform 1 0 17572 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1636993656
transform 1 0 18676 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1636993656
transform 1 0 19780 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1636993656
transform 1 0 20884 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 25201
transform 1 0 21988 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 25201
transform 1 0 22540 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1636993656
transform 1 0 22724 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1636993656
transform 1 0 23828 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1636993656
transform 1 0 24932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1636993656
transform 1 0 26036 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 25201
transform 1 0 27140 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 25201
transform 1 0 27692 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1636993656
transform 1 0 27876 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1636993656
transform 1 0 28980 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1636993656
transform 1 0 30084 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1636993656
transform 1 0 31188 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 25201
transform 1 0 32292 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 25201
transform 1 0 32844 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1636993656
transform 1 0 33028 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1636993656
transform 1 0 34132 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1636993656
transform 1 0 35236 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1636993656
transform 1 0 36340 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 25201
transform 1 0 37444 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 25201
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1636993656
transform 1 0 38180 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1636993656
transform 1 0 39284 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1636993656
transform 1 0 40388 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1636993656
transform 1 0 41492 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 25201
transform 1 0 42596 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 25201
transform 1 0 43148 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1636993656
transform 1 0 43332 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1636993656
transform 1 0 44436 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1636993656
transform 1 0 45540 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1636993656
transform 1 0 46644 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 25201
transform 1 0 47748 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 25201
transform 1 0 48300 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1636993656
transform 1 0 48484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1636993656
transform 1 0 49588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1636993656
transform 1 0 50692 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1636993656
transform 1 0 51796 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 25201
transform 1 0 52900 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 25201
transform 1 0 53452 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1636993656
transform 1 0 53636 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1636993656
transform 1 0 54740 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1636993656
transform 1 0 55844 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1636993656
transform 1 0 56948 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 25201
transform 1 0 58052 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 25201
transform 1 0 58604 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_617
timestamp 1636993656
transform 1 0 58788 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_629
timestamp 1636993656
transform 1 0 59892 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_641
timestamp 1636993656
transform 1 0 60996 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_653
timestamp 1636993656
transform 1 0 62100 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 25201
transform 1 0 63204 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 25201
transform 1 0 63756 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_673
timestamp 1636993656
transform 1 0 63940 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_685
timestamp 1636993656
transform 1 0 65044 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_697
timestamp 1636993656
transform 1 0 66148 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_709
timestamp 1636993656
transform 1 0 67252 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 25201
transform 1 0 68356 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 25201
transform 1 0 68908 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_729
timestamp 1636993656
transform 1 0 69092 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_741
timestamp 1636993656
transform 1 0 70196 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_753
timestamp 1636993656
transform 1 0 71300 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_765
timestamp 1636993656
transform 1 0 72404 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_777
timestamp 25201
transform 1 0 73508 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_783
timestamp 25201
transform 1 0 74060 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_785
timestamp 1636993656
transform 1 0 74244 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_797
timestamp 1636993656
transform 1 0 75348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_809
timestamp 1636993656
transform 1 0 76452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_821
timestamp 25201
transform 1 0 77556 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1636993656
transform 1 0 2300 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1636993656
transform 1 0 3404 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 25201
transform 1 0 4508 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636993656
transform 1 0 4692 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1636993656
transform 1 0 5796 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1636993656
transform 1 0 6900 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1636993656
transform 1 0 8004 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 25201
transform 1 0 9108 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 25201
transform 1 0 9660 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1636993656
transform 1 0 9844 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1636993656
transform 1 0 10948 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1636993656
transform 1 0 12052 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1636993656
transform 1 0 13156 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 25201
transform 1 0 14260 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 25201
transform 1 0 14812 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1636993656
transform 1 0 14996 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1636993656
transform 1 0 16100 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1636993656
transform 1 0 17204 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1636993656
transform 1 0 18308 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 25201
transform 1 0 19412 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 25201
transform 1 0 19964 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1636993656
transform 1 0 20148 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1636993656
transform 1 0 21252 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1636993656
transform 1 0 22356 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1636993656
transform 1 0 23460 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 25201
transform 1 0 24564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 25201
transform 1 0 25116 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1636993656
transform 1 0 25300 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1636993656
transform 1 0 26404 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1636993656
transform 1 0 27508 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1636993656
transform 1 0 28612 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 25201
transform 1 0 29716 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 25201
transform 1 0 30268 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1636993656
transform 1 0 30452 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1636993656
transform 1 0 31556 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1636993656
transform 1 0 32660 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1636993656
transform 1 0 33764 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 25201
transform 1 0 34868 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 25201
transform 1 0 35420 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1636993656
transform 1 0 35604 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1636993656
transform 1 0 36708 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1636993656
transform 1 0 37812 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1636993656
transform 1 0 38916 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 25201
transform 1 0 40020 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 25201
transform 1 0 40572 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1636993656
transform 1 0 40756 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1636993656
transform 1 0 41860 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1636993656
transform 1 0 42964 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1636993656
transform 1 0 44068 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 25201
transform 1 0 45172 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 25201
transform 1 0 45724 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1636993656
transform 1 0 45908 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1636993656
transform 1 0 47012 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1636993656
transform 1 0 48116 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1636993656
transform 1 0 49220 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 25201
transform 1 0 50324 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 25201
transform 1 0 50876 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1636993656
transform 1 0 51060 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1636993656
transform 1 0 52164 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1636993656
transform 1 0 53268 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1636993656
transform 1 0 54372 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 25201
transform 1 0 55476 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 25201
transform 1 0 56028 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1636993656
transform 1 0 56212 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1636993656
transform 1 0 57316 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1636993656
transform 1 0 58420 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_625
timestamp 1636993656
transform 1 0 59524 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 25201
transform 1 0 60628 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 25201
transform 1 0 61180 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_645
timestamp 1636993656
transform 1 0 61364 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_657
timestamp 1636993656
transform 1 0 62468 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_669
timestamp 1636993656
transform 1 0 63572 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_681
timestamp 1636993656
transform 1 0 64676 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 25201
transform 1 0 65780 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 25201
transform 1 0 66332 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_701
timestamp 1636993656
transform 1 0 66516 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_713
timestamp 1636993656
transform 1 0 67620 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_725
timestamp 1636993656
transform 1 0 68724 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_737
timestamp 1636993656
transform 1 0 69828 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_749
timestamp 25201
transform 1 0 70932 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_755
timestamp 25201
transform 1 0 71484 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_757
timestamp 1636993656
transform 1 0 71668 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_769
timestamp 1636993656
transform 1 0 72772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_781
timestamp 1636993656
transform 1 0 73876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_793
timestamp 1636993656
transform 1 0 74980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_805
timestamp 25201
transform 1 0 76084 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_811
timestamp 25201
transform 1 0 76636 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_813
timestamp 25201
transform 1 0 76820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_821
timestamp 25201
transform 1 0 77556 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636993656
transform 1 0 2300 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636993656
transform 1 0 3404 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1636993656
transform 1 0 4508 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1636993656
transform 1 0 5612 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 25201
transform 1 0 6716 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 25201
transform 1 0 7084 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1636993656
transform 1 0 7268 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1636993656
transform 1 0 8372 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1636993656
transform 1 0 9476 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1636993656
transform 1 0 10580 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 25201
transform 1 0 11684 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 25201
transform 1 0 12236 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1636993656
transform 1 0 12420 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1636993656
transform 1 0 13524 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1636993656
transform 1 0 14628 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1636993656
transform 1 0 15732 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 25201
transform 1 0 16836 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 25201
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1636993656
transform 1 0 17572 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1636993656
transform 1 0 18676 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1636993656
transform 1 0 19780 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1636993656
transform 1 0 20884 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 25201
transform 1 0 21988 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 25201
transform 1 0 22540 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1636993656
transform 1 0 22724 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1636993656
transform 1 0 23828 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1636993656
transform 1 0 24932 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1636993656
transform 1 0 26036 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 25201
transform 1 0 27140 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 25201
transform 1 0 27692 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1636993656
transform 1 0 27876 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1636993656
transform 1 0 28980 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1636993656
transform 1 0 30084 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1636993656
transform 1 0 31188 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 25201
transform 1 0 32292 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 25201
transform 1 0 32844 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1636993656
transform 1 0 33028 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1636993656
transform 1 0 34132 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1636993656
transform 1 0 35236 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1636993656
transform 1 0 36340 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 25201
transform 1 0 37444 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 25201
transform 1 0 37996 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1636993656
transform 1 0 38180 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1636993656
transform 1 0 39284 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1636993656
transform 1 0 40388 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1636993656
transform 1 0 41492 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 25201
transform 1 0 42596 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 25201
transform 1 0 43148 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1636993656
transform 1 0 43332 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1636993656
transform 1 0 44436 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1636993656
transform 1 0 45540 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1636993656
transform 1 0 46644 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 25201
transform 1 0 47748 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 25201
transform 1 0 48300 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1636993656
transform 1 0 48484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1636993656
transform 1 0 49588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1636993656
transform 1 0 50692 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1636993656
transform 1 0 51796 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 25201
transform 1 0 52900 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 25201
transform 1 0 53452 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1636993656
transform 1 0 53636 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1636993656
transform 1 0 54740 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1636993656
transform 1 0 55844 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1636993656
transform 1 0 56948 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 25201
transform 1 0 58052 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 25201
transform 1 0 58604 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_617
timestamp 1636993656
transform 1 0 58788 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_629
timestamp 1636993656
transform 1 0 59892 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_641
timestamp 1636993656
transform 1 0 60996 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_653
timestamp 1636993656
transform 1 0 62100 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 25201
transform 1 0 63204 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 25201
transform 1 0 63756 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_673
timestamp 1636993656
transform 1 0 63940 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_685
timestamp 1636993656
transform 1 0 65044 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_697
timestamp 1636993656
transform 1 0 66148 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_709
timestamp 1636993656
transform 1 0 67252 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 25201
transform 1 0 68356 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 25201
transform 1 0 68908 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_729
timestamp 1636993656
transform 1 0 69092 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_741
timestamp 1636993656
transform 1 0 70196 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_753
timestamp 1636993656
transform 1 0 71300 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_765
timestamp 1636993656
transform 1 0 72404 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_777
timestamp 25201
transform 1 0 73508 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_783
timestamp 25201
transform 1 0 74060 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_785
timestamp 1636993656
transform 1 0 74244 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_797
timestamp 1636993656
transform 1 0 75348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_809
timestamp 1636993656
transform 1 0 76452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_821
timestamp 25201
transform 1 0 77556 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636993656
transform 1 0 2300 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636993656
transform 1 0 3404 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 25201
transform 1 0 4508 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636993656
transform 1 0 4692 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1636993656
transform 1 0 5796 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1636993656
transform 1 0 6900 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1636993656
transform 1 0 8004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 25201
transform 1 0 9108 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 25201
transform 1 0 9660 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1636993656
transform 1 0 9844 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1636993656
transform 1 0 10948 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1636993656
transform 1 0 12052 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1636993656
transform 1 0 13156 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 25201
transform 1 0 14260 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 25201
transform 1 0 14812 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1636993656
transform 1 0 14996 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1636993656
transform 1 0 16100 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1636993656
transform 1 0 17204 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1636993656
transform 1 0 18308 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 25201
transform 1 0 19412 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 25201
transform 1 0 19964 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1636993656
transform 1 0 20148 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1636993656
transform 1 0 21252 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1636993656
transform 1 0 22356 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1636993656
transform 1 0 23460 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 25201
transform 1 0 24564 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 25201
transform 1 0 25116 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1636993656
transform 1 0 25300 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1636993656
transform 1 0 26404 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1636993656
transform 1 0 27508 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1636993656
transform 1 0 28612 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 25201
transform 1 0 29716 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 25201
transform 1 0 30268 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1636993656
transform 1 0 30452 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1636993656
transform 1 0 31556 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1636993656
transform 1 0 32660 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1636993656
transform 1 0 33764 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 25201
transform 1 0 34868 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 25201
transform 1 0 35420 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1636993656
transform 1 0 35604 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1636993656
transform 1 0 36708 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1636993656
transform 1 0 37812 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1636993656
transform 1 0 38916 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 25201
transform 1 0 40020 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 25201
transform 1 0 40572 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1636993656
transform 1 0 40756 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1636993656
transform 1 0 41860 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1636993656
transform 1 0 42964 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1636993656
transform 1 0 44068 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 25201
transform 1 0 45172 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 25201
transform 1 0 45724 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1636993656
transform 1 0 45908 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1636993656
transform 1 0 47012 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1636993656
transform 1 0 48116 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1636993656
transform 1 0 49220 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 25201
transform 1 0 50324 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 25201
transform 1 0 50876 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1636993656
transform 1 0 51060 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1636993656
transform 1 0 52164 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1636993656
transform 1 0 53268 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1636993656
transform 1 0 54372 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 25201
transform 1 0 55476 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 25201
transform 1 0 56028 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1636993656
transform 1 0 56212 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1636993656
transform 1 0 57316 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1636993656
transform 1 0 58420 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_625
timestamp 1636993656
transform 1 0 59524 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 25201
transform 1 0 60628 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 25201
transform 1 0 61180 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_645
timestamp 1636993656
transform 1 0 61364 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_657
timestamp 1636993656
transform 1 0 62468 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_669
timestamp 1636993656
transform 1 0 63572 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_681
timestamp 1636993656
transform 1 0 64676 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 25201
transform 1 0 65780 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 25201
transform 1 0 66332 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_701
timestamp 1636993656
transform 1 0 66516 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_713
timestamp 1636993656
transform 1 0 67620 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_725
timestamp 1636993656
transform 1 0 68724 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_737
timestamp 1636993656
transform 1 0 69828 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_749
timestamp 25201
transform 1 0 70932 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_755
timestamp 25201
transform 1 0 71484 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_757
timestamp 1636993656
transform 1 0 71668 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_769
timestamp 1636993656
transform 1 0 72772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_781
timestamp 1636993656
transform 1 0 73876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_793
timestamp 1636993656
transform 1 0 74980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_805
timestamp 25201
transform 1 0 76084 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_811
timestamp 25201
transform 1 0 76636 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_813
timestamp 25201
transform 1 0 76820 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_821
timestamp 25201
transform 1 0 77556 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636993656
transform 1 0 2300 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636993656
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636993656
transform 1 0 4508 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1636993656
transform 1 0 5612 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 25201
transform 1 0 6716 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 25201
transform 1 0 7084 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1636993656
transform 1 0 7268 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1636993656
transform 1 0 8372 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1636993656
transform 1 0 9476 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1636993656
transform 1 0 10580 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 25201
transform 1 0 11684 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 25201
transform 1 0 12236 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1636993656
transform 1 0 12420 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1636993656
transform 1 0 13524 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1636993656
transform 1 0 14628 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1636993656
transform 1 0 15732 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 25201
transform 1 0 16836 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 25201
transform 1 0 17388 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1636993656
transform 1 0 17572 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1636993656
transform 1 0 18676 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1636993656
transform 1 0 19780 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1636993656
transform 1 0 20884 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 25201
transform 1 0 21988 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 25201
transform 1 0 22540 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1636993656
transform 1 0 22724 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1636993656
transform 1 0 23828 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1636993656
transform 1 0 24932 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1636993656
transform 1 0 26036 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 25201
transform 1 0 27140 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 25201
transform 1 0 27692 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1636993656
transform 1 0 27876 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1636993656
transform 1 0 28980 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1636993656
transform 1 0 30084 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1636993656
transform 1 0 31188 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 25201
transform 1 0 32292 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 25201
transform 1 0 32844 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1636993656
transform 1 0 33028 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1636993656
transform 1 0 34132 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1636993656
transform 1 0 35236 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1636993656
transform 1 0 36340 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 25201
transform 1 0 37444 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 25201
transform 1 0 37996 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1636993656
transform 1 0 38180 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1636993656
transform 1 0 39284 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1636993656
transform 1 0 40388 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1636993656
transform 1 0 41492 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 25201
transform 1 0 42596 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 25201
transform 1 0 43148 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1636993656
transform 1 0 43332 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1636993656
transform 1 0 44436 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1636993656
transform 1 0 45540 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1636993656
transform 1 0 46644 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 25201
transform 1 0 47748 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 25201
transform 1 0 48300 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1636993656
transform 1 0 48484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1636993656
transform 1 0 49588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1636993656
transform 1 0 50692 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1636993656
transform 1 0 51796 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 25201
transform 1 0 52900 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 25201
transform 1 0 53452 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1636993656
transform 1 0 53636 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1636993656
transform 1 0 54740 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1636993656
transform 1 0 55844 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1636993656
transform 1 0 56948 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 25201
transform 1 0 58052 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 25201
transform 1 0 58604 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_617
timestamp 1636993656
transform 1 0 58788 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_629
timestamp 1636993656
transform 1 0 59892 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_641
timestamp 1636993656
transform 1 0 60996 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_653
timestamp 1636993656
transform 1 0 62100 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 25201
transform 1 0 63204 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 25201
transform 1 0 63756 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_673
timestamp 1636993656
transform 1 0 63940 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_685
timestamp 1636993656
transform 1 0 65044 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_697
timestamp 1636993656
transform 1 0 66148 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_709
timestamp 1636993656
transform 1 0 67252 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 25201
transform 1 0 68356 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 25201
transform 1 0 68908 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_729
timestamp 1636993656
transform 1 0 69092 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_741
timestamp 1636993656
transform 1 0 70196 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_753
timestamp 1636993656
transform 1 0 71300 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_765
timestamp 1636993656
transform 1 0 72404 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_777
timestamp 25201
transform 1 0 73508 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_783
timestamp 25201
transform 1 0 74060 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_785
timestamp 1636993656
transform 1 0 74244 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_797
timestamp 1636993656
transform 1 0 75348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_809
timestamp 1636993656
transform 1 0 76452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_821
timestamp 25201
transform 1 0 77556 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636993656
transform 1 0 2300 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636993656
transform 1 0 3404 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 25201
transform 1 0 4508 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1636993656
transform 1 0 4692 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1636993656
transform 1 0 5796 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1636993656
transform 1 0 6900 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1636993656
transform 1 0 8004 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 25201
transform 1 0 9108 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 25201
transform 1 0 9660 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1636993656
transform 1 0 9844 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1636993656
transform 1 0 10948 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1636993656
transform 1 0 12052 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1636993656
transform 1 0 13156 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 25201
transform 1 0 14260 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 25201
transform 1 0 14812 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1636993656
transform 1 0 14996 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1636993656
transform 1 0 16100 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1636993656
transform 1 0 17204 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1636993656
transform 1 0 18308 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 25201
transform 1 0 19412 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 25201
transform 1 0 19964 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1636993656
transform 1 0 20148 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1636993656
transform 1 0 21252 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1636993656
transform 1 0 22356 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1636993656
transform 1 0 23460 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 25201
transform 1 0 24564 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 25201
transform 1 0 25116 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1636993656
transform 1 0 25300 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1636993656
transform 1 0 26404 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1636993656
transform 1 0 27508 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1636993656
transform 1 0 28612 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 25201
transform 1 0 29716 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 25201
transform 1 0 30268 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1636993656
transform 1 0 30452 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1636993656
transform 1 0 31556 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1636993656
transform 1 0 32660 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1636993656
transform 1 0 33764 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 25201
transform 1 0 34868 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 25201
transform 1 0 35420 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1636993656
transform 1 0 35604 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1636993656
transform 1 0 36708 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1636993656
transform 1 0 37812 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1636993656
transform 1 0 38916 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 25201
transform 1 0 40020 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 25201
transform 1 0 40572 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1636993656
transform 1 0 40756 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1636993656
transform 1 0 41860 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1636993656
transform 1 0 42964 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1636993656
transform 1 0 44068 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 25201
transform 1 0 45172 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 25201
transform 1 0 45724 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1636993656
transform 1 0 45908 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1636993656
transform 1 0 47012 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1636993656
transform 1 0 48116 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1636993656
transform 1 0 49220 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 25201
transform 1 0 50324 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 25201
transform 1 0 50876 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1636993656
transform 1 0 51060 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1636993656
transform 1 0 52164 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1636993656
transform 1 0 53268 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1636993656
transform 1 0 54372 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 25201
transform 1 0 55476 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 25201
transform 1 0 56028 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1636993656
transform 1 0 56212 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1636993656
transform 1 0 57316 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1636993656
transform 1 0 58420 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_625
timestamp 1636993656
transform 1 0 59524 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 25201
transform 1 0 60628 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 25201
transform 1 0 61180 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_645
timestamp 1636993656
transform 1 0 61364 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_657
timestamp 1636993656
transform 1 0 62468 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_669
timestamp 1636993656
transform 1 0 63572 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_681
timestamp 1636993656
transform 1 0 64676 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 25201
transform 1 0 65780 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 25201
transform 1 0 66332 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_701
timestamp 1636993656
transform 1 0 66516 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_713
timestamp 1636993656
transform 1 0 67620 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_725
timestamp 1636993656
transform 1 0 68724 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_737
timestamp 1636993656
transform 1 0 69828 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_749
timestamp 25201
transform 1 0 70932 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_755
timestamp 25201
transform 1 0 71484 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_757
timestamp 1636993656
transform 1 0 71668 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_769
timestamp 1636993656
transform 1 0 72772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_781
timestamp 1636993656
transform 1 0 73876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_793
timestamp 1636993656
transform 1 0 74980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_805
timestamp 25201
transform 1 0 76084 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_811
timestamp 25201
transform 1 0 76636 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_813
timestamp 25201
transform 1 0 76820 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_821
timestamp 25201
transform 1 0 77556 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1636993656
transform 1 0 2300 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1636993656
transform 1 0 3404 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1636993656
transform 1 0 4508 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1636993656
transform 1 0 5612 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 25201
transform 1 0 6716 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 25201
transform 1 0 7084 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1636993656
transform 1 0 7268 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1636993656
transform 1 0 8372 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1636993656
transform 1 0 9476 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1636993656
transform 1 0 10580 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 25201
transform 1 0 11684 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 25201
transform 1 0 12236 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1636993656
transform 1 0 12420 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1636993656
transform 1 0 13524 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1636993656
transform 1 0 14628 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1636993656
transform 1 0 15732 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 25201
transform 1 0 16836 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 25201
transform 1 0 17388 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1636993656
transform 1 0 17572 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1636993656
transform 1 0 18676 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1636993656
transform 1 0 19780 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1636993656
transform 1 0 20884 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 25201
transform 1 0 21988 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 25201
transform 1 0 22540 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1636993656
transform 1 0 22724 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1636993656
transform 1 0 23828 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1636993656
transform 1 0 24932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1636993656
transform 1 0 26036 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 25201
transform 1 0 27140 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 25201
transform 1 0 27692 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1636993656
transform 1 0 27876 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1636993656
transform 1 0 28980 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1636993656
transform 1 0 30084 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1636993656
transform 1 0 31188 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 25201
transform 1 0 32292 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 25201
transform 1 0 32844 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1636993656
transform 1 0 33028 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1636993656
transform 1 0 34132 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1636993656
transform 1 0 35236 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1636993656
transform 1 0 36340 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 25201
transform 1 0 37444 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 25201
transform 1 0 37996 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1636993656
transform 1 0 38180 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1636993656
transform 1 0 39284 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1636993656
transform 1 0 40388 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1636993656
transform 1 0 41492 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 25201
transform 1 0 42596 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 25201
transform 1 0 43148 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1636993656
transform 1 0 43332 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1636993656
transform 1 0 44436 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1636993656
transform 1 0 45540 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1636993656
transform 1 0 46644 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 25201
transform 1 0 47748 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 25201
transform 1 0 48300 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1636993656
transform 1 0 48484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1636993656
transform 1 0 49588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1636993656
transform 1 0 50692 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1636993656
transform 1 0 51796 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 25201
transform 1 0 52900 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 25201
transform 1 0 53452 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1636993656
transform 1 0 53636 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1636993656
transform 1 0 54740 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1636993656
transform 1 0 55844 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1636993656
transform 1 0 56948 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 25201
transform 1 0 58052 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 25201
transform 1 0 58604 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_617
timestamp 1636993656
transform 1 0 58788 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_629
timestamp 1636993656
transform 1 0 59892 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_641
timestamp 1636993656
transform 1 0 60996 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_653
timestamp 1636993656
transform 1 0 62100 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 25201
transform 1 0 63204 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 25201
transform 1 0 63756 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_673
timestamp 1636993656
transform 1 0 63940 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_685
timestamp 1636993656
transform 1 0 65044 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_697
timestamp 1636993656
transform 1 0 66148 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_709
timestamp 1636993656
transform 1 0 67252 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_721
timestamp 25201
transform 1 0 68356 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_727
timestamp 25201
transform 1 0 68908 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_729
timestamp 1636993656
transform 1 0 69092 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_741
timestamp 1636993656
transform 1 0 70196 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_753
timestamp 1636993656
transform 1 0 71300 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_765
timestamp 1636993656
transform 1 0 72404 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_777
timestamp 25201
transform 1 0 73508 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_783
timestamp 25201
transform 1 0 74060 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_785
timestamp 1636993656
transform 1 0 74244 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_797
timestamp 1636993656
transform 1 0 75348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_809
timestamp 1636993656
transform 1 0 76452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_821
timestamp 25201
transform 1 0 77556 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636993656
transform 1 0 2300 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636993656
transform 1 0 3404 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 25201
transform 1 0 4508 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636993656
transform 1 0 4692 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1636993656
transform 1 0 5796 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1636993656
transform 1 0 6900 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1636993656
transform 1 0 8004 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 25201
transform 1 0 9108 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 25201
transform 1 0 9660 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1636993656
transform 1 0 9844 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1636993656
transform 1 0 10948 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1636993656
transform 1 0 12052 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1636993656
transform 1 0 13156 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 25201
transform 1 0 14260 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 25201
transform 1 0 14812 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1636993656
transform 1 0 14996 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1636993656
transform 1 0 16100 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1636993656
transform 1 0 17204 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1636993656
transform 1 0 18308 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 25201
transform 1 0 19412 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 25201
transform 1 0 19964 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1636993656
transform 1 0 20148 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1636993656
transform 1 0 21252 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1636993656
transform 1 0 22356 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1636993656
transform 1 0 23460 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 25201
transform 1 0 24564 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 25201
transform 1 0 25116 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1636993656
transform 1 0 25300 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1636993656
transform 1 0 26404 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1636993656
transform 1 0 27508 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1636993656
transform 1 0 28612 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 25201
transform 1 0 29716 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 25201
transform 1 0 30268 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1636993656
transform 1 0 30452 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1636993656
transform 1 0 31556 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1636993656
transform 1 0 32660 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1636993656
transform 1 0 33764 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 25201
transform 1 0 34868 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 25201
transform 1 0 35420 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1636993656
transform 1 0 35604 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1636993656
transform 1 0 36708 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1636993656
transform 1 0 37812 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1636993656
transform 1 0 38916 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 25201
transform 1 0 40020 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 25201
transform 1 0 40572 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1636993656
transform 1 0 40756 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1636993656
transform 1 0 41860 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1636993656
transform 1 0 42964 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1636993656
transform 1 0 44068 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 25201
transform 1 0 45172 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 25201
transform 1 0 45724 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1636993656
transform 1 0 45908 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1636993656
transform 1 0 47012 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1636993656
transform 1 0 48116 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1636993656
transform 1 0 49220 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 25201
transform 1 0 50324 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 25201
transform 1 0 50876 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1636993656
transform 1 0 51060 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1636993656
transform 1 0 52164 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1636993656
transform 1 0 53268 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1636993656
transform 1 0 54372 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 25201
transform 1 0 55476 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 25201
transform 1 0 56028 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1636993656
transform 1 0 56212 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1636993656
transform 1 0 57316 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1636993656
transform 1 0 58420 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_625
timestamp 1636993656
transform 1 0 59524 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 25201
transform 1 0 60628 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 25201
transform 1 0 61180 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_645
timestamp 1636993656
transform 1 0 61364 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_657
timestamp 1636993656
transform 1 0 62468 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_669
timestamp 1636993656
transform 1 0 63572 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_681
timestamp 1636993656
transform 1 0 64676 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 25201
transform 1 0 65780 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 25201
transform 1 0 66332 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_701
timestamp 1636993656
transform 1 0 66516 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_713
timestamp 1636993656
transform 1 0 67620 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_725
timestamp 1636993656
transform 1 0 68724 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_737
timestamp 1636993656
transform 1 0 69828 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_749
timestamp 25201
transform 1 0 70932 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_755
timestamp 25201
transform 1 0 71484 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_757
timestamp 1636993656
transform 1 0 71668 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_769
timestamp 1636993656
transform 1 0 72772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_781
timestamp 1636993656
transform 1 0 73876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_793
timestamp 1636993656
transform 1 0 74980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_805
timestamp 25201
transform 1 0 76084 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_811
timestamp 25201
transform 1 0 76636 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_813
timestamp 25201
transform 1 0 76820 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_821
timestamp 25201
transform 1 0 77556 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1636993656
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1636993656
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1636993656
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1636993656
transform 1 0 5612 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 25201
transform 1 0 6716 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 25201
transform 1 0 7084 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1636993656
transform 1 0 7268 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1636993656
transform 1 0 8372 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1636993656
transform 1 0 9476 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1636993656
transform 1 0 10580 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 25201
transform 1 0 11684 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 25201
transform 1 0 12236 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1636993656
transform 1 0 12420 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1636993656
transform 1 0 13524 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1636993656
transform 1 0 14628 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1636993656
transform 1 0 15732 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 25201
transform 1 0 16836 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 25201
transform 1 0 17388 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1636993656
transform 1 0 17572 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1636993656
transform 1 0 18676 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1636993656
transform 1 0 19780 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1636993656
transform 1 0 20884 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 25201
transform 1 0 21988 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 25201
transform 1 0 22540 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1636993656
transform 1 0 22724 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1636993656
transform 1 0 23828 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1636993656
transform 1 0 24932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1636993656
transform 1 0 26036 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 25201
transform 1 0 27140 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 25201
transform 1 0 27692 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1636993656
transform 1 0 27876 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1636993656
transform 1 0 28980 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1636993656
transform 1 0 30084 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1636993656
transform 1 0 31188 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 25201
transform 1 0 32292 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 25201
transform 1 0 32844 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1636993656
transform 1 0 33028 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1636993656
transform 1 0 34132 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1636993656
transform 1 0 35236 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1636993656
transform 1 0 36340 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 25201
transform 1 0 37444 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 25201
transform 1 0 37996 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1636993656
transform 1 0 38180 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1636993656
transform 1 0 39284 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1636993656
transform 1 0 40388 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1636993656
transform 1 0 41492 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 25201
transform 1 0 42596 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 25201
transform 1 0 43148 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1636993656
transform 1 0 43332 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1636993656
transform 1 0 44436 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1636993656
transform 1 0 45540 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1636993656
transform 1 0 46644 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 25201
transform 1 0 47748 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 25201
transform 1 0 48300 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1636993656
transform 1 0 48484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1636993656
transform 1 0 49588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1636993656
transform 1 0 50692 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1636993656
transform 1 0 51796 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 25201
transform 1 0 52900 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 25201
transform 1 0 53452 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1636993656
transform 1 0 53636 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1636993656
transform 1 0 54740 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1636993656
transform 1 0 55844 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1636993656
transform 1 0 56948 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 25201
transform 1 0 58052 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 25201
transform 1 0 58604 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_617
timestamp 1636993656
transform 1 0 58788 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_629
timestamp 1636993656
transform 1 0 59892 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_641
timestamp 1636993656
transform 1 0 60996 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_653
timestamp 1636993656
transform 1 0 62100 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 25201
transform 1 0 63204 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 25201
transform 1 0 63756 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_673
timestamp 1636993656
transform 1 0 63940 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_685
timestamp 1636993656
transform 1 0 65044 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_697
timestamp 1636993656
transform 1 0 66148 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_709
timestamp 1636993656
transform 1 0 67252 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 25201
transform 1 0 68356 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 25201
transform 1 0 68908 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_729
timestamp 1636993656
transform 1 0 69092 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_741
timestamp 1636993656
transform 1 0 70196 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_753
timestamp 1636993656
transform 1 0 71300 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_765
timestamp 1636993656
transform 1 0 72404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_777
timestamp 25201
transform 1 0 73508 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_783
timestamp 25201
transform 1 0 74060 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_785
timestamp 1636993656
transform 1 0 74244 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_797
timestamp 1636993656
transform 1 0 75348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_809
timestamp 1636993656
transform 1 0 76452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_821
timestamp 25201
transform 1 0 77556 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636993656
transform 1 0 2300 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636993656
transform 1 0 3404 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 25201
transform 1 0 4508 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636993656
transform 1 0 4692 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1636993656
transform 1 0 5796 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1636993656
transform 1 0 6900 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1636993656
transform 1 0 8004 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 25201
transform 1 0 9108 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 25201
transform 1 0 9660 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1636993656
transform 1 0 9844 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1636993656
transform 1 0 10948 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1636993656
transform 1 0 12052 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1636993656
transform 1 0 13156 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 25201
transform 1 0 14260 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 25201
transform 1 0 14812 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1636993656
transform 1 0 14996 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1636993656
transform 1 0 16100 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1636993656
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1636993656
transform 1 0 18308 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 25201
transform 1 0 19412 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 25201
transform 1 0 19964 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1636993656
transform 1 0 20148 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1636993656
transform 1 0 21252 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1636993656
transform 1 0 22356 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1636993656
transform 1 0 23460 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 25201
transform 1 0 24564 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 25201
transform 1 0 25116 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1636993656
transform 1 0 25300 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1636993656
transform 1 0 26404 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1636993656
transform 1 0 27508 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1636993656
transform 1 0 28612 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 25201
transform 1 0 29716 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 25201
transform 1 0 30268 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1636993656
transform 1 0 30452 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1636993656
transform 1 0 31556 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1636993656
transform 1 0 32660 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1636993656
transform 1 0 33764 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 25201
transform 1 0 34868 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 25201
transform 1 0 35420 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1636993656
transform 1 0 35604 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1636993656
transform 1 0 36708 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1636993656
transform 1 0 37812 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1636993656
transform 1 0 38916 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 25201
transform 1 0 40020 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 25201
transform 1 0 40572 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1636993656
transform 1 0 40756 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1636993656
transform 1 0 41860 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1636993656
transform 1 0 42964 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1636993656
transform 1 0 44068 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 25201
transform 1 0 45172 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 25201
transform 1 0 45724 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1636993656
transform 1 0 45908 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1636993656
transform 1 0 47012 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1636993656
transform 1 0 48116 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1636993656
transform 1 0 49220 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 25201
transform 1 0 50324 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 25201
transform 1 0 50876 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1636993656
transform 1 0 51060 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1636993656
transform 1 0 52164 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1636993656
transform 1 0 53268 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1636993656
transform 1 0 54372 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 25201
transform 1 0 55476 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 25201
transform 1 0 56028 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1636993656
transform 1 0 56212 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1636993656
transform 1 0 57316 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1636993656
transform 1 0 58420 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_625
timestamp 1636993656
transform 1 0 59524 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 25201
transform 1 0 60628 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 25201
transform 1 0 61180 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_645
timestamp 1636993656
transform 1 0 61364 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_657
timestamp 1636993656
transform 1 0 62468 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_669
timestamp 1636993656
transform 1 0 63572 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_681
timestamp 1636993656
transform 1 0 64676 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 25201
transform 1 0 65780 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 25201
transform 1 0 66332 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_701
timestamp 1636993656
transform 1 0 66516 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_713
timestamp 1636993656
transform 1 0 67620 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_725
timestamp 1636993656
transform 1 0 68724 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_737
timestamp 1636993656
transform 1 0 69828 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_749
timestamp 25201
transform 1 0 70932 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_755
timestamp 25201
transform 1 0 71484 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_757
timestamp 1636993656
transform 1 0 71668 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_769
timestamp 1636993656
transform 1 0 72772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_781
timestamp 1636993656
transform 1 0 73876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_793
timestamp 1636993656
transform 1 0 74980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_805
timestamp 25201
transform 1 0 76084 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_811
timestamp 25201
transform 1 0 76636 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_813
timestamp 25201
transform 1 0 76820 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_821
timestamp 25201
transform 1 0 77556 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636993656
transform 1 0 2300 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636993656
transform 1 0 3404 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1636993656
transform 1 0 4508 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1636993656
transform 1 0 5612 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 25201
transform 1 0 6716 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 25201
transform 1 0 7084 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1636993656
transform 1 0 7268 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1636993656
transform 1 0 8372 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1636993656
transform 1 0 9476 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1636993656
transform 1 0 10580 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 25201
transform 1 0 11684 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 25201
transform 1 0 12236 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1636993656
transform 1 0 12420 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1636993656
transform 1 0 13524 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1636993656
transform 1 0 14628 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1636993656
transform 1 0 15732 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 25201
transform 1 0 16836 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 25201
transform 1 0 17388 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1636993656
transform 1 0 17572 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1636993656
transform 1 0 18676 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1636993656
transform 1 0 19780 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1636993656
transform 1 0 20884 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 25201
transform 1 0 21988 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 25201
transform 1 0 22540 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1636993656
transform 1 0 22724 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1636993656
transform 1 0 23828 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1636993656
transform 1 0 24932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1636993656
transform 1 0 26036 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 25201
transform 1 0 27140 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 25201
transform 1 0 27692 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1636993656
transform 1 0 27876 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1636993656
transform 1 0 28980 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1636993656
transform 1 0 30084 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1636993656
transform 1 0 31188 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 25201
transform 1 0 32292 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 25201
transform 1 0 32844 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1636993656
transform 1 0 33028 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1636993656
transform 1 0 34132 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1636993656
transform 1 0 35236 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1636993656
transform 1 0 36340 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 25201
transform 1 0 37444 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 25201
transform 1 0 37996 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1636993656
transform 1 0 38180 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1636993656
transform 1 0 39284 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1636993656
transform 1 0 40388 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1636993656
transform 1 0 41492 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 25201
transform 1 0 42596 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 25201
transform 1 0 43148 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1636993656
transform 1 0 43332 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1636993656
transform 1 0 44436 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1636993656
transform 1 0 45540 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1636993656
transform 1 0 46644 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 25201
transform 1 0 47748 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 25201
transform 1 0 48300 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1636993656
transform 1 0 48484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1636993656
transform 1 0 49588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1636993656
transform 1 0 50692 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1636993656
transform 1 0 51796 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 25201
transform 1 0 52900 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 25201
transform 1 0 53452 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1636993656
transform 1 0 53636 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1636993656
transform 1 0 54740 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1636993656
transform 1 0 55844 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1636993656
transform 1 0 56948 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 25201
transform 1 0 58052 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 25201
transform 1 0 58604 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_617
timestamp 1636993656
transform 1 0 58788 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_629
timestamp 1636993656
transform 1 0 59892 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_641
timestamp 1636993656
transform 1 0 60996 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_653
timestamp 1636993656
transform 1 0 62100 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 25201
transform 1 0 63204 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 25201
transform 1 0 63756 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_673
timestamp 1636993656
transform 1 0 63940 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_685
timestamp 1636993656
transform 1 0 65044 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_697
timestamp 1636993656
transform 1 0 66148 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_709
timestamp 1636993656
transform 1 0 67252 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 25201
transform 1 0 68356 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 25201
transform 1 0 68908 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_729
timestamp 1636993656
transform 1 0 69092 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_741
timestamp 1636993656
transform 1 0 70196 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_753
timestamp 1636993656
transform 1 0 71300 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_765
timestamp 1636993656
transform 1 0 72404 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_777
timestamp 25201
transform 1 0 73508 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_783
timestamp 25201
transform 1 0 74060 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_785
timestamp 1636993656
transform 1 0 74244 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_797
timestamp 1636993656
transform 1 0 75348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_809
timestamp 1636993656
transform 1 0 76452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_821
timestamp 25201
transform 1 0 77556 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1636993656
transform 1 0 2300 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1636993656
transform 1 0 3404 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 25201
transform 1 0 4508 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636993656
transform 1 0 4692 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1636993656
transform 1 0 5796 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1636993656
transform 1 0 6900 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1636993656
transform 1 0 8004 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 25201
transform 1 0 9108 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 25201
transform 1 0 9660 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1636993656
transform 1 0 9844 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1636993656
transform 1 0 10948 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1636993656
transform 1 0 12052 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1636993656
transform 1 0 13156 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 25201
transform 1 0 14260 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 25201
transform 1 0 14812 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1636993656
transform 1 0 14996 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1636993656
transform 1 0 16100 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1636993656
transform 1 0 17204 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1636993656
transform 1 0 18308 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 25201
transform 1 0 19412 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 25201
transform 1 0 19964 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1636993656
transform 1 0 20148 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1636993656
transform 1 0 21252 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1636993656
transform 1 0 22356 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1636993656
transform 1 0 23460 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 25201
transform 1 0 24564 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 25201
transform 1 0 25116 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1636993656
transform 1 0 25300 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1636993656
transform 1 0 26404 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1636993656
transform 1 0 27508 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1636993656
transform 1 0 28612 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 25201
transform 1 0 29716 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 25201
transform 1 0 30268 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1636993656
transform 1 0 30452 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1636993656
transform 1 0 31556 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1636993656
transform 1 0 32660 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1636993656
transform 1 0 33764 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 25201
transform 1 0 34868 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 25201
transform 1 0 35420 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1636993656
transform 1 0 35604 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1636993656
transform 1 0 36708 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1636993656
transform 1 0 37812 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1636993656
transform 1 0 38916 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 25201
transform 1 0 40020 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 25201
transform 1 0 40572 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1636993656
transform 1 0 40756 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1636993656
transform 1 0 41860 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1636993656
transform 1 0 42964 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1636993656
transform 1 0 44068 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 25201
transform 1 0 45172 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 25201
transform 1 0 45724 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1636993656
transform 1 0 45908 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1636993656
transform 1 0 47012 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1636993656
transform 1 0 48116 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1636993656
transform 1 0 49220 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 25201
transform 1 0 50324 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 25201
transform 1 0 50876 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1636993656
transform 1 0 51060 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1636993656
transform 1 0 52164 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1636993656
transform 1 0 53268 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1636993656
transform 1 0 54372 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 25201
transform 1 0 55476 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 25201
transform 1 0 56028 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1636993656
transform 1 0 56212 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1636993656
transform 1 0 57316 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1636993656
transform 1 0 58420 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_625
timestamp 1636993656
transform 1 0 59524 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 25201
transform 1 0 60628 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 25201
transform 1 0 61180 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_645
timestamp 1636993656
transform 1 0 61364 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_657
timestamp 1636993656
transform 1 0 62468 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_669
timestamp 1636993656
transform 1 0 63572 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_681
timestamp 1636993656
transform 1 0 64676 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 25201
transform 1 0 65780 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 25201
transform 1 0 66332 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_701
timestamp 1636993656
transform 1 0 66516 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_713
timestamp 1636993656
transform 1 0 67620 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_725
timestamp 1636993656
transform 1 0 68724 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_737
timestamp 1636993656
transform 1 0 69828 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_749
timestamp 25201
transform 1 0 70932 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_755
timestamp 25201
transform 1 0 71484 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_757
timestamp 1636993656
transform 1 0 71668 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_769
timestamp 1636993656
transform 1 0 72772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_781
timestamp 1636993656
transform 1 0 73876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_793
timestamp 1636993656
transform 1 0 74980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_805
timestamp 25201
transform 1 0 76084 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_811
timestamp 25201
transform 1 0 76636 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_813
timestamp 25201
transform 1 0 76820 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_821
timestamp 25201
transform 1 0 77556 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1636993656
transform 1 0 2300 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1636993656
transform 1 0 3404 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1636993656
transform 1 0 4508 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1636993656
transform 1 0 5612 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 25201
transform 1 0 6716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 25201
transform 1 0 7084 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1636993656
transform 1 0 7268 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1636993656
transform 1 0 8372 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1636993656
transform 1 0 9476 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1636993656
transform 1 0 10580 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 25201
transform 1 0 11684 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 25201
transform 1 0 12236 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1636993656
transform 1 0 12420 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1636993656
transform 1 0 13524 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1636993656
transform 1 0 14628 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1636993656
transform 1 0 15732 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 25201
transform 1 0 16836 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 25201
transform 1 0 17388 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1636993656
transform 1 0 17572 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1636993656
transform 1 0 18676 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1636993656
transform 1 0 19780 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1636993656
transform 1 0 20884 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 25201
transform 1 0 21988 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 25201
transform 1 0 22540 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1636993656
transform 1 0 22724 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1636993656
transform 1 0 23828 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1636993656
transform 1 0 24932 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1636993656
transform 1 0 26036 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 25201
transform 1 0 27140 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 25201
transform 1 0 27692 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1636993656
transform 1 0 27876 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1636993656
transform 1 0 28980 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1636993656
transform 1 0 30084 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1636993656
transform 1 0 31188 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 25201
transform 1 0 32292 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 25201
transform 1 0 32844 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1636993656
transform 1 0 33028 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1636993656
transform 1 0 34132 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1636993656
transform 1 0 35236 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1636993656
transform 1 0 36340 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 25201
transform 1 0 37444 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 25201
transform 1 0 37996 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1636993656
transform 1 0 38180 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1636993656
transform 1 0 39284 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1636993656
transform 1 0 40388 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1636993656
transform 1 0 41492 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 25201
transform 1 0 42596 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 25201
transform 1 0 43148 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1636993656
transform 1 0 43332 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1636993656
transform 1 0 44436 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1636993656
transform 1 0 45540 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1636993656
transform 1 0 46644 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 25201
transform 1 0 47748 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 25201
transform 1 0 48300 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1636993656
transform 1 0 48484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1636993656
transform 1 0 49588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1636993656
transform 1 0 50692 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1636993656
transform 1 0 51796 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 25201
transform 1 0 52900 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 25201
transform 1 0 53452 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1636993656
transform 1 0 53636 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1636993656
transform 1 0 54740 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1636993656
transform 1 0 55844 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1636993656
transform 1 0 56948 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 25201
transform 1 0 58052 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 25201
transform 1 0 58604 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_617
timestamp 1636993656
transform 1 0 58788 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_629
timestamp 1636993656
transform 1 0 59892 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_641
timestamp 1636993656
transform 1 0 60996 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_653
timestamp 1636993656
transform 1 0 62100 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 25201
transform 1 0 63204 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 25201
transform 1 0 63756 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_673
timestamp 1636993656
transform 1 0 63940 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_685
timestamp 1636993656
transform 1 0 65044 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_697
timestamp 1636993656
transform 1 0 66148 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_709
timestamp 1636993656
transform 1 0 67252 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 25201
transform 1 0 68356 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 25201
transform 1 0 68908 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_729
timestamp 1636993656
transform 1 0 69092 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_741
timestamp 1636993656
transform 1 0 70196 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_753
timestamp 1636993656
transform 1 0 71300 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_765
timestamp 1636993656
transform 1 0 72404 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_777
timestamp 25201
transform 1 0 73508 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_783
timestamp 25201
transform 1 0 74060 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_785
timestamp 1636993656
transform 1 0 74244 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_797
timestamp 1636993656
transform 1 0 75348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_809
timestamp 1636993656
transform 1 0 76452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_821
timestamp 25201
transform 1 0 77556 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636993656
transform 1 0 2300 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636993656
transform 1 0 3404 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 25201
transform 1 0 4508 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1636993656
transform 1 0 4692 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1636993656
transform 1 0 5796 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1636993656
transform 1 0 6900 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1636993656
transform 1 0 8004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 25201
transform 1 0 9108 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 25201
transform 1 0 9660 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1636993656
transform 1 0 9844 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1636993656
transform 1 0 10948 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1636993656
transform 1 0 12052 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1636993656
transform 1 0 13156 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 25201
transform 1 0 14260 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 25201
transform 1 0 14812 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1636993656
transform 1 0 14996 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1636993656
transform 1 0 16100 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1636993656
transform 1 0 17204 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1636993656
transform 1 0 18308 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 25201
transform 1 0 19412 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 25201
transform 1 0 19964 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1636993656
transform 1 0 20148 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1636993656
transform 1 0 21252 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1636993656
transform 1 0 22356 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1636993656
transform 1 0 23460 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 25201
transform 1 0 24564 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 25201
transform 1 0 25116 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1636993656
transform 1 0 25300 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1636993656
transform 1 0 26404 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1636993656
transform 1 0 27508 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1636993656
transform 1 0 28612 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 25201
transform 1 0 29716 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 25201
transform 1 0 30268 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1636993656
transform 1 0 30452 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1636993656
transform 1 0 31556 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1636993656
transform 1 0 32660 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1636993656
transform 1 0 33764 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 25201
transform 1 0 34868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 25201
transform 1 0 35420 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1636993656
transform 1 0 35604 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1636993656
transform 1 0 36708 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1636993656
transform 1 0 37812 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1636993656
transform 1 0 38916 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 25201
transform 1 0 40020 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 25201
transform 1 0 40572 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1636993656
transform 1 0 40756 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1636993656
transform 1 0 41860 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1636993656
transform 1 0 42964 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1636993656
transform 1 0 44068 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 25201
transform 1 0 45172 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 25201
transform 1 0 45724 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1636993656
transform 1 0 45908 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1636993656
transform 1 0 47012 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1636993656
transform 1 0 48116 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1636993656
transform 1 0 49220 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 25201
transform 1 0 50324 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 25201
transform 1 0 50876 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1636993656
transform 1 0 51060 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1636993656
transform 1 0 52164 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1636993656
transform 1 0 53268 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1636993656
transform 1 0 54372 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 25201
transform 1 0 55476 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 25201
transform 1 0 56028 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1636993656
transform 1 0 56212 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1636993656
transform 1 0 57316 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1636993656
transform 1 0 58420 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_625
timestamp 1636993656
transform 1 0 59524 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 25201
transform 1 0 60628 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 25201
transform 1 0 61180 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_645
timestamp 1636993656
transform 1 0 61364 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_657
timestamp 1636993656
transform 1 0 62468 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_669
timestamp 1636993656
transform 1 0 63572 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_681
timestamp 1636993656
transform 1 0 64676 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 25201
transform 1 0 65780 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 25201
transform 1 0 66332 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_701
timestamp 1636993656
transform 1 0 66516 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_713
timestamp 1636993656
transform 1 0 67620 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_725
timestamp 1636993656
transform 1 0 68724 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_737
timestamp 1636993656
transform 1 0 69828 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_749
timestamp 25201
transform 1 0 70932 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_755
timestamp 25201
transform 1 0 71484 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_757
timestamp 1636993656
transform 1 0 71668 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_769
timestamp 1636993656
transform 1 0 72772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_781
timestamp 1636993656
transform 1 0 73876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_793
timestamp 1636993656
transform 1 0 74980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_805
timestamp 25201
transform 1 0 76084 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_811
timestamp 25201
transform 1 0 76636 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_813
timestamp 25201
transform 1 0 76820 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_821
timestamp 25201
transform 1 0 77556 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636993656
transform 1 0 2300 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_15
timestamp 25201
transform 1 0 3404 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1636993656
transform 1 0 5612 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 25201
transform 1 0 6716 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 25201
transform 1 0 7084 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_57
timestamp 25201
transform 1 0 7268 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_63
timestamp 1636993656
transform 1 0 7820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_75
timestamp 25201
transform 1 0 8924 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_99
timestamp 25201
transform 1 0 11132 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 25201
transform 1 0 12144 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1636993656
transform 1 0 12420 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1636993656
transform 1 0 13524 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_137
timestamp 25201
transform 1 0 14628 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_143
timestamp 1636993656
transform 1 0 15180 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_155
timestamp 1636993656
transform 1 0 16284 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 25201
transform 1 0 17388 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_188
timestamp 1636993656
transform 1 0 19320 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_200
timestamp 1636993656
transform 1 0 20424 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_212
timestamp 25201
transform 1 0 21528 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 25201
transform 1 0 22540 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1636993656
transform 1 0 22724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_237
timestamp 25201
transform 1 0 23828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_259
timestamp 25201
transform 1 0 25852 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_263
timestamp 1636993656
transform 1 0 26220 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_275
timestamp 25201
transform 1 0 27324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 25201
transform 1 0 27692 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1636993656
transform 1 0 27876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_293
timestamp 25201
transform 1 0 28980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_299
timestamp 25201
transform 1 0 29532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_319
timestamp 1636993656
transform 1 0 31372 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_331
timestamp 25201
transform 1 0 32476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 25201
transform 1 0 32844 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 25201
transform 1 0 33028 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_348
timestamp 1636993656
transform 1 0 34040 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_360
timestamp 25201
transform 1 0 35144 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_379
timestamp 25201
transform 1 0 36892 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_383
timestamp 25201
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 25201
transform 1 0 37996 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1636993656
transform 1 0 38180 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1636993656
transform 1 0 39284 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_417
timestamp 25201
transform 1 0 40388 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_423
timestamp 1636993656
transform 1 0 40940 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_435
timestamp 1636993656
transform 1 0 42044 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 25201
transform 1 0 43148 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_449
timestamp 25201
transform 1 0 43332 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_457
timestamp 25201
transform 1 0 44068 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_479
timestamp 1636993656
transform 1 0 46092 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_491
timestamp 25201
transform 1 0 47196 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_499
timestamp 25201
transform 1 0 47932 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 25201
transform 1 0 48300 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1636993656
transform 1 0 48484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_517
timestamp 25201
transform 1 0 49588 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_539
timestamp 25201
transform 1 0 51612 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_543
timestamp 1636993656
transform 1 0 51980 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_555
timestamp 25201
transform 1 0 53084 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 25201
transform 1 0 53452 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1636993656
transform 1 0 53636 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_573
timestamp 25201
transform 1 0 54740 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_579
timestamp 25201
transform 1 0 55292 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_583
timestamp 1636993656
transform 1 0 55660 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_595
timestamp 1636993656
transform 1 0 56764 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_607
timestamp 25201
transform 1 0 57868 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_617
timestamp 25201
transform 1 0 58788 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_639
timestamp 1636993656
transform 1 0 60812 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_651
timestamp 1636993656
transform 1 0 61916 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_663
timestamp 25201
transform 1 0 63020 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 25201
transform 1 0 63756 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_673
timestamp 1636993656
transform 1 0 63940 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_685
timestamp 1636993656
transform 1 0 65044 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_697
timestamp 1636993656
transform 1 0 66148 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_709
timestamp 1636993656
transform 1 0 67252 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 25201
transform 1 0 68356 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 25201
transform 1 0 68908 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_729
timestamp 1636993656
transform 1 0 69092 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_741
timestamp 1636993656
transform 1 0 70196 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_753
timestamp 1636993656
transform 1 0 71300 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_765
timestamp 1636993656
transform 1 0 72404 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_777
timestamp 25201
transform 1 0 73508 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_783
timestamp 25201
transform 1 0 74060 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_785
timestamp 1636993656
transform 1 0 74244 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_797
timestamp 1636993656
transform 1 0 75348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_809
timestamp 1636993656
transform 1 0 76452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_821
timestamp 25201
transform 1 0 77556 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_19
timestamp 25201
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 25201
transform 1 0 4508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_29
timestamp 25201
transform 1 0 4692 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_37
timestamp 25201
transform 1 0 5428 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_57
timestamp 25201
transform 1 0 7268 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_79
timestamp 25201
transform 1 0 9292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 25201
transform 1 0 9660 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 25201
transform 1 0 9844 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_93
timestamp 25201
transform 1 0 10580 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_113
timestamp 25201
transform 1 0 12420 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_121
timestamp 25201
transform 1 0 13156 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 25201
transform 1 0 14812 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 25201
transform 1 0 14996 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_159
timestamp 25201
transform 1 0 16652 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 25201
transform 1 0 17388 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_169
timestamp 25201
transform 1 0 17572 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_177
timestamp 25201
transform 1 0 18308 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_197
timestamp 25201
transform 1 0 20148 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_219
timestamp 25201
transform 1 0 22172 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 25201
transform 1 0 22540 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_241
timestamp 25201
transform 1 0 24196 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 25201
transform 1 0 24932 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_253
timestamp 25201
transform 1 0 25300 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_261
timestamp 25201
transform 1 0 26036 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 25201
transform 1 0 27692 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 25201
transform 1 0 27876 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_299
timestamp 25201
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 25201
transform 1 0 30268 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 25201
transform 1 0 30452 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_317
timestamp 25201
transform 1 0 31188 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_337
timestamp 25201
transform 1 0 33028 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_359
timestamp 25201
transform 1 0 35052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 25201
transform 1 0 35420 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_365
timestamp 25201
transform 1 0 35604 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_373
timestamp 25201
transform 1 0 36340 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_393
timestamp 25201
transform 1 0 38180 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_401
timestamp 25201
transform 1 0 38916 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 25201
transform 1 0 40572 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_421
timestamp 25201
transform 1 0 40756 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_439
timestamp 25201
transform 1 0 42412 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_447
timestamp 25201
transform 1 0 43148 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_465
timestamp 25201
transform 1 0 44804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_473
timestamp 25201
transform 1 0 45540 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_477
timestamp 25201
transform 1 0 45908 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_499
timestamp 25201
transform 1 0 47932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_503
timestamp 25201
transform 1 0 48300 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_521
timestamp 25201
transform 1 0 49956 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_529
timestamp 25201
transform 1 0 50692 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_533
timestamp 25201
transform 1 0 51060 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_541
timestamp 25201
transform 1 0 51796 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_559
timestamp 25201
transform 1 0 53452 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_561
timestamp 25201
transform 1 0 53636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_579
timestamp 25201
transform 1 0 55292 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 25201
transform 1 0 56028 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_605
timestamp 25201
transform 1 0 57684 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_613
timestamp 25201
transform 1 0 58420 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_633
timestamp 25201
transform 1 0 60260 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_641
timestamp 25201
transform 1 0 60996 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_645
timestamp 1636993656
transform 1 0 61364 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_657
timestamp 1636993656
transform 1 0 62468 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_669
timestamp 25201
transform 1 0 63572 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_673
timestamp 1636993656
transform 1 0 63940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_685
timestamp 1636993656
transform 1 0 65044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_697
timestamp 25201
transform 1 0 66148 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_701
timestamp 1636993656
transform 1 0 66516 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_713
timestamp 1636993656
transform 1 0 67620 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_725
timestamp 25201
transform 1 0 68724 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_729
timestamp 1636993656
transform 1 0 69092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_741
timestamp 1636993656
transform 1 0 70196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_753
timestamp 25201
transform 1 0 71300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_757
timestamp 1636993656
transform 1 0 71668 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_769
timestamp 1636993656
transform 1 0 72772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_781
timestamp 25201
transform 1 0 73876 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_785
timestamp 1636993656
transform 1 0 74244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_797
timestamp 1636993656
transform 1 0 75348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_809
timestamp 25201
transform 1 0 76452 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_813
timestamp 25201
transform 1 0 76820 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_821
timestamp 25201
transform 1 0 77556 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 25201
transform -1 0 34960 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 25201
transform 1 0 21896 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 25201
transform -1 0 33580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 25201
transform 1 0 12696 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 25201
transform -1 0 12328 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 25201
transform 1 0 14168 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 25201
transform 1 0 24840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 25201
transform -1 0 36524 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 25201
transform 1 0 27048 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 25201
transform 1 0 3864 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 25201
transform 1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 25201
transform -1 0 18584 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 25201
transform -1 0 48116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 25201
transform 1 0 38456 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 25201
transform 1 0 41308 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 25201
transform -1 0 38916 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 25201
transform 1 0 30728 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 25201
transform 1 0 30728 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 25201
transform 1 0 48852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 25201
transform -1 0 48116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 25201
transform -1 0 45632 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 25201
transform -1 0 16652 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 25201
transform 1 0 7544 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 25201
transform 1 0 7912 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 25201
transform -1 0 29900 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 25201
transform -1 0 29624 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 25201
transform 1 0 29624 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 25201
transform -1 0 24104 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 25201
transform 1 0 12696 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 25201
transform 1 0 23644 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 25201
transform -1 0 28612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 25201
transform -1 0 28980 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 25201
transform -1 0 28152 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 25201
transform 1 0 29440 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 25201
transform 1 0 24472 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 25201
transform 1 0 31096 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 25201
transform -1 0 16008 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 25201
transform 1 0 7544 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 25201
transform 1 0 17112 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 25201
transform 1 0 47012 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 25201
transform -1 0 47380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 25201
transform -1 0 44436 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 25201
transform -1 0 41492 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 25201
transform 1 0 39560 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 25201
transform 1 0 34040 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 25201
transform -1 0 6624 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 25201
transform 1 0 11592 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 25201
transform 1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 25201
transform 1 0 5704 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 25201
transform 1 0 7728 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 25201
transform -1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 25201
transform 1 0 11224 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 25201
transform -1 0 17848 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 25201
transform -1 0 14168 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 25201
transform -1 0 26036 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 25201
transform 1 0 15088 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 25201
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 25201
transform -1 0 27048 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 25201
transform 1 0 25576 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 25201
transform 1 0 25944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 25201
transform -1 0 14168 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 25201
transform 1 0 16744 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 25201
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 25201
transform 1 0 42228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 25201
transform -1 0 40388 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 25201
transform 1 0 35604 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 25201
transform 1 0 16744 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 25201
transform 1 0 31832 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 25201
transform -1 0 33764 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 25201
transform -1 0 27784 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 25201
transform 1 0 31096 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 25201
transform 1 0 34776 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 25201
transform 1 0 21896 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 25201
transform 1 0 28704 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 25201
transform 1 0 28888 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 25201
transform 1 0 5704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 25201
transform 1 0 17480 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 25201
transform 1 0 23736 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 25201
transform 1 0 8464 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 25201
transform 1 0 13064 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 25201
transform -1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 25201
transform -1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 25201
transform 1 0 11592 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 25201
transform 1 0 21896 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 25201
transform 1 0 45908 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 25201
transform -1 0 44252 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 25201
transform 1 0 37352 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 25201
transform 1 0 15088 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 25201
transform 1 0 27416 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 25201
transform -1 0 28888 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 25201
transform 1 0 25208 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 25201
transform 1 0 48484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 25201
transform -1 0 43700 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 25201
transform -1 0 31096 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 25201
transform 1 0 29624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 25201
transform 1 0 21896 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 25201
transform 1 0 24472 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 25201
transform -1 0 29624 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 25201
transform 1 0 28152 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 25201
transform -1 0 51520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 25201
transform -1 0 43516 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 25201
transform -1 0 37352 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 25201
transform 1 0 37352 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 25201
transform -1 0 13432 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 25201
transform 1 0 11224 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 25201
transform -1 0 16376 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 25201
transform 1 0 17848 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 25201
transform -1 0 21988 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 25201
transform -1 0 16744 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 25201
transform -1 0 14904 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold111
timestamp 25201
transform -1 0 14904 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 25201
transform 1 0 38732 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 25201
transform 1 0 33672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 25201
transform 1 0 36616 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 25201
transform -1 0 36616 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 25201
transform -1 0 21528 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 25201
transform 1 0 14536 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 25201
transform -1 0 19320 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 25201
transform 1 0 35604 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold120
timestamp 25201
transform 1 0 45172 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 25201
transform -1 0 23736 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 25201
transform 1 0 16560 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 25201
transform -1 0 30360 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 25201
transform -1 0 32200 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold125
timestamp 25201
transform 1 0 31464 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 25201
transform -1 0 31648 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 25201
transform 1 0 22264 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold128
timestamp 25201
transform -1 0 30360 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 25201
transform 1 0 28888 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 25201
transform 1 0 24288 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold131
timestamp 25201
transform 1 0 28888 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 25201
transform -1 0 37352 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 25201
transform 1 0 38824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold134
timestamp 25201
transform 1 0 38548 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 25201
transform 1 0 27968 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 25201
transform 1 0 13432 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold137
timestamp 25201
transform -1 0 26956 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 25201
transform -1 0 36616 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 25201
transform 1 0 28152 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold140
timestamp 25201
transform 1 0 36616 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 25201
transform -1 0 23920 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 25201
transform -1 0 19688 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold143
timestamp 25201
transform -1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 25201
transform -1 0 34776 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 25201
transform -1 0 35052 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold146
timestamp 25201
transform -1 0 35512 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 25201
transform -1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 25201
transform 1 0 10856 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold149
timestamp 25201
transform 1 0 23368 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 25201
transform -1 0 42228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 25201
transform -1 0 42688 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold152
timestamp 25201
transform 1 0 43332 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 25201
transform -1 0 44988 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 25201
transform -1 0 41308 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold155
timestamp 25201
transform 1 0 39192 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 25201
transform -1 0 19872 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 25201
transform 1 0 18216 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold158
timestamp 25201
transform 1 0 20332 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 25201
transform 1 0 39376 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 25201
transform 1 0 44068 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold161
timestamp 25201
transform 1 0 46644 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 25201
transform 1 0 20608 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 25201
transform -1 0 16744 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold164
timestamp 25201
transform 1 0 18216 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 25201
transform 1 0 26312 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 25201
transform 1 0 69184 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold170
timestamp 25201
transform -1 0 76728 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 25201
transform -1 0 34040 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 25201
transform -1 0 58880 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 25201
transform -1 0 62836 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 25201
transform 1 0 74520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold177
timestamp 25201
transform -1 0 76728 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 25201
transform 1 0 6440 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 25201
transform 1 0 8280 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 25201
transform 1 0 19872 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 25201
transform -1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 25201
transform -1 0 29624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 25201
transform -1 0 68632 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 25201
transform 1 0 53728 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  hold187
timestamp 25201
transform 1 0 41492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 25201
transform 1 0 57408 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold189
timestamp 25201
transform 1 0 58788 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 25201
transform 1 0 25576 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 25201
transform -1 0 53176 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 25201
transform -1 0 73140 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 25201
transform 1 0 64768 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold197
timestamp 25201
transform 1 0 65504 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 25201
transform 1 0 8648 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 25201
transform 1 0 64400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 25201
transform -1 0 53912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold205
timestamp 25201
transform 1 0 52072 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 25201
transform 1 0 9016 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 25201
transform 1 0 54648 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold213
timestamp 25201
transform 1 0 54004 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 25201
transform -1 0 42596 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 25201
transform -1 0 69368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold221
timestamp 25201
transform 1 0 67528 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 25201
transform -1 0 42412 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 25201
transform 1 0 60996 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold229
timestamp 25201
transform 1 0 61732 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 25201
transform 1 0 9016 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 25201
transform -1 0 24380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 25201
transform 1 0 70104 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold238
timestamp 25201
transform 1 0 69460 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 25201
transform -1 0 42228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 25201
transform 1 0 71392 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold246
timestamp 25201
transform -1 0 73232 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 25201
transform -1 0 9752 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 25201
transform 1 0 11132 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  hold249
timestamp 25201
transform -1 0 10488 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 25201
transform 1 0 10120 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 25201
transform -1 0 45724 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 25201
transform -1 0 44068 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 25201
transform 1 0 48852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold259
timestamp 25201
transform -1 0 50048 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 25201
transform 1 0 31832 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 25201
transform -1 0 36800 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 25201
transform 1 0 23736 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 25201
transform 1 0 25944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 25201
transform 1 0 20424 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 25201
transform 1 0 18216 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 25201
transform 1 0 18216 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold267
timestamp 25201
transform 1 0 29624 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 25201
transform 1 0 23736 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 25201
transform -1 0 29624 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 25201
transform 1 0 30360 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 25201
transform 1 0 3128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 25201
transform 1 0 11960 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 25201
transform -1 0 13524 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 25201
transform 1 0 9016 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 25201
transform -1 0 11592 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 25201
transform 1 0 6624 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 25201
transform -1 0 26680 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 25201
transform 1 0 19320 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 25201
transform -1 0 19136 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 25201
transform -1 0 26220 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 25201
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 25201
transform -1 0 30360 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 25201
transform -1 0 30360 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 25201
transform 1 0 17296 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 25201
transform 1 0 28152 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 25201
transform 1 0 26680 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 25201
transform -1 0 28704 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 25201
transform -1 0 26680 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 25201
transform 1 0 16744 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 25201
transform 1 0 38180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold291
timestamp 25201
transform -1 0 35880 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 25201
transform -1 0 25208 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 25201
transform -1 0 22080 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold294
timestamp 25201
transform 1 0 15640 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 25201
transform 1 0 18952 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold296
timestamp 25201
transform -1 0 37352 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold297
timestamp 25201
transform -1 0 35144 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold298
timestamp 25201
transform -1 0 37536 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 25201
transform -1 0 37444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 25201
transform 1 0 33304 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold301
timestamp 25201
transform -1 0 31372 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold302
timestamp 25201
transform 1 0 34132 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold303
timestamp 25201
transform 1 0 33396 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 25201
transform -1 0 41952 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 25201
transform 1 0 40848 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold306
timestamp 25201
transform 1 0 36340 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold307
timestamp 25201
transform -1 0 43056 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold308
timestamp 25201
transform -1 0 25208 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold309
timestamp 25201
transform -1 0 18952 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 25201
transform 1 0 9752 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 25201
transform 1 0 19320 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold312
timestamp 25201
transform 1 0 39192 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold313
timestamp 25201
transform -1 0 39376 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 25201
transform -1 0 21896 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold315
timestamp 25201
transform -1 0 23736 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold316
timestamp 25201
transform 1 0 10120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold317
timestamp 25201
transform 1 0 6440 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 25201
transform 1 0 21160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold319
timestamp 25201
transform -1 0 27416 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold320
timestamp 25201
transform -1 0 34316 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold321
timestamp 25201
transform 1 0 22632 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 25201
transform -1 0 16008 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold325
timestamp 25201
transform -1 0 26956 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold326
timestamp 25201
transform -1 0 17112 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold327
timestamp 25201
transform 1 0 10120 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold330
timestamp 25201
transform 1 0 20792 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold331
timestamp 25201
transform -1 0 22264 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold332
timestamp 25201
transform -1 0 30636 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold333
timestamp 25201
transform 1 0 24472 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold336
timestamp 25201
transform -1 0 28888 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold337
timestamp 25201
transform -1 0 36616 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold338
timestamp 25201
transform 1 0 35052 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold339
timestamp 25201
transform 1 0 28888 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold342
timestamp 25201
transform -1 0 42780 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold343
timestamp 25201
transform 1 0 28152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold344
timestamp 25201
transform -1 0 38272 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold345
timestamp 25201
transform -1 0 38916 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold348
timestamp 25201
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold349
timestamp 25201
transform 1 0 3128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold350
timestamp 25201
transform -1 0 9936 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold351
timestamp 25201
transform 1 0 14536 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold354
timestamp 25201
transform 1 0 44068 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold355
timestamp 25201
transform -1 0 50692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold356
timestamp 25201
transform 1 0 45540 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold357
timestamp 25201
transform -1 0 45540 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold360
timestamp 25201
transform -1 0 17480 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold361
timestamp 25201
transform 1 0 4968 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold362
timestamp 25201
transform -1 0 19320 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold363
timestamp 25201
transform 1 0 11960 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s4s_1  hold366
timestamp 25201
transform -1 0 9200 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold367
timestamp 25201
transform 1 0 11960 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold368
timestamp 25201
transform -1 0 16008 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold369
timestamp 25201
transform -1 0 25392 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold372
timestamp 25201
transform 1 0 35880 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold373
timestamp 25201
transform -1 0 46644 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold374
timestamp 25201
transform -1 0 41860 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold375
timestamp 25201
transform -1 0 45540 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold378
timestamp 25201
transform 1 0 39928 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold379
timestamp 25201
transform 1 0 26312 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold380
timestamp 25201
transform 1 0 33304 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold381
timestamp 25201
transform -1 0 47104 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold384
timestamp 25201
transform 1 0 27048 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold385
timestamp 25201
transform 1 0 26680 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold386
timestamp 25201
transform 1 0 16744 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold387
timestamp 25201
transform 1 0 26312 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold390
timestamp 25201
transform -1 0 31464 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold391
timestamp 25201
transform -1 0 32384 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold392
timestamp 25201
transform -1 0 32936 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold393
timestamp 25201
transform -1 0 32752 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold396
timestamp 25201
transform 1 0 10856 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold397
timestamp 25201
transform 1 0 9384 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold398
timestamp 25201
transform -1 0 17480 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold399
timestamp 25201
transform -1 0 22540 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold402
timestamp 25201
transform -1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold403
timestamp 25201
transform 1 0 2392 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold404
timestamp 25201
transform 1 0 4968 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold405
timestamp 25201
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold408
timestamp 25201
transform 1 0 45908 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold409
timestamp 25201
transform -1 0 50784 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold410
timestamp 25201
transform -1 0 47012 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold411
timestamp 25201
transform -1 0 45172 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold416
timestamp 25201
transform -1 0 77648 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold417
timestamp 25201
transform 1 0 74704 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold418
timestamp 25201
transform -1 0 13432 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold419
timestamp 25201
transform 1 0 16376 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold420
timestamp 25201
transform 1 0 15272 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold421
timestamp 25201
transform 1 0 10488 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold422
timestamp 25201
transform -1 0 16744 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold423
timestamp 25201
transform 1 0 5704 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold424
timestamp 25201
transform -1 0 23828 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold425
timestamp 25201
transform 1 0 10856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold426
timestamp 25201
transform -1 0 23092 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold427
timestamp 25201
transform 1 0 19688 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold428
timestamp 25201
transform 1 0 14536 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold429
timestamp 25201
transform -1 0 18400 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold430
timestamp 25201
transform -1 0 17848 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold431
timestamp 25201
transform 1 0 20608 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold432
timestamp 25201
transform -1 0 27876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold433
timestamp 25201
transform 1 0 17848 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold434
timestamp 25201
transform -1 0 27784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold435
timestamp 25201
transform 1 0 27048 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold436
timestamp 25201
transform 1 0 33304 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold437
timestamp 25201
transform -1 0 47380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold438
timestamp 25201
transform 1 0 35604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold439
timestamp 25201
transform 1 0 34776 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold440
timestamp 25201
transform -1 0 14536 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold441
timestamp 25201
transform 1 0 8280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold442
timestamp 25201
transform 1 0 14168 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold443
timestamp 25201
transform -1 0 23644 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold444
timestamp 25201
transform -1 0 30268 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold445
timestamp 25201
transform -1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold446
timestamp 25201
transform 1 0 21896 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold447
timestamp 25201
transform -1 0 29624 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold448
timestamp 25201
transform -1 0 35696 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold449
timestamp 25201
transform -1 0 34776 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold450
timestamp 25201
transform 1 0 29624 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold451
timestamp 25201
transform 1 0 32568 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold452
timestamp 25201
transform -1 0 37352 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold453
timestamp 25201
transform 1 0 21896 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold454
timestamp 25201
transform 1 0 28888 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold455
timestamp 25201
transform -1 0 36432 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold456
timestamp 25201
transform 1 0 9016 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold457
timestamp 25201
transform -1 0 7176 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold458
timestamp 25201
transform -1 0 20056 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold459
timestamp 25201
transform 1 0 21160 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold460
timestamp 25201
transform 1 0 43332 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold461
timestamp 25201
transform -1 0 48852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold462
timestamp 25201
transform 1 0 41308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold463
timestamp 25201
transform -1 0 42964 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold466
timestamp 25201
transform -1 0 75256 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold467
timestamp 25201
transform -1 0 77464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold468
timestamp 25201
transform -1 0 77556 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold469
timestamp 25201
transform -1 0 33764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold470
timestamp 25201
transform -1 0 34224 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold471
timestamp 25201
transform 1 0 25944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold472
timestamp 25201
transform 1 0 20148 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold473
timestamp 25201
transform -1 0 31280 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold474
timestamp 25201
transform 1 0 20148 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold475
timestamp 25201
transform 1 0 47380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold476
timestamp 25201
transform -1 0 48852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold477
timestamp 25201
transform -1 0 46368 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold478
timestamp 25201
transform -1 0 40204 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold479
timestamp 25201
transform -1 0 39928 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold480
timestamp 25201
transform -1 0 34040 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold484
timestamp 25201
transform 1 0 51704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold485
timestamp 25201
transform 1 0 52072 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold489
timestamp 25201
transform 1 0 53912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold490
timestamp 25201
transform -1 0 56212 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold494
timestamp 25201
transform -1 0 58144 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold495
timestamp 25201
transform -1 0 59616 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold499
timestamp 25201
transform -1 0 65872 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold500
timestamp 25201
transform 1 0 65504 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold504
timestamp 25201
transform -1 0 62100 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold505
timestamp 25201
transform -1 0 63572 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold509
timestamp 25201
transform 1 0 69368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold510
timestamp 25201
transform -1 0 71668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold514
timestamp 25201
transform 1 0 67160 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold515
timestamp 25201
transform 1 0 67528 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold519
timestamp 25201
transform -1 0 72404 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold520
timestamp 25201
transform -1 0 73876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold521
timestamp 25201
transform 1 0 49220 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold522
timestamp 25201
transform -1 0 50324 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold523
timestamp 25201
transform -1 0 47840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold524
timestamp 25201
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold525
timestamp 25201
transform 1 0 4232 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold526
timestamp 25201
transform 1 0 5152 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold530
timestamp 25201
transform -1 0 44896 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold531
timestamp 25201
transform 1 0 18584 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold532
timestamp 25201
transform 1 0 15824 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold533
timestamp 25201
transform 1 0 18584 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold534
timestamp 25201
transform 1 0 10488 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold535
timestamp 25201
transform 1 0 25208 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold536
timestamp 25201
transform 1 0 25576 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold537
timestamp 25201
transform -1 0 38088 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold538
timestamp 25201
transform 1 0 41584 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold539
timestamp 25201
transform 1 0 40756 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold540
timestamp 25201
transform 1 0 40756 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold541
timestamp 25201
transform 1 0 40480 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold542
timestamp 25201
transform -1 0 41492 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold543
timestamp 25201
transform -1 0 40296 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold544
timestamp 25201
transform -1 0 40664 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold545
timestamp 25201
transform -1 0 40848 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold546
timestamp 25201
transform -1 0 34776 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold547
timestamp 25201
transform -1 0 35512 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold548
timestamp 25201
transform 1 0 33304 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold549
timestamp 25201
transform 1 0 30636 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold552
timestamp 25201
transform 1 0 76912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold553
timestamp 25201
transform -1 0 77648 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold554
timestamp 25201
transform 1 0 73416 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold555
timestamp 25201
transform -1 0 37720 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold556
timestamp 25201
transform -1 0 26312 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold557
timestamp 25201
transform -1 0 32108 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold558
timestamp 25201
transform -1 0 26772 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold559
timestamp 25201
transform -1 0 34776 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold560
timestamp 25201
transform -1 0 32476 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold561
timestamp 25201
transform -1 0 28888 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold562
timestamp 25201
transform -1 0 23920 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold563
timestamp 25201
transform -1 0 32936 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold564
timestamp 25201
transform 1 0 31832 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold733
timestamp 25201
transform 1 0 19320 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold734
timestamp 25201
transform -1 0 20424 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold735
timestamp 25201
transform 1 0 38088 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold736
timestamp 25201
transform -1 0 39652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold737
timestamp 25201
transform -1 0 37076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold900
timestamp 25201
transform -1 0 28152 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold920
timestamp 25201
transform -1 0 19688 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold921
timestamp 25201
transform 1 0 11224 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1098
timestamp 25201
transform -1 0 21620 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1099
timestamp 25201
transform -1 0 21252 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1100
timestamp 25201
transform 1 0 13616 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1101
timestamp 25201
transform 1 0 16008 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1278
timestamp 25201
transform 1 0 16744 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1279
timestamp 25201
transform -1 0 21160 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1280
timestamp 25201
transform -1 0 22356 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1458
timestamp 25201
transform -1 0 22264 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1459
timestamp 25201
transform 1 0 12880 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 25201
transform 1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 25201
transform -1 0 28152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 25201
transform -1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 25201
transform 1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 25201
transform 1 0 42044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 25201
transform -1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 25201
transform 1 0 48116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 25201
transform 1 0 13524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 25201
transform 1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 25201
transform 1 0 20240 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 25201
transform 1 0 23460 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 25201
transform -1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 25201
transform 1 0 27876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 25201
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 25201
transform -1 0 21160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 25201
transform -1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 25201
transform -1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 25201
transform -1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 25201
transform 1 0 19688 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 25201
transform 1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 25201
transform 1 0 30452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 25201
transform 1 0 38272 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 25201
transform 1 0 40848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 25201
transform 1 0 45540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 25201
transform -1 0 48392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 25201
transform 1 0 47840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 25201
transform -1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 25201
transform 1 0 22264 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 25201
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 25201
transform -1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 25201
transform -1 0 25576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 25201
transform -1 0 20148 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 25201
transform -1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 25201
transform -1 0 25116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 25201
transform 1 0 32016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 25201
transform -1 0 12696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap102
timestamp 25201
transform -1 0 23092 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output37
timestamp 25201
transform -1 0 14904 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output38
timestamp 25201
transform 1 0 36156 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output39
timestamp 25201
transform -1 0 39192 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output40
timestamp 25201
transform -1 0 40664 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output41
timestamp 25201
transform 1 0 41768 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output42
timestamp 25201
transform 1 0 43884 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output43
timestamp 25201
transform 1 0 45908 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output44
timestamp 25201
transform -1 0 49956 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output45
timestamp 25201
transform -1 0 53084 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output46
timestamp 25201
transform -1 0 55108 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output47
timestamp 25201
transform 1 0 15272 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output48
timestamp 25201
transform -1 0 58696 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output49
timestamp 25201
transform -1 0 62836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output50
timestamp 25201
transform -1 0 66424 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output51
timestamp 25201
transform -1 0 68540 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output52
timestamp 25201
transform -1 0 70564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output53
timestamp 25201
transform -1 0 73140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output54
timestamp 25201
transform -1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output55
timestamp 25201
transform -1 0 76268 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output56
timestamp 25201
transform 1 0 76176 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output57
timestamp 25201
transform 1 0 22264 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output58
timestamp 25201
transform -1 0 25208 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output59
timestamp 25201
transform 1 0 26312 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output60
timestamp 25201
transform 1 0 28428 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output61
timestamp 25201
transform -1 0 31924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output62
timestamp 25201
transform 1 0 31464 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output63
timestamp 25201
transform 1 0 34040 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 25201
transform 1 0 59340 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 25201
transform 1 0 22724 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 25201
transform 1 0 18584 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 25201
transform 1 0 15180 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 25201
transform -1 0 12328 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 25201
transform 1 0 7820 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 25201
transform -1 0 5612 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 25201
transform 1 0 56212 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 25201
transform 1 0 51980 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 25201
transform 1 0 48484 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 25201
transform 1 0 44620 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 25201
transform 1 0 40940 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 25201
transform 1 0 36616 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 25201
transform 1 0 33580 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 25201
transform 1 0 29900 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 25201
transform 1 0 26220 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 25201
transform 1 0 58788 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 25201
transform -1 0 22172 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 25201
transform -1 0 19044 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 25201
transform -1 0 14812 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 25201
transform -1 0 11132 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 25201
transform -1 0 7176 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 25201
transform -1 0 3772 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 25201
transform 1 0 53820 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 25201
transform 1 0 50140 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 25201
transform 1 0 46460 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 25201
transform 1 0 43332 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 25201
transform 1 0 39100 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 25201
transform 1 0 35420 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 25201
transform -1 0 32936 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 25201
transform -1 0 29532 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 25201
transform -1 0 25852 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_65
timestamp 25201
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 25201
transform -1 0 77924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_66
timestamp 25201
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 25201
transform -1 0 77924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_67
timestamp 25201
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 25201
transform -1 0 77924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_68
timestamp 25201
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 25201
transform -1 0 77924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_69
timestamp 25201
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 25201
transform -1 0 77924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_70
timestamp 25201
transform 1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 25201
transform -1 0 77924 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_71
timestamp 25201
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 25201
transform -1 0 77924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_72
timestamp 25201
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 25201
transform -1 0 77924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_73
timestamp 25201
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 25201
transform -1 0 77924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_74
timestamp 25201
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 25201
transform -1 0 77924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_75
timestamp 25201
transform 1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 25201
transform -1 0 77924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_76
timestamp 25201
transform 1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 25201
transform -1 0 77924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_77
timestamp 25201
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 25201
transform -1 0 77924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_78
timestamp 25201
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 25201
transform -1 0 77924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_79
timestamp 25201
transform 1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 25201
transform -1 0 77924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_80
timestamp 25201
transform 1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 25201
transform -1 0 77924 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_81
timestamp 25201
transform 1 0 2024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 25201
transform -1 0 77924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_82
timestamp 25201
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 25201
transform -1 0 77924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_83
timestamp 25201
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 25201
transform -1 0 77924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_84
timestamp 25201
transform 1 0 2024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 25201
transform -1 0 77924 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_85
timestamp 25201
transform 1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 25201
transform -1 0 77924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_86
timestamp 25201
transform 1 0 2024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 25201
transform -1 0 77924 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_87
timestamp 25201
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 25201
transform -1 0 77924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_88
timestamp 25201
transform 1 0 2024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 25201
transform -1 0 77924 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_89
timestamp 25201
transform 1 0 2024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 25201
transform -1 0 77924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_90
timestamp 25201
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 25201
transform -1 0 77924 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_91
timestamp 25201
transform 1 0 2024 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 25201
transform -1 0 77924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_92
timestamp 25201
transform 1 0 2024 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 25201
transform -1 0 77924 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_93
timestamp 25201
transform 1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 25201
transform -1 0 77924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_94
timestamp 25201
transform 1 0 2024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 25201
transform -1 0 77924 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_95
timestamp 25201
transform 1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 25201
transform -1 0 77924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_96
timestamp 25201
transform 1 0 2024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 25201
transform -1 0 77924 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_97
timestamp 25201
transform 1 0 2024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 25201
transform -1 0 77924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_98
timestamp 25201
transform 1 0 2024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 25201
transform -1 0 77924 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_99
timestamp 25201
transform 1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 25201
transform -1 0 77924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_100
timestamp 25201
transform 1 0 2024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 25201
transform -1 0 77924 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_101
timestamp 25201
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 25201
transform -1 0 77924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_102
timestamp 25201
transform 1 0 2024 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 25201
transform -1 0 77924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_103
timestamp 25201
transform 1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 25201
transform -1 0 77924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_104
timestamp 25201
transform 1 0 2024 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 25201
transform -1 0 77924 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_105
timestamp 25201
transform 1 0 2024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 25201
transform -1 0 77924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_106
timestamp 25201
transform 1 0 2024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 25201
transform -1 0 77924 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_107
timestamp 25201
transform 1 0 2024 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 25201
transform -1 0 77924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_108
timestamp 25201
transform 1 0 2024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 25201
transform -1 0 77924 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_109
timestamp 25201
transform 1 0 2024 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 25201
transform -1 0 77924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_110
timestamp 25201
transform 1 0 2024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 25201
transform -1 0 77924 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_111
timestamp 25201
transform 1 0 2024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 25201
transform -1 0 77924 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_112
timestamp 25201
transform 1 0 2024 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 25201
transform -1 0 77924 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_113
timestamp 25201
transform 1 0 2024 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 25201
transform -1 0 77924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_114
timestamp 25201
transform 1 0 2024 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 25201
transform -1 0 77924 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_115
timestamp 25201
transform 1 0 2024 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 25201
transform -1 0 77924 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_116
timestamp 25201
transform 1 0 2024 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 25201
transform -1 0 77924 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_117
timestamp 25201
transform 1 0 2024 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 25201
transform -1 0 77924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_118
timestamp 25201
transform 1 0 2024 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 25201
transform -1 0 77924 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_119
timestamp 25201
transform 1 0 2024 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 25201
transform -1 0 77924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_120
timestamp 25201
transform 1 0 2024 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 25201
transform -1 0 77924 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_121
timestamp 25201
transform 1 0 2024 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 25201
transform -1 0 77924 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_122
timestamp 25201
transform 1 0 2024 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 25201
transform -1 0 77924 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_123
timestamp 25201
transform 1 0 2024 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 25201
transform -1 0 77924 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_124
timestamp 25201
transform 1 0 2024 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 25201
transform -1 0 77924 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_125
timestamp 25201
transform 1 0 2024 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 25201
transform -1 0 77924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_126
timestamp 25201
transform 1 0 2024 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 25201
transform -1 0 77924 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_127
timestamp 25201
transform 1 0 2024 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 25201
transform -1 0 77924 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_128
timestamp 25201
transform 1 0 2024 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 25201
transform -1 0 77924 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_129
timestamp 25201
transform 1 0 2024 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 25201
transform -1 0 77924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_130
timestamp 25201
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_131
timestamp 25201
transform 1 0 7176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp 25201
transform 1 0 9752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp 25201
transform 1 0 12328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp 25201
transform 1 0 14904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp 25201
transform 1 0 17480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp 25201
transform 1 0 20056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_137
timestamp 25201
transform 1 0 22632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138
timestamp 25201
transform 1 0 25208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 25201
transform 1 0 27784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 25201
transform 1 0 30360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 25201
transform 1 0 32936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 25201
transform 1 0 35512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_143
timestamp 25201
transform 1 0 38088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_144
timestamp 25201
transform 1 0 40664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_145
timestamp 25201
transform 1 0 43240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_146
timestamp 25201
transform 1 0 45816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_147
timestamp 25201
transform 1 0 48392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_148
timestamp 25201
transform 1 0 50968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_149
timestamp 25201
transform 1 0 53544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_150
timestamp 25201
transform 1 0 56120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_151
timestamp 25201
transform 1 0 58696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_152
timestamp 25201
transform 1 0 61272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_153
timestamp 25201
transform 1 0 63848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_154
timestamp 25201
transform 1 0 66424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_155
timestamp 25201
transform 1 0 69000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_156
timestamp 25201
transform 1 0 71576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_157
timestamp 25201
transform 1 0 74152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_158
timestamp 25201
transform 1 0 76728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_159
timestamp 25201
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_160
timestamp 25201
transform 1 0 12328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_161
timestamp 25201
transform 1 0 17480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_162
timestamp 25201
transform 1 0 22632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_163
timestamp 25201
transform 1 0 27784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_164
timestamp 25201
transform 1 0 32936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_165
timestamp 25201
transform 1 0 38088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_166
timestamp 25201
transform 1 0 43240 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_167
timestamp 25201
transform 1 0 48392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_168
timestamp 25201
transform 1 0 53544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_169
timestamp 25201
transform 1 0 58696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_170
timestamp 25201
transform 1 0 63848 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_171
timestamp 25201
transform 1 0 69000 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_172
timestamp 25201
transform 1 0 74152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_173
timestamp 25201
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_174
timestamp 25201
transform 1 0 9752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_175
timestamp 25201
transform 1 0 14904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_176
timestamp 25201
transform 1 0 20056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_177
timestamp 25201
transform 1 0 25208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_178
timestamp 25201
transform 1 0 30360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_179
timestamp 25201
transform 1 0 35512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_180
timestamp 25201
transform 1 0 40664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_181
timestamp 25201
transform 1 0 45816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_182
timestamp 25201
transform 1 0 50968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_183
timestamp 25201
transform 1 0 56120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_184
timestamp 25201
transform 1 0 61272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_185
timestamp 25201
transform 1 0 66424 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_186
timestamp 25201
transform 1 0 71576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_187
timestamp 25201
transform 1 0 76728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_188
timestamp 25201
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_189
timestamp 25201
transform 1 0 12328 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_190
timestamp 25201
transform 1 0 17480 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_191
timestamp 25201
transform 1 0 22632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_192
timestamp 25201
transform 1 0 27784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_193
timestamp 25201
transform 1 0 32936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_194
timestamp 25201
transform 1 0 38088 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_195
timestamp 25201
transform 1 0 43240 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_196
timestamp 25201
transform 1 0 48392 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_197
timestamp 25201
transform 1 0 53544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_198
timestamp 25201
transform 1 0 58696 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_199
timestamp 25201
transform 1 0 63848 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_200
timestamp 25201
transform 1 0 69000 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_201
timestamp 25201
transform 1 0 74152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_202
timestamp 25201
transform 1 0 4600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_203
timestamp 25201
transform 1 0 9752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_204
timestamp 25201
transform 1 0 14904 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_205
timestamp 25201
transform 1 0 20056 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_206
timestamp 25201
transform 1 0 25208 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_207
timestamp 25201
transform 1 0 30360 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_208
timestamp 25201
transform 1 0 35512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_209
timestamp 25201
transform 1 0 40664 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_210
timestamp 25201
transform 1 0 45816 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_211
timestamp 25201
transform 1 0 50968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_212
timestamp 25201
transform 1 0 56120 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_213
timestamp 25201
transform 1 0 61272 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_214
timestamp 25201
transform 1 0 66424 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_215
timestamp 25201
transform 1 0 71576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_216
timestamp 25201
transform 1 0 76728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_217
timestamp 25201
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_218
timestamp 25201
transform 1 0 12328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_219
timestamp 25201
transform 1 0 17480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_220
timestamp 25201
transform 1 0 22632 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_221
timestamp 25201
transform 1 0 27784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_222
timestamp 25201
transform 1 0 32936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_223
timestamp 25201
transform 1 0 38088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_224
timestamp 25201
transform 1 0 43240 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_225
timestamp 25201
transform 1 0 48392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_226
timestamp 25201
transform 1 0 53544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_227
timestamp 25201
transform 1 0 58696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_228
timestamp 25201
transform 1 0 63848 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_229
timestamp 25201
transform 1 0 69000 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_230
timestamp 25201
transform 1 0 74152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_231
timestamp 25201
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_232
timestamp 25201
transform 1 0 9752 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_233
timestamp 25201
transform 1 0 14904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_234
timestamp 25201
transform 1 0 20056 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_235
timestamp 25201
transform 1 0 25208 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_236
timestamp 25201
transform 1 0 30360 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_237
timestamp 25201
transform 1 0 35512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_238
timestamp 25201
transform 1 0 40664 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_239
timestamp 25201
transform 1 0 45816 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_240
timestamp 25201
transform 1 0 50968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_241
timestamp 25201
transform 1 0 56120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_242
timestamp 25201
transform 1 0 61272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_243
timestamp 25201
transform 1 0 66424 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_244
timestamp 25201
transform 1 0 71576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_245
timestamp 25201
transform 1 0 76728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_246
timestamp 25201
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_247
timestamp 25201
transform 1 0 12328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_248
timestamp 25201
transform 1 0 17480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_249
timestamp 25201
transform 1 0 22632 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_250
timestamp 25201
transform 1 0 27784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_251
timestamp 25201
transform 1 0 32936 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_252
timestamp 25201
transform 1 0 38088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_253
timestamp 25201
transform 1 0 43240 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_254
timestamp 25201
transform 1 0 48392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_255
timestamp 25201
transform 1 0 53544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_256
timestamp 25201
transform 1 0 58696 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_257
timestamp 25201
transform 1 0 63848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_258
timestamp 25201
transform 1 0 69000 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_259
timestamp 25201
transform 1 0 74152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_260
timestamp 25201
transform 1 0 4600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_261
timestamp 25201
transform 1 0 9752 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_262
timestamp 25201
transform 1 0 14904 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_263
timestamp 25201
transform 1 0 20056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_264
timestamp 25201
transform 1 0 25208 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_265
timestamp 25201
transform 1 0 30360 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_266
timestamp 25201
transform 1 0 35512 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_267
timestamp 25201
transform 1 0 40664 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_268
timestamp 25201
transform 1 0 45816 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_269
timestamp 25201
transform 1 0 50968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_270
timestamp 25201
transform 1 0 56120 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_271
timestamp 25201
transform 1 0 61272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_272
timestamp 25201
transform 1 0 66424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_273
timestamp 25201
transform 1 0 71576 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_274
timestamp 25201
transform 1 0 76728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_275
timestamp 25201
transform 1 0 7176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_276
timestamp 25201
transform 1 0 12328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_277
timestamp 25201
transform 1 0 17480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_278
timestamp 25201
transform 1 0 22632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_279
timestamp 25201
transform 1 0 27784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_280
timestamp 25201
transform 1 0 32936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_281
timestamp 25201
transform 1 0 38088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_282
timestamp 25201
transform 1 0 43240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_283
timestamp 25201
transform 1 0 48392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_284
timestamp 25201
transform 1 0 53544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_285
timestamp 25201
transform 1 0 58696 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_286
timestamp 25201
transform 1 0 63848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_287
timestamp 25201
transform 1 0 69000 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_288
timestamp 25201
transform 1 0 74152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_289
timestamp 25201
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_290
timestamp 25201
transform 1 0 9752 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_291
timestamp 25201
transform 1 0 14904 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_292
timestamp 25201
transform 1 0 20056 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_293
timestamp 25201
transform 1 0 25208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_294
timestamp 25201
transform 1 0 30360 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_295
timestamp 25201
transform 1 0 35512 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_296
timestamp 25201
transform 1 0 40664 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_297
timestamp 25201
transform 1 0 45816 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_298
timestamp 25201
transform 1 0 50968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_299
timestamp 25201
transform 1 0 56120 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_300
timestamp 25201
transform 1 0 61272 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_301
timestamp 25201
transform 1 0 66424 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_302
timestamp 25201
transform 1 0 71576 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_303
timestamp 25201
transform 1 0 76728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_304
timestamp 25201
transform 1 0 7176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_305
timestamp 25201
transform 1 0 12328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_306
timestamp 25201
transform 1 0 17480 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_307
timestamp 25201
transform 1 0 22632 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_308
timestamp 25201
transform 1 0 27784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_309
timestamp 25201
transform 1 0 32936 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_310
timestamp 25201
transform 1 0 38088 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_311
timestamp 25201
transform 1 0 43240 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_312
timestamp 25201
transform 1 0 48392 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_313
timestamp 25201
transform 1 0 53544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_314
timestamp 25201
transform 1 0 58696 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_315
timestamp 25201
transform 1 0 63848 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_316
timestamp 25201
transform 1 0 69000 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_317
timestamp 25201
transform 1 0 74152 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_318
timestamp 25201
transform 1 0 4600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_319
timestamp 25201
transform 1 0 9752 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_320
timestamp 25201
transform 1 0 14904 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_321
timestamp 25201
transform 1 0 20056 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_322
timestamp 25201
transform 1 0 25208 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_323
timestamp 25201
transform 1 0 30360 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_324
timestamp 25201
transform 1 0 35512 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_325
timestamp 25201
transform 1 0 40664 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_326
timestamp 25201
transform 1 0 45816 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_327
timestamp 25201
transform 1 0 50968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_328
timestamp 25201
transform 1 0 56120 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_329
timestamp 25201
transform 1 0 61272 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_330
timestamp 25201
transform 1 0 66424 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_331
timestamp 25201
transform 1 0 71576 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_332
timestamp 25201
transform 1 0 76728 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_333
timestamp 25201
transform 1 0 7176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_334
timestamp 25201
transform 1 0 12328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_335
timestamp 25201
transform 1 0 17480 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_336
timestamp 25201
transform 1 0 22632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_337
timestamp 25201
transform 1 0 27784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_338
timestamp 25201
transform 1 0 32936 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_339
timestamp 25201
transform 1 0 38088 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_340
timestamp 25201
transform 1 0 43240 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_341
timestamp 25201
transform 1 0 48392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_342
timestamp 25201
transform 1 0 53544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_343
timestamp 25201
transform 1 0 58696 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_344
timestamp 25201
transform 1 0 63848 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_345
timestamp 25201
transform 1 0 69000 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_346
timestamp 25201
transform 1 0 74152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_347
timestamp 25201
transform 1 0 4600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_348
timestamp 25201
transform 1 0 9752 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_349
timestamp 25201
transform 1 0 14904 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_350
timestamp 25201
transform 1 0 20056 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_351
timestamp 25201
transform 1 0 25208 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_352
timestamp 25201
transform 1 0 30360 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_353
timestamp 25201
transform 1 0 35512 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_354
timestamp 25201
transform 1 0 40664 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_355
timestamp 25201
transform 1 0 45816 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_356
timestamp 25201
transform 1 0 50968 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_357
timestamp 25201
transform 1 0 56120 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_358
timestamp 25201
transform 1 0 61272 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_359
timestamp 25201
transform 1 0 66424 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_360
timestamp 25201
transform 1 0 71576 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_361
timestamp 25201
transform 1 0 76728 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_362
timestamp 25201
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_363
timestamp 25201
transform 1 0 12328 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_364
timestamp 25201
transform 1 0 17480 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_365
timestamp 25201
transform 1 0 22632 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_366
timestamp 25201
transform 1 0 27784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_367
timestamp 25201
transform 1 0 32936 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_368
timestamp 25201
transform 1 0 38088 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_369
timestamp 25201
transform 1 0 43240 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_370
timestamp 25201
transform 1 0 48392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_371
timestamp 25201
transform 1 0 53544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_372
timestamp 25201
transform 1 0 58696 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_373
timestamp 25201
transform 1 0 63848 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_374
timestamp 25201
transform 1 0 69000 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_375
timestamp 25201
transform 1 0 74152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_376
timestamp 25201
transform 1 0 4600 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_377
timestamp 25201
transform 1 0 9752 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_378
timestamp 25201
transform 1 0 14904 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_379
timestamp 25201
transform 1 0 20056 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_380
timestamp 25201
transform 1 0 25208 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_381
timestamp 25201
transform 1 0 30360 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_382
timestamp 25201
transform 1 0 35512 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_383
timestamp 25201
transform 1 0 40664 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_384
timestamp 25201
transform 1 0 45816 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_385
timestamp 25201
transform 1 0 50968 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_386
timestamp 25201
transform 1 0 56120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_387
timestamp 25201
transform 1 0 61272 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_388
timestamp 25201
transform 1 0 66424 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_389
timestamp 25201
transform 1 0 71576 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_390
timestamp 25201
transform 1 0 76728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_391
timestamp 25201
transform 1 0 7176 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_392
timestamp 25201
transform 1 0 12328 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_393
timestamp 25201
transform 1 0 17480 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_394
timestamp 25201
transform 1 0 22632 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_395
timestamp 25201
transform 1 0 27784 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_396
timestamp 25201
transform 1 0 32936 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_397
timestamp 25201
transform 1 0 38088 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_398
timestamp 25201
transform 1 0 43240 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_399
timestamp 25201
transform 1 0 48392 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_400
timestamp 25201
transform 1 0 53544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_401
timestamp 25201
transform 1 0 58696 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_402
timestamp 25201
transform 1 0 63848 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_403
timestamp 25201
transform 1 0 69000 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_404
timestamp 25201
transform 1 0 74152 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_405
timestamp 25201
transform 1 0 4600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_406
timestamp 25201
transform 1 0 9752 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_407
timestamp 25201
transform 1 0 14904 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_408
timestamp 25201
transform 1 0 20056 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_409
timestamp 25201
transform 1 0 25208 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_410
timestamp 25201
transform 1 0 30360 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_411
timestamp 25201
transform 1 0 35512 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_412
timestamp 25201
transform 1 0 40664 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_413
timestamp 25201
transform 1 0 45816 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_414
timestamp 25201
transform 1 0 50968 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_415
timestamp 25201
transform 1 0 56120 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_416
timestamp 25201
transform 1 0 61272 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_417
timestamp 25201
transform 1 0 66424 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_418
timestamp 25201
transform 1 0 71576 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_419
timestamp 25201
transform 1 0 76728 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_420
timestamp 25201
transform 1 0 7176 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_421
timestamp 25201
transform 1 0 12328 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_422
timestamp 25201
transform 1 0 17480 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_423
timestamp 25201
transform 1 0 22632 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_424
timestamp 25201
transform 1 0 27784 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_425
timestamp 25201
transform 1 0 32936 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_426
timestamp 25201
transform 1 0 38088 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_427
timestamp 25201
transform 1 0 43240 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_428
timestamp 25201
transform 1 0 48392 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_429
timestamp 25201
transform 1 0 53544 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_430
timestamp 25201
transform 1 0 58696 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_431
timestamp 25201
transform 1 0 63848 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_432
timestamp 25201
transform 1 0 69000 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_433
timestamp 25201
transform 1 0 74152 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_434
timestamp 25201
transform 1 0 4600 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_435
timestamp 25201
transform 1 0 9752 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_436
timestamp 25201
transform 1 0 14904 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_437
timestamp 25201
transform 1 0 20056 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_438
timestamp 25201
transform 1 0 25208 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_439
timestamp 25201
transform 1 0 30360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_440
timestamp 25201
transform 1 0 35512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_441
timestamp 25201
transform 1 0 40664 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_442
timestamp 25201
transform 1 0 45816 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_443
timestamp 25201
transform 1 0 50968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_444
timestamp 25201
transform 1 0 56120 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_445
timestamp 25201
transform 1 0 61272 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_446
timestamp 25201
transform 1 0 66424 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_447
timestamp 25201
transform 1 0 71576 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_448
timestamp 25201
transform 1 0 76728 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_449
timestamp 25201
transform 1 0 7176 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_450
timestamp 25201
transform 1 0 12328 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_451
timestamp 25201
transform 1 0 17480 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_452
timestamp 25201
transform 1 0 22632 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_453
timestamp 25201
transform 1 0 27784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_454
timestamp 25201
transform 1 0 32936 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_455
timestamp 25201
transform 1 0 38088 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_456
timestamp 25201
transform 1 0 43240 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_457
timestamp 25201
transform 1 0 48392 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_458
timestamp 25201
transform 1 0 53544 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_459
timestamp 25201
transform 1 0 58696 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_460
timestamp 25201
transform 1 0 63848 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_461
timestamp 25201
transform 1 0 69000 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_462
timestamp 25201
transform 1 0 74152 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_463
timestamp 25201
transform 1 0 4600 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_464
timestamp 25201
transform 1 0 9752 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_465
timestamp 25201
transform 1 0 14904 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_466
timestamp 25201
transform 1 0 20056 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_467
timestamp 25201
transform 1 0 25208 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_468
timestamp 25201
transform 1 0 30360 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_469
timestamp 25201
transform 1 0 35512 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_470
timestamp 25201
transform 1 0 40664 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_471
timestamp 25201
transform 1 0 45816 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_472
timestamp 25201
transform 1 0 50968 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_473
timestamp 25201
transform 1 0 56120 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_474
timestamp 25201
transform 1 0 61272 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_475
timestamp 25201
transform 1 0 66424 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_476
timestamp 25201
transform 1 0 71576 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_477
timestamp 25201
transform 1 0 76728 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_478
timestamp 25201
transform 1 0 7176 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_479
timestamp 25201
transform 1 0 12328 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_480
timestamp 25201
transform 1 0 17480 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_481
timestamp 25201
transform 1 0 22632 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_482
timestamp 25201
transform 1 0 27784 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_483
timestamp 25201
transform 1 0 32936 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_484
timestamp 25201
transform 1 0 38088 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_485
timestamp 25201
transform 1 0 43240 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_486
timestamp 25201
transform 1 0 48392 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_487
timestamp 25201
transform 1 0 53544 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_488
timestamp 25201
transform 1 0 58696 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_489
timestamp 25201
transform 1 0 63848 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_490
timestamp 25201
transform 1 0 69000 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_491
timestamp 25201
transform 1 0 74152 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_492
timestamp 25201
transform 1 0 4600 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_493
timestamp 25201
transform 1 0 9752 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_494
timestamp 25201
transform 1 0 14904 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_495
timestamp 25201
transform 1 0 20056 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_496
timestamp 25201
transform 1 0 25208 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_497
timestamp 25201
transform 1 0 30360 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_498
timestamp 25201
transform 1 0 35512 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_499
timestamp 25201
transform 1 0 40664 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_500
timestamp 25201
transform 1 0 45816 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_501
timestamp 25201
transform 1 0 50968 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_502
timestamp 25201
transform 1 0 56120 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_503
timestamp 25201
transform 1 0 61272 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_504
timestamp 25201
transform 1 0 66424 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_505
timestamp 25201
transform 1 0 71576 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_506
timestamp 25201
transform 1 0 76728 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_507
timestamp 25201
transform 1 0 7176 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_508
timestamp 25201
transform 1 0 12328 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_509
timestamp 25201
transform 1 0 17480 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_510
timestamp 25201
transform 1 0 22632 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_511
timestamp 25201
transform 1 0 27784 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_512
timestamp 25201
transform 1 0 32936 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_513
timestamp 25201
transform 1 0 38088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_514
timestamp 25201
transform 1 0 43240 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_515
timestamp 25201
transform 1 0 48392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_516
timestamp 25201
transform 1 0 53544 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_517
timestamp 25201
transform 1 0 58696 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_518
timestamp 25201
transform 1 0 63848 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_519
timestamp 25201
transform 1 0 69000 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_520
timestamp 25201
transform 1 0 74152 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_521
timestamp 25201
transform 1 0 4600 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_522
timestamp 25201
transform 1 0 9752 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_523
timestamp 25201
transform 1 0 14904 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_524
timestamp 25201
transform 1 0 20056 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_525
timestamp 25201
transform 1 0 25208 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_526
timestamp 25201
transform 1 0 30360 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_527
timestamp 25201
transform 1 0 35512 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_528
timestamp 25201
transform 1 0 40664 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_529
timestamp 25201
transform 1 0 45816 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_530
timestamp 25201
transform 1 0 50968 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_531
timestamp 25201
transform 1 0 56120 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_532
timestamp 25201
transform 1 0 61272 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_533
timestamp 25201
transform 1 0 66424 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_534
timestamp 25201
transform 1 0 71576 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_535
timestamp 25201
transform 1 0 76728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_536
timestamp 25201
transform 1 0 7176 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_537
timestamp 25201
transform 1 0 12328 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_538
timestamp 25201
transform 1 0 17480 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_539
timestamp 25201
transform 1 0 22632 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_540
timestamp 25201
transform 1 0 27784 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_541
timestamp 25201
transform 1 0 32936 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_542
timestamp 25201
transform 1 0 38088 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_543
timestamp 25201
transform 1 0 43240 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_544
timestamp 25201
transform 1 0 48392 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_545
timestamp 25201
transform 1 0 53544 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_546
timestamp 25201
transform 1 0 58696 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_547
timestamp 25201
transform 1 0 63848 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_548
timestamp 25201
transform 1 0 69000 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_549
timestamp 25201
transform 1 0 74152 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_550
timestamp 25201
transform 1 0 4600 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_551
timestamp 25201
transform 1 0 9752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_552
timestamp 25201
transform 1 0 14904 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_553
timestamp 25201
transform 1 0 20056 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_554
timestamp 25201
transform 1 0 25208 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_555
timestamp 25201
transform 1 0 30360 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_556
timestamp 25201
transform 1 0 35512 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_557
timestamp 25201
transform 1 0 40664 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_558
timestamp 25201
transform 1 0 45816 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_559
timestamp 25201
transform 1 0 50968 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_560
timestamp 25201
transform 1 0 56120 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_561
timestamp 25201
transform 1 0 61272 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_562
timestamp 25201
transform 1 0 66424 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_563
timestamp 25201
transform 1 0 71576 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_564
timestamp 25201
transform 1 0 76728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_565
timestamp 25201
transform 1 0 7176 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_566
timestamp 25201
transform 1 0 12328 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_567
timestamp 25201
transform 1 0 17480 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_568
timestamp 25201
transform 1 0 22632 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_569
timestamp 25201
transform 1 0 27784 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_570
timestamp 25201
transform 1 0 32936 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_571
timestamp 25201
transform 1 0 38088 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_572
timestamp 25201
transform 1 0 43240 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_573
timestamp 25201
transform 1 0 48392 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_574
timestamp 25201
transform 1 0 53544 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_575
timestamp 25201
transform 1 0 58696 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_576
timestamp 25201
transform 1 0 63848 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_577
timestamp 25201
transform 1 0 69000 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_578
timestamp 25201
transform 1 0 74152 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_579
timestamp 25201
transform 1 0 4600 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_580
timestamp 25201
transform 1 0 9752 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_581
timestamp 25201
transform 1 0 14904 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_582
timestamp 25201
transform 1 0 20056 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_583
timestamp 25201
transform 1 0 25208 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_584
timestamp 25201
transform 1 0 30360 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_585
timestamp 25201
transform 1 0 35512 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_586
timestamp 25201
transform 1 0 40664 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_587
timestamp 25201
transform 1 0 45816 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_588
timestamp 25201
transform 1 0 50968 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_589
timestamp 25201
transform 1 0 56120 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_590
timestamp 25201
transform 1 0 61272 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_591
timestamp 25201
transform 1 0 66424 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_592
timestamp 25201
transform 1 0 71576 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_593
timestamp 25201
transform 1 0 76728 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_594
timestamp 25201
transform 1 0 7176 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_595
timestamp 25201
transform 1 0 12328 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_596
timestamp 25201
transform 1 0 17480 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_597
timestamp 25201
transform 1 0 22632 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_598
timestamp 25201
transform 1 0 27784 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_599
timestamp 25201
transform 1 0 32936 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_600
timestamp 25201
transform 1 0 38088 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_601
timestamp 25201
transform 1 0 43240 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_602
timestamp 25201
transform 1 0 48392 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_603
timestamp 25201
transform 1 0 53544 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_604
timestamp 25201
transform 1 0 58696 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_605
timestamp 25201
transform 1 0 63848 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_606
timestamp 25201
transform 1 0 69000 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_607
timestamp 25201
transform 1 0 74152 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_608
timestamp 25201
transform 1 0 4600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_609
timestamp 25201
transform 1 0 9752 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_610
timestamp 25201
transform 1 0 14904 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_611
timestamp 25201
transform 1 0 20056 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_612
timestamp 25201
transform 1 0 25208 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_613
timestamp 25201
transform 1 0 30360 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_614
timestamp 25201
transform 1 0 35512 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_615
timestamp 25201
transform 1 0 40664 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_616
timestamp 25201
transform 1 0 45816 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_617
timestamp 25201
transform 1 0 50968 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_618
timestamp 25201
transform 1 0 56120 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_619
timestamp 25201
transform 1 0 61272 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_620
timestamp 25201
transform 1 0 66424 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_621
timestamp 25201
transform 1 0 71576 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_622
timestamp 25201
transform 1 0 76728 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_623
timestamp 25201
transform 1 0 7176 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_624
timestamp 25201
transform 1 0 12328 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_625
timestamp 25201
transform 1 0 17480 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_626
timestamp 25201
transform 1 0 22632 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_627
timestamp 25201
transform 1 0 27784 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_628
timestamp 25201
transform 1 0 32936 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_629
timestamp 25201
transform 1 0 38088 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_630
timestamp 25201
transform 1 0 43240 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_631
timestamp 25201
transform 1 0 48392 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_632
timestamp 25201
transform 1 0 53544 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_633
timestamp 25201
transform 1 0 58696 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_634
timestamp 25201
transform 1 0 63848 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_635
timestamp 25201
transform 1 0 69000 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_636
timestamp 25201
transform 1 0 74152 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_637
timestamp 25201
transform 1 0 4600 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_638
timestamp 25201
transform 1 0 9752 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_639
timestamp 25201
transform 1 0 14904 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_640
timestamp 25201
transform 1 0 20056 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_641
timestamp 25201
transform 1 0 25208 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_642
timestamp 25201
transform 1 0 30360 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_643
timestamp 25201
transform 1 0 35512 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_644
timestamp 25201
transform 1 0 40664 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_645
timestamp 25201
transform 1 0 45816 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_646
timestamp 25201
transform 1 0 50968 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_647
timestamp 25201
transform 1 0 56120 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_648
timestamp 25201
transform 1 0 61272 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_649
timestamp 25201
transform 1 0 66424 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_650
timestamp 25201
transform 1 0 71576 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_651
timestamp 25201
transform 1 0 76728 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_652
timestamp 25201
transform 1 0 7176 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_653
timestamp 25201
transform 1 0 12328 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_654
timestamp 25201
transform 1 0 17480 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_655
timestamp 25201
transform 1 0 22632 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_656
timestamp 25201
transform 1 0 27784 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_657
timestamp 25201
transform 1 0 32936 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_658
timestamp 25201
transform 1 0 38088 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_659
timestamp 25201
transform 1 0 43240 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_660
timestamp 25201
transform 1 0 48392 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_661
timestamp 25201
transform 1 0 53544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_662
timestamp 25201
transform 1 0 58696 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_663
timestamp 25201
transform 1 0 63848 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_664
timestamp 25201
transform 1 0 69000 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_665
timestamp 25201
transform 1 0 74152 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_666
timestamp 25201
transform 1 0 4600 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_667
timestamp 25201
transform 1 0 9752 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_668
timestamp 25201
transform 1 0 14904 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_669
timestamp 25201
transform 1 0 20056 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_670
timestamp 25201
transform 1 0 25208 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_671
timestamp 25201
transform 1 0 30360 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_672
timestamp 25201
transform 1 0 35512 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_673
timestamp 25201
transform 1 0 40664 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_674
timestamp 25201
transform 1 0 45816 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_675
timestamp 25201
transform 1 0 50968 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_676
timestamp 25201
transform 1 0 56120 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_677
timestamp 25201
transform 1 0 61272 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_678
timestamp 25201
transform 1 0 66424 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_679
timestamp 25201
transform 1 0 71576 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_680
timestamp 25201
transform 1 0 76728 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_681
timestamp 25201
transform 1 0 7176 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_682
timestamp 25201
transform 1 0 12328 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_683
timestamp 25201
transform 1 0 17480 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_684
timestamp 25201
transform 1 0 22632 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_685
timestamp 25201
transform 1 0 27784 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_686
timestamp 25201
transform 1 0 32936 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_687
timestamp 25201
transform 1 0 38088 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_688
timestamp 25201
transform 1 0 43240 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_689
timestamp 25201
transform 1 0 48392 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_690
timestamp 25201
transform 1 0 53544 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_691
timestamp 25201
transform 1 0 58696 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_692
timestamp 25201
transform 1 0 63848 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_693
timestamp 25201
transform 1 0 69000 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_694
timestamp 25201
transform 1 0 74152 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_695
timestamp 25201
transform 1 0 4600 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_696
timestamp 25201
transform 1 0 9752 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_697
timestamp 25201
transform 1 0 14904 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_698
timestamp 25201
transform 1 0 20056 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_699
timestamp 25201
transform 1 0 25208 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_700
timestamp 25201
transform 1 0 30360 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_701
timestamp 25201
transform 1 0 35512 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_702
timestamp 25201
transform 1 0 40664 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_703
timestamp 25201
transform 1 0 45816 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_704
timestamp 25201
transform 1 0 50968 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_705
timestamp 25201
transform 1 0 56120 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_706
timestamp 25201
transform 1 0 61272 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_707
timestamp 25201
transform 1 0 66424 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_708
timestamp 25201
transform 1 0 71576 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_709
timestamp 25201
transform 1 0 76728 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_710
timestamp 25201
transform 1 0 7176 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_711
timestamp 25201
transform 1 0 12328 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_712
timestamp 25201
transform 1 0 17480 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_713
timestamp 25201
transform 1 0 22632 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_714
timestamp 25201
transform 1 0 27784 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_715
timestamp 25201
transform 1 0 32936 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_716
timestamp 25201
transform 1 0 38088 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_717
timestamp 25201
transform 1 0 43240 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_718
timestamp 25201
transform 1 0 48392 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_719
timestamp 25201
transform 1 0 53544 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_720
timestamp 25201
transform 1 0 58696 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_721
timestamp 25201
transform 1 0 63848 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_722
timestamp 25201
transform 1 0 69000 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_723
timestamp 25201
transform 1 0 74152 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_724
timestamp 25201
transform 1 0 4600 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_725
timestamp 25201
transform 1 0 9752 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_726
timestamp 25201
transform 1 0 14904 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_727
timestamp 25201
transform 1 0 20056 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_728
timestamp 25201
transform 1 0 25208 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_729
timestamp 25201
transform 1 0 30360 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_730
timestamp 25201
transform 1 0 35512 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_731
timestamp 25201
transform 1 0 40664 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_732
timestamp 25201
transform 1 0 45816 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_733
timestamp 25201
transform 1 0 50968 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_734
timestamp 25201
transform 1 0 56120 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_735
timestamp 25201
transform 1 0 61272 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_736
timestamp 25201
transform 1 0 66424 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_737
timestamp 25201
transform 1 0 71576 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_738
timestamp 25201
transform 1 0 76728 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_739
timestamp 25201
transform 1 0 7176 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_740
timestamp 25201
transform 1 0 12328 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_741
timestamp 25201
transform 1 0 17480 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_742
timestamp 25201
transform 1 0 22632 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_743
timestamp 25201
transform 1 0 27784 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_744
timestamp 25201
transform 1 0 32936 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_745
timestamp 25201
transform 1 0 38088 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_746
timestamp 25201
transform 1 0 43240 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_747
timestamp 25201
transform 1 0 48392 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_748
timestamp 25201
transform 1 0 53544 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_749
timestamp 25201
transform 1 0 58696 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_750
timestamp 25201
transform 1 0 63848 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_751
timestamp 25201
transform 1 0 69000 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_752
timestamp 25201
transform 1 0 74152 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_753
timestamp 25201
transform 1 0 4600 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_754
timestamp 25201
transform 1 0 9752 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_755
timestamp 25201
transform 1 0 14904 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_756
timestamp 25201
transform 1 0 20056 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_757
timestamp 25201
transform 1 0 25208 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_758
timestamp 25201
transform 1 0 30360 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_759
timestamp 25201
transform 1 0 35512 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_760
timestamp 25201
transform 1 0 40664 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_761
timestamp 25201
transform 1 0 45816 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_762
timestamp 25201
transform 1 0 50968 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_763
timestamp 25201
transform 1 0 56120 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_764
timestamp 25201
transform 1 0 61272 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_765
timestamp 25201
transform 1 0 66424 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_766
timestamp 25201
transform 1 0 71576 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_767
timestamp 25201
transform 1 0 76728 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_768
timestamp 25201
transform 1 0 7176 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_769
timestamp 25201
transform 1 0 12328 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_770
timestamp 25201
transform 1 0 17480 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_771
timestamp 25201
transform 1 0 22632 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_772
timestamp 25201
transform 1 0 27784 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_773
timestamp 25201
transform 1 0 32936 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_774
timestamp 25201
transform 1 0 38088 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_775
timestamp 25201
transform 1 0 43240 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_776
timestamp 25201
transform 1 0 48392 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_777
timestamp 25201
transform 1 0 53544 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_778
timestamp 25201
transform 1 0 58696 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_779
timestamp 25201
transform 1 0 63848 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_780
timestamp 25201
transform 1 0 69000 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_781
timestamp 25201
transform 1 0 74152 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_782
timestamp 25201
transform 1 0 4600 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_783
timestamp 25201
transform 1 0 9752 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_784
timestamp 25201
transform 1 0 14904 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_785
timestamp 25201
transform 1 0 20056 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_786
timestamp 25201
transform 1 0 25208 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_787
timestamp 25201
transform 1 0 30360 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_788
timestamp 25201
transform 1 0 35512 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_789
timestamp 25201
transform 1 0 40664 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_790
timestamp 25201
transform 1 0 45816 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_791
timestamp 25201
transform 1 0 50968 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_792
timestamp 25201
transform 1 0 56120 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_793
timestamp 25201
transform 1 0 61272 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_794
timestamp 25201
transform 1 0 66424 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_795
timestamp 25201
transform 1 0 71576 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_796
timestamp 25201
transform 1 0 76728 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_797
timestamp 25201
transform 1 0 7176 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_798
timestamp 25201
transform 1 0 12328 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_799
timestamp 25201
transform 1 0 17480 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_800
timestamp 25201
transform 1 0 22632 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_801
timestamp 25201
transform 1 0 27784 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_802
timestamp 25201
transform 1 0 32936 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_803
timestamp 25201
transform 1 0 38088 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_804
timestamp 25201
transform 1 0 43240 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_805
timestamp 25201
transform 1 0 48392 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_806
timestamp 25201
transform 1 0 53544 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_807
timestamp 25201
transform 1 0 58696 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_808
timestamp 25201
transform 1 0 63848 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_809
timestamp 25201
transform 1 0 69000 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_810
timestamp 25201
transform 1 0 74152 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_811
timestamp 25201
transform 1 0 4600 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_812
timestamp 25201
transform 1 0 9752 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_813
timestamp 25201
transform 1 0 14904 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_814
timestamp 25201
transform 1 0 20056 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_815
timestamp 25201
transform 1 0 25208 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_816
timestamp 25201
transform 1 0 30360 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_817
timestamp 25201
transform 1 0 35512 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_818
timestamp 25201
transform 1 0 40664 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_819
timestamp 25201
transform 1 0 45816 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_820
timestamp 25201
transform 1 0 50968 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_821
timestamp 25201
transform 1 0 56120 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_822
timestamp 25201
transform 1 0 61272 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_823
timestamp 25201
transform 1 0 66424 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_824
timestamp 25201
transform 1 0 71576 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_825
timestamp 25201
transform 1 0 76728 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_826
timestamp 25201
transform 1 0 7176 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_827
timestamp 25201
transform 1 0 12328 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_828
timestamp 25201
transform 1 0 17480 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_829
timestamp 25201
transform 1 0 22632 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_830
timestamp 25201
transform 1 0 27784 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_831
timestamp 25201
transform 1 0 32936 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_832
timestamp 25201
transform 1 0 38088 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_833
timestamp 25201
transform 1 0 43240 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_834
timestamp 25201
transform 1 0 48392 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_835
timestamp 25201
transform 1 0 53544 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_836
timestamp 25201
transform 1 0 58696 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_837
timestamp 25201
transform 1 0 63848 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_838
timestamp 25201
transform 1 0 69000 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_839
timestamp 25201
transform 1 0 74152 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_840
timestamp 25201
transform 1 0 4600 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_841
timestamp 25201
transform 1 0 9752 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_842
timestamp 25201
transform 1 0 14904 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_843
timestamp 25201
transform 1 0 20056 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_844
timestamp 25201
transform 1 0 25208 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_845
timestamp 25201
transform 1 0 30360 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_846
timestamp 25201
transform 1 0 35512 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_847
timestamp 25201
transform 1 0 40664 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_848
timestamp 25201
transform 1 0 45816 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_849
timestamp 25201
transform 1 0 50968 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_850
timestamp 25201
transform 1 0 56120 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_851
timestamp 25201
transform 1 0 61272 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_852
timestamp 25201
transform 1 0 66424 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_853
timestamp 25201
transform 1 0 71576 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_854
timestamp 25201
transform 1 0 76728 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_855
timestamp 25201
transform 1 0 7176 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_856
timestamp 25201
transform 1 0 12328 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_857
timestamp 25201
transform 1 0 17480 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_858
timestamp 25201
transform 1 0 22632 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_859
timestamp 25201
transform 1 0 27784 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_860
timestamp 25201
transform 1 0 32936 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_861
timestamp 25201
transform 1 0 38088 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_862
timestamp 25201
transform 1 0 43240 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_863
timestamp 25201
transform 1 0 48392 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_864
timestamp 25201
transform 1 0 53544 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_865
timestamp 25201
transform 1 0 58696 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_866
timestamp 25201
transform 1 0 63848 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_867
timestamp 25201
transform 1 0 69000 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_868
timestamp 25201
transform 1 0 74152 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_869
timestamp 25201
transform 1 0 4600 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_870
timestamp 25201
transform 1 0 9752 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_871
timestamp 25201
transform 1 0 14904 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_872
timestamp 25201
transform 1 0 20056 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_873
timestamp 25201
transform 1 0 25208 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_874
timestamp 25201
transform 1 0 30360 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_875
timestamp 25201
transform 1 0 35512 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_876
timestamp 25201
transform 1 0 40664 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_877
timestamp 25201
transform 1 0 45816 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_878
timestamp 25201
transform 1 0 50968 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_879
timestamp 25201
transform 1 0 56120 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_880
timestamp 25201
transform 1 0 61272 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_881
timestamp 25201
transform 1 0 66424 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_882
timestamp 25201
transform 1 0 71576 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_883
timestamp 25201
transform 1 0 76728 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_884
timestamp 25201
transform 1 0 7176 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_885
timestamp 25201
transform 1 0 12328 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_886
timestamp 25201
transform 1 0 17480 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_887
timestamp 25201
transform 1 0 22632 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_888
timestamp 25201
transform 1 0 27784 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_889
timestamp 25201
transform 1 0 32936 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_890
timestamp 25201
transform 1 0 38088 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_891
timestamp 25201
transform 1 0 43240 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_892
timestamp 25201
transform 1 0 48392 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_893
timestamp 25201
transform 1 0 53544 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_894
timestamp 25201
transform 1 0 58696 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_895
timestamp 25201
transform 1 0 63848 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_896
timestamp 25201
transform 1 0 69000 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_897
timestamp 25201
transform 1 0 74152 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_898
timestamp 25201
transform 1 0 4600 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_899
timestamp 25201
transform 1 0 9752 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_900
timestamp 25201
transform 1 0 14904 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_901
timestamp 25201
transform 1 0 20056 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_902
timestamp 25201
transform 1 0 25208 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_903
timestamp 25201
transform 1 0 30360 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_904
timestamp 25201
transform 1 0 35512 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_905
timestamp 25201
transform 1 0 40664 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_906
timestamp 25201
transform 1 0 45816 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_907
timestamp 25201
transform 1 0 50968 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_908
timestamp 25201
transform 1 0 56120 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_909
timestamp 25201
transform 1 0 61272 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_910
timestamp 25201
transform 1 0 66424 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_911
timestamp 25201
transform 1 0 71576 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_912
timestamp 25201
transform 1 0 76728 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_913
timestamp 25201
transform 1 0 7176 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_914
timestamp 25201
transform 1 0 12328 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_915
timestamp 25201
transform 1 0 17480 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_916
timestamp 25201
transform 1 0 22632 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_917
timestamp 25201
transform 1 0 27784 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_918
timestamp 25201
transform 1 0 32936 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_919
timestamp 25201
transform 1 0 38088 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_920
timestamp 25201
transform 1 0 43240 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_921
timestamp 25201
transform 1 0 48392 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_922
timestamp 25201
transform 1 0 53544 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_923
timestamp 25201
transform 1 0 58696 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_924
timestamp 25201
transform 1 0 63848 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_925
timestamp 25201
transform 1 0 69000 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_926
timestamp 25201
transform 1 0 74152 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_927
timestamp 25201
transform 1 0 4600 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_928
timestamp 25201
transform 1 0 9752 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_929
timestamp 25201
transform 1 0 14904 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_930
timestamp 25201
transform 1 0 20056 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_931
timestamp 25201
transform 1 0 25208 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_932
timestamp 25201
transform 1 0 30360 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_933
timestamp 25201
transform 1 0 35512 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_934
timestamp 25201
transform 1 0 40664 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_935
timestamp 25201
transform 1 0 45816 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_936
timestamp 25201
transform 1 0 50968 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_937
timestamp 25201
transform 1 0 56120 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_938
timestamp 25201
transform 1 0 61272 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_939
timestamp 25201
transform 1 0 66424 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_940
timestamp 25201
transform 1 0 71576 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_941
timestamp 25201
transform 1 0 76728 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_942
timestamp 25201
transform 1 0 7176 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_943
timestamp 25201
transform 1 0 12328 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_944
timestamp 25201
transform 1 0 17480 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_945
timestamp 25201
transform 1 0 22632 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_946
timestamp 25201
transform 1 0 27784 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_947
timestamp 25201
transform 1 0 32936 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_948
timestamp 25201
transform 1 0 38088 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_949
timestamp 25201
transform 1 0 43240 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_950
timestamp 25201
transform 1 0 48392 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_951
timestamp 25201
transform 1 0 53544 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_952
timestamp 25201
transform 1 0 58696 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_953
timestamp 25201
transform 1 0 63848 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_954
timestamp 25201
transform 1 0 69000 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_955
timestamp 25201
transform 1 0 74152 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_956
timestamp 25201
transform 1 0 4600 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_957
timestamp 25201
transform 1 0 9752 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_958
timestamp 25201
transform 1 0 14904 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_959
timestamp 25201
transform 1 0 20056 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_960
timestamp 25201
transform 1 0 25208 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_961
timestamp 25201
transform 1 0 30360 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_962
timestamp 25201
transform 1 0 35512 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_963
timestamp 25201
transform 1 0 40664 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_964
timestamp 25201
transform 1 0 45816 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_965
timestamp 25201
transform 1 0 50968 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_966
timestamp 25201
transform 1 0 56120 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_967
timestamp 25201
transform 1 0 61272 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_968
timestamp 25201
transform 1 0 66424 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_969
timestamp 25201
transform 1 0 71576 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_970
timestamp 25201
transform 1 0 76728 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_971
timestamp 25201
transform 1 0 7176 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_972
timestamp 25201
transform 1 0 12328 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_973
timestamp 25201
transform 1 0 17480 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_974
timestamp 25201
transform 1 0 22632 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_975
timestamp 25201
transform 1 0 27784 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_976
timestamp 25201
transform 1 0 32936 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_977
timestamp 25201
transform 1 0 38088 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_978
timestamp 25201
transform 1 0 43240 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_979
timestamp 25201
transform 1 0 48392 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_980
timestamp 25201
transform 1 0 53544 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_981
timestamp 25201
transform 1 0 58696 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_982
timestamp 25201
transform 1 0 63848 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_983
timestamp 25201
transform 1 0 69000 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_984
timestamp 25201
transform 1 0 74152 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_985
timestamp 25201
transform 1 0 4600 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_986
timestamp 25201
transform 1 0 9752 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_987
timestamp 25201
transform 1 0 14904 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_988
timestamp 25201
transform 1 0 20056 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_989
timestamp 25201
transform 1 0 25208 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_990
timestamp 25201
transform 1 0 30360 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_991
timestamp 25201
transform 1 0 35512 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_992
timestamp 25201
transform 1 0 40664 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_993
timestamp 25201
transform 1 0 45816 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_994
timestamp 25201
transform 1 0 50968 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_995
timestamp 25201
transform 1 0 56120 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_996
timestamp 25201
transform 1 0 61272 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_997
timestamp 25201
transform 1 0 66424 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_998
timestamp 25201
transform 1 0 71576 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_999
timestamp 25201
transform 1 0 76728 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1000
timestamp 25201
transform 1 0 7176 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1001
timestamp 25201
transform 1 0 12328 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1002
timestamp 25201
transform 1 0 17480 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1003
timestamp 25201
transform 1 0 22632 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1004
timestamp 25201
transform 1 0 27784 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1005
timestamp 25201
transform 1 0 32936 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1006
timestamp 25201
transform 1 0 38088 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1007
timestamp 25201
transform 1 0 43240 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1008
timestamp 25201
transform 1 0 48392 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1009
timestamp 25201
transform 1 0 53544 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1010
timestamp 25201
transform 1 0 58696 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1011
timestamp 25201
transform 1 0 63848 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1012
timestamp 25201
transform 1 0 69000 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1013
timestamp 25201
transform 1 0 74152 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1014
timestamp 25201
transform 1 0 4600 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1015
timestamp 25201
transform 1 0 9752 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1016
timestamp 25201
transform 1 0 14904 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1017
timestamp 25201
transform 1 0 20056 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1018
timestamp 25201
transform 1 0 25208 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1019
timestamp 25201
transform 1 0 30360 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1020
timestamp 25201
transform 1 0 35512 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1021
timestamp 25201
transform 1 0 40664 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1022
timestamp 25201
transform 1 0 45816 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1023
timestamp 25201
transform 1 0 50968 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1024
timestamp 25201
transform 1 0 56120 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1025
timestamp 25201
transform 1 0 61272 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1026
timestamp 25201
transform 1 0 66424 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1027
timestamp 25201
transform 1 0 71576 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1028
timestamp 25201
transform 1 0 76728 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1029
timestamp 25201
transform 1 0 7176 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1030
timestamp 25201
transform 1 0 12328 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1031
timestamp 25201
transform 1 0 17480 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1032
timestamp 25201
transform 1 0 22632 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1033
timestamp 25201
transform 1 0 27784 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1034
timestamp 25201
transform 1 0 32936 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1035
timestamp 25201
transform 1 0 38088 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1036
timestamp 25201
transform 1 0 43240 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1037
timestamp 25201
transform 1 0 48392 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1038
timestamp 25201
transform 1 0 53544 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1039
timestamp 25201
transform 1 0 58696 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1040
timestamp 25201
transform 1 0 63848 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1041
timestamp 25201
transform 1 0 69000 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1042
timestamp 25201
transform 1 0 74152 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1043
timestamp 25201
transform 1 0 4600 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1044
timestamp 25201
transform 1 0 9752 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1045
timestamp 25201
transform 1 0 14904 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1046
timestamp 25201
transform 1 0 20056 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1047
timestamp 25201
transform 1 0 25208 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1048
timestamp 25201
transform 1 0 30360 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1049
timestamp 25201
transform 1 0 35512 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1050
timestamp 25201
transform 1 0 40664 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1051
timestamp 25201
transform 1 0 45816 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1052
timestamp 25201
transform 1 0 50968 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1053
timestamp 25201
transform 1 0 56120 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1054
timestamp 25201
transform 1 0 61272 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1055
timestamp 25201
transform 1 0 66424 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1056
timestamp 25201
transform 1 0 71576 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1057
timestamp 25201
transform 1 0 76728 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1058
timestamp 25201
transform 1 0 7176 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1059
timestamp 25201
transform 1 0 12328 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1060
timestamp 25201
transform 1 0 17480 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1061
timestamp 25201
transform 1 0 22632 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1062
timestamp 25201
transform 1 0 27784 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1063
timestamp 25201
transform 1 0 32936 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1064
timestamp 25201
transform 1 0 38088 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1065
timestamp 25201
transform 1 0 43240 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1066
timestamp 25201
transform 1 0 48392 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1067
timestamp 25201
transform 1 0 53544 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1068
timestamp 25201
transform 1 0 58696 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1069
timestamp 25201
transform 1 0 63848 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1070
timestamp 25201
transform 1 0 69000 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1071
timestamp 25201
transform 1 0 74152 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1072
timestamp 25201
transform 1 0 4600 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1073
timestamp 25201
transform 1 0 7176 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1074
timestamp 25201
transform 1 0 9752 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1075
timestamp 25201
transform 1 0 12328 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1076
timestamp 25201
transform 1 0 14904 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1077
timestamp 25201
transform 1 0 17480 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1078
timestamp 25201
transform 1 0 20056 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1079
timestamp 25201
transform 1 0 22632 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1080
timestamp 25201
transform 1 0 25208 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1081
timestamp 25201
transform 1 0 27784 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1082
timestamp 25201
transform 1 0 30360 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1083
timestamp 25201
transform 1 0 32936 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1084
timestamp 25201
transform 1 0 35512 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1085
timestamp 25201
transform 1 0 38088 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1086
timestamp 25201
transform 1 0 40664 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1087
timestamp 25201
transform 1 0 43240 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1088
timestamp 25201
transform 1 0 45816 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1089
timestamp 25201
transform 1 0 48392 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1090
timestamp 25201
transform 1 0 50968 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1091
timestamp 25201
transform 1 0 53544 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1092
timestamp 25201
transform 1 0 56120 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1093
timestamp 25201
transform 1 0 58696 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1094
timestamp 25201
transform 1 0 61272 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1095
timestamp 25201
transform 1 0 63848 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1096
timestamp 25201
transform 1 0 66424 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1097
timestamp 25201
transform 1 0 69000 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1098
timestamp 25201
transform 1 0 71576 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1099
timestamp 25201
transform 1 0 74152 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1100
timestamp 25201
transform 1 0 76728 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire103
timestamp 25201
transform -1 0 24840 0 -1 5440
box -38 -48 314 592
<< labels >>
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 HADDR[0]
port 0 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 HADDR[10]
port 1 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 HADDR[11]
port 2 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 HADDR[12]
port 3 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 HADDR[13]
port 4 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 HADDR[14]
port 5 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 HADDR[15]
port 6 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 HADDR[16]
port 7 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 HADDR[17]
port 8 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 HADDR[18]
port 9 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 HADDR[19]
port 10 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 HADDR[1]
port 11 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 HADDR[20]
port 12 nsew signal input
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 HADDR[21]
port 13 nsew signal input
flabel metal2 s 58622 0 58678 800 0 FreeSans 224 90 0 0 HADDR[22]
port 14 nsew signal input
flabel metal2 s 60554 0 60610 800 0 FreeSans 224 90 0 0 HADDR[23]
port 15 nsew signal input
flabel metal2 s 62486 0 62542 800 0 FreeSans 224 90 0 0 HADDR[24]
port 16 nsew signal input
flabel metal2 s 64418 0 64474 800 0 FreeSans 224 90 0 0 HADDR[25]
port 17 nsew signal input
flabel metal2 s 66350 0 66406 800 0 FreeSans 224 90 0 0 HADDR[26]
port 18 nsew signal input
flabel metal2 s 68282 0 68338 800 0 FreeSans 224 90 0 0 HADDR[27]
port 19 nsew signal input
flabel metal2 s 70214 0 70270 800 0 FreeSans 224 90 0 0 HADDR[28]
port 20 nsew signal input
flabel metal2 s 72146 0 72202 800 0 FreeSans 224 90 0 0 HADDR[29]
port 21 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 HADDR[2]
port 22 nsew signal input
flabel metal2 s 74078 0 74134 800 0 FreeSans 224 90 0 0 HADDR[30]
port 23 nsew signal input
flabel metal2 s 76010 0 76066 800 0 FreeSans 224 90 0 0 HADDR[31]
port 24 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 HADDR[3]
port 25 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 HADDR[4]
port 26 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 HADDR[5]
port 27 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 HADDR[6]
port 28 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 HADDR[7]
port 29 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 HADDR[8]
port 30 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 HADDR[9]
port 31 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 HCLK
port 32 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 HRDATA[0]
port 33 nsew signal output
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 HRDATA[10]
port 34 nsew signal output
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 HRDATA[11]
port 35 nsew signal output
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 HRDATA[12]
port 36 nsew signal output
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 HRDATA[13]
port 37 nsew signal output
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 HRDATA[14]
port 38 nsew signal output
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 HRDATA[15]
port 39 nsew signal output
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 HRDATA[16]
port 40 nsew signal output
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 HRDATA[17]
port 41 nsew signal output
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 HRDATA[18]
port 42 nsew signal output
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 HRDATA[19]
port 43 nsew signal output
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 HRDATA[1]
port 44 nsew signal output
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 HRDATA[20]
port 45 nsew signal output
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 HRDATA[21]
port 46 nsew signal output
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 HRDATA[22]
port 47 nsew signal output
flabel metal2 s 61198 0 61254 800 0 FreeSans 224 90 0 0 HRDATA[23]
port 48 nsew signal output
flabel metal2 s 63130 0 63186 800 0 FreeSans 224 90 0 0 HRDATA[24]
port 49 nsew signal output
flabel metal2 s 65062 0 65118 800 0 FreeSans 224 90 0 0 HRDATA[25]
port 50 nsew signal output
flabel metal2 s 66994 0 67050 800 0 FreeSans 224 90 0 0 HRDATA[26]
port 51 nsew signal output
flabel metal2 s 68926 0 68982 800 0 FreeSans 224 90 0 0 HRDATA[27]
port 52 nsew signal output
flabel metal2 s 70858 0 70914 800 0 FreeSans 224 90 0 0 HRDATA[28]
port 53 nsew signal output
flabel metal2 s 72790 0 72846 800 0 FreeSans 224 90 0 0 HRDATA[29]
port 54 nsew signal output
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 HRDATA[2]
port 55 nsew signal output
flabel metal2 s 74722 0 74778 800 0 FreeSans 224 90 0 0 HRDATA[30]
port 56 nsew signal output
flabel metal2 s 76654 0 76710 800 0 FreeSans 224 90 0 0 HRDATA[31]
port 57 nsew signal output
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 HRDATA[3]
port 58 nsew signal output
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 HRDATA[4]
port 59 nsew signal output
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 HRDATA[5]
port 60 nsew signal output
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 HRDATA[6]
port 61 nsew signal output
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 HRDATA[7]
port 62 nsew signal output
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 HRDATA[8]
port 63 nsew signal output
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 HRDATA[9]
port 64 nsew signal output
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 HREADY
port 65 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 HREADYOUT
port 66 nsew signal output
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 HRESETn
port 67 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 HSEL
port 68 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 HSIZE[0]
port 69 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 HSIZE[1]
port 70 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 HSIZE[2]
port 71 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 HTRANS[0]
port 72 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 HTRANS[1]
port 73 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 HWDATA[0]
port 74 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 HWDATA[10]
port 75 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 HWDATA[11]
port 76 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 HWDATA[12]
port 77 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 HWDATA[13]
port 78 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 HWDATA[14]
port 79 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 HWDATA[15]
port 80 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 HWDATA[16]
port 81 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 HWDATA[17]
port 82 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 HWDATA[18]
port 83 nsew signal input
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 HWDATA[19]
port 84 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 HWDATA[1]
port 85 nsew signal input
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 HWDATA[20]
port 86 nsew signal input
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 HWDATA[21]
port 87 nsew signal input
flabel metal2 s 59910 0 59966 800 0 FreeSans 224 90 0 0 HWDATA[22]
port 88 nsew signal input
flabel metal2 s 61842 0 61898 800 0 FreeSans 224 90 0 0 HWDATA[23]
port 89 nsew signal input
flabel metal2 s 63774 0 63830 800 0 FreeSans 224 90 0 0 HWDATA[24]
port 90 nsew signal input
flabel metal2 s 65706 0 65762 800 0 FreeSans 224 90 0 0 HWDATA[25]
port 91 nsew signal input
flabel metal2 s 67638 0 67694 800 0 FreeSans 224 90 0 0 HWDATA[26]
port 92 nsew signal input
flabel metal2 s 69570 0 69626 800 0 FreeSans 224 90 0 0 HWDATA[27]
port 93 nsew signal input
flabel metal2 s 71502 0 71558 800 0 FreeSans 224 90 0 0 HWDATA[28]
port 94 nsew signal input
flabel metal2 s 73434 0 73490 800 0 FreeSans 224 90 0 0 HWDATA[29]
port 95 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 HWDATA[2]
port 96 nsew signal input
flabel metal2 s 75366 0 75422 800 0 FreeSans 224 90 0 0 HWDATA[30]
port 97 nsew signal input
flabel metal2 s 77298 0 77354 800 0 FreeSans 224 90 0 0 HWDATA[31]
port 98 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 HWDATA[3]
port 99 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 HWDATA[4]
port 100 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 HWDATA[5]
port 101 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 HWDATA[6]
port 102 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 HWDATA[7]
port 103 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 HWDATA[8]
port 104 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 HWDATA[9]
port 105 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 HWRITE
port 106 nsew signal input
flabel metal2 s 59266 39200 59322 40000 0 FreeSans 224 90 0 0 gpio_oeb[0]
port 107 nsew signal output
flabel metal2 s 22466 39200 22522 40000 0 FreeSans 224 90 0 0 gpio_oeb[10]
port 108 nsew signal output
flabel metal2 s 18786 39200 18842 40000 0 FreeSans 224 90 0 0 gpio_oeb[11]
port 109 nsew signal output
flabel metal2 s 15106 39200 15162 40000 0 FreeSans 224 90 0 0 gpio_oeb[12]
port 110 nsew signal output
flabel metal2 s 11426 39200 11482 40000 0 FreeSans 224 90 0 0 gpio_oeb[13]
port 111 nsew signal output
flabel metal2 s 7746 39200 7802 40000 0 FreeSans 224 90 0 0 gpio_oeb[14]
port 112 nsew signal output
flabel metal2 s 4066 39200 4122 40000 0 FreeSans 224 90 0 0 gpio_oeb[15]
port 113 nsew signal output
flabel metal2 s 55586 39200 55642 40000 0 FreeSans 224 90 0 0 gpio_oeb[1]
port 114 nsew signal output
flabel metal2 s 51906 39200 51962 40000 0 FreeSans 224 90 0 0 gpio_oeb[2]
port 115 nsew signal output
flabel metal2 s 48226 39200 48282 40000 0 FreeSans 224 90 0 0 gpio_oeb[3]
port 116 nsew signal output
flabel metal2 s 44546 39200 44602 40000 0 FreeSans 224 90 0 0 gpio_oeb[4]
port 117 nsew signal output
flabel metal2 s 40866 39200 40922 40000 0 FreeSans 224 90 0 0 gpio_oeb[5]
port 118 nsew signal output
flabel metal2 s 37186 39200 37242 40000 0 FreeSans 224 90 0 0 gpio_oeb[6]
port 119 nsew signal output
flabel metal2 s 33506 39200 33562 40000 0 FreeSans 224 90 0 0 gpio_oeb[7]
port 120 nsew signal output
flabel metal2 s 29826 39200 29882 40000 0 FreeSans 224 90 0 0 gpio_oeb[8]
port 121 nsew signal output
flabel metal2 s 26146 39200 26202 40000 0 FreeSans 224 90 0 0 gpio_oeb[9]
port 122 nsew signal output
flabel metal2 s 57426 39200 57482 40000 0 FreeSans 224 90 0 0 gpio_out[0]
port 123 nsew signal output
flabel metal2 s 20626 39200 20682 40000 0 FreeSans 224 90 0 0 gpio_out[10]
port 124 nsew signal output
flabel metal2 s 16946 39200 17002 40000 0 FreeSans 224 90 0 0 gpio_out[11]
port 125 nsew signal output
flabel metal2 s 13266 39200 13322 40000 0 FreeSans 224 90 0 0 gpio_out[12]
port 126 nsew signal output
flabel metal2 s 9586 39200 9642 40000 0 FreeSans 224 90 0 0 gpio_out[13]
port 127 nsew signal output
flabel metal2 s 5906 39200 5962 40000 0 FreeSans 224 90 0 0 gpio_out[14]
port 128 nsew signal output
flabel metal2 s 2226 39200 2282 40000 0 FreeSans 224 90 0 0 gpio_out[15]
port 129 nsew signal output
flabel metal2 s 53746 39200 53802 40000 0 FreeSans 224 90 0 0 gpio_out[1]
port 130 nsew signal output
flabel metal2 s 50066 39200 50122 40000 0 FreeSans 224 90 0 0 gpio_out[2]
port 131 nsew signal output
flabel metal2 s 46386 39200 46442 40000 0 FreeSans 224 90 0 0 gpio_out[3]
port 132 nsew signal output
flabel metal2 s 42706 39200 42762 40000 0 FreeSans 224 90 0 0 gpio_out[4]
port 133 nsew signal output
flabel metal2 s 39026 39200 39082 40000 0 FreeSans 224 90 0 0 gpio_out[5]
port 134 nsew signal output
flabel metal2 s 35346 39200 35402 40000 0 FreeSans 224 90 0 0 gpio_out[6]
port 135 nsew signal output
flabel metal2 s 31666 39200 31722 40000 0 FreeSans 224 90 0 0 gpio_out[7]
port 136 nsew signal output
flabel metal2 s 27986 39200 28042 40000 0 FreeSans 224 90 0 0 gpio_out[8]
port 137 nsew signal output
flabel metal2 s 24306 39200 24362 40000 0 FreeSans 224 90 0 0 gpio_out[9]
port 138 nsew signal output
flabel metal4 s 5128 2128 5448 37584 0 FreeSans 1920 90 0 0 vccd1
port 139 nsew power bidirectional
flabel metal4 s 35848 2128 36168 37584 0 FreeSans 1920 90 0 0 vccd1
port 139 nsew power bidirectional
flabel metal4 s 66568 2128 66888 37584 0 FreeSans 1920 90 0 0 vccd1
port 139 nsew power bidirectional
flabel metal4 s 5788 2128 6108 37584 0 FreeSans 1920 90 0 0 vssd1
port 140 nsew ground bidirectional
flabel metal4 s 36508 2128 36828 37584 0 FreeSans 1920 90 0 0 vssd1
port 140 nsew ground bidirectional
flabel metal4 s 67228 2128 67548 37584 0 FreeSans 1920 90 0 0 vssd1
port 140 nsew ground bidirectional
rlabel metal1 39974 37536 39974 37536 0 vccd1
rlabel metal1 39974 36992 39974 36992 0 vssd1
rlabel metal1 21666 9486 21666 9486 0 CTRL_REG
rlabel metal2 12466 4318 12466 4318 0 HADDR[0]
rlabel metal2 35466 1027 35466 1027 0 HADDR[10]
rlabel metal2 37398 823 37398 823 0 HADDR[11]
rlabel metal2 39376 5270 39376 5270 0 HADDR[12]
rlabel metal2 41262 1027 41262 1027 0 HADDR[13]
rlabel metal2 43240 5100 43240 5100 0 HADDR[14]
rlabel metal2 45172 5746 45172 5746 0 HADDR[15]
rlabel metal2 16146 1044 16146 1044 0 HADDR[1]
rlabel metal2 19366 1044 19366 1044 0 HADDR[2]
rlabel metal2 21850 561 21850 561 0 HADDR[3]
rlabel metal2 9614 1258 9614 1258 0 HADDR[4]
rlabel metal2 25806 976 25806 976 0 HADDR[5]
rlabel metal2 27738 1163 27738 1163 0 HADDR[6]
rlabel metal1 21068 5678 21068 5678 0 HADDR[7]
rlabel metal1 31142 10506 31142 10506 0 HADDR[8]
rlabel metal2 33442 527 33442 527 0 HADDR[9]
rlabel metal2 9154 476 9154 476 0 HCLK
rlabel metal2 13570 1554 13570 1554 0 HRDATA[0]
rlabel metal2 36110 1622 36110 1622 0 HRDATA[10]
rlabel metal2 38042 1761 38042 1761 0 HRDATA[11]
rlabel metal2 39974 1622 39974 1622 0 HRDATA[12]
rlabel metal2 41906 1554 41906 1554 0 HRDATA[13]
rlabel metal2 43838 823 43838 823 0 HRDATA[14]
rlabel metal1 46460 2958 46460 2958 0 HRDATA[15]
rlabel metal1 48254 2958 48254 2958 0 HRDATA[16]
rlabel metal2 51566 1826 51566 1826 0 HRDATA[18]
rlabel metal2 53498 1860 53498 1860 0 HRDATA[19]
rlabel metal1 17250 3570 17250 3570 0 HRDATA[1]
rlabel metal2 57362 1554 57362 1554 0 HRDATA[21]
rlabel metal2 61226 1860 61226 1860 0 HRDATA[23]
rlabel metal2 65090 1860 65090 1860 0 HRDATA[25]
rlabel metal2 67022 1826 67022 1826 0 HRDATA[26]
rlabel metal2 68954 1860 68954 1860 0 HRDATA[27]
rlabel metal2 70886 1860 70886 1860 0 HRDATA[28]
rlabel metal2 20010 959 20010 959 0 HRDATA[2]
rlabel metal2 74750 1860 74750 1860 0 HRDATA[30]
rlabel metal2 76682 1435 76682 1435 0 HRDATA[31]
rlabel metal1 22356 2482 22356 2482 0 HRDATA[3]
rlabel metal2 24518 1520 24518 1520 0 HRDATA[4]
rlabel metal2 26450 1860 26450 1860 0 HRDATA[5]
rlabel metal2 28382 1095 28382 1095 0 HRDATA[6]
rlabel metal2 30314 959 30314 959 0 HRDATA[7]
rlabel metal2 32246 1622 32246 1622 0 HRDATA[8]
rlabel metal2 34178 1554 34178 1554 0 HRDATA[9]
rlabel metal2 9706 1078 9706 1078 0 HREADY
rlabel metal2 10994 1027 10994 1027 0 HRESETn
rlabel metal2 11638 1588 11638 1588 0 HSEL
rlabel metal2 18078 1010 18078 1010 0 HTRANS[1]
rlabel metal1 15134 6290 15134 6290 0 HWDATA[0]
rlabel metal2 36754 1095 36754 1095 0 HWDATA[10]
rlabel metal2 38686 1761 38686 1761 0 HWDATA[11]
rlabel metal2 40618 1384 40618 1384 0 HWDATA[12]
rlabel metal2 42550 1761 42550 1761 0 HWDATA[13]
rlabel metal1 44804 4454 44804 4454 0 HWDATA[14]
rlabel metal1 47840 3910 47840 3910 0 HWDATA[15]
rlabel metal2 18722 1367 18722 1367 0 HWDATA[1]
rlabel metal2 21298 1078 21298 1078 0 HWDATA[2]
rlabel metal2 23230 1078 23230 1078 0 HWDATA[3]
rlabel via2 14674 5117 14674 5117 0 HWDATA[4]
rlabel metal2 27002 8449 27002 8449 0 HWDATA[5]
rlabel metal2 29026 1761 29026 1761 0 HWDATA[6]
rlabel metal2 20562 2417 20562 2417 0 HWDATA[7]
rlabel metal1 33258 10574 33258 10574 0 HWDATA[8]
rlabel via3 34845 5100 34845 5100 0 HWDATA[9]
rlabel metal2 12282 1095 12282 1095 0 HWRITE
rlabel metal2 15962 3264 15962 3264 0 _000_
rlabel metal1 20792 5338 20792 5338 0 _001_
rlabel metal1 21442 6970 21442 6970 0 _002_
rlabel metal2 22310 8636 22310 8636 0 _003_
rlabel metal1 21068 7514 21068 7514 0 _004_
rlabel metal1 24426 4794 24426 4794 0 _005_
rlabel metal1 23828 6834 23828 6834 0 _006_
rlabel metal1 26818 6426 26818 6426 0 _007_
rlabel metal1 28336 7514 28336 7514 0 _008_
rlabel metal1 28336 7310 28336 7310 0 _009_
rlabel metal2 25346 5984 25346 5984 0 _010_
rlabel metal2 32246 7990 32246 7990 0 _011_
rlabel metal2 33626 6630 33626 6630 0 _012_
rlabel metal1 36570 7412 36570 7412 0 _013_
rlabel metal1 36708 4794 36708 4794 0 _014_
rlabel metal1 36800 5338 36800 5338 0 _015_
rlabel metal2 29026 3502 29026 3502 0 _016_
rlabel metal1 34914 5814 34914 5814 0 _017_
rlabel metal1 11178 2278 11178 2278 0 _018_
rlabel metal1 12282 2618 12282 2618 0 _019_
rlabel metal1 13846 3468 13846 3468 0 _020_
rlabel metal2 17618 2108 17618 2108 0 _021_
rlabel metal2 19090 5083 19090 5083 0 _022_
rlabel metal1 20700 3910 20700 3910 0 _023_
rlabel metal1 23322 4794 23322 4794 0 _024_
rlabel via2 25714 3349 25714 3349 0 _025_
rlabel metal1 27968 4794 27968 4794 0 _026_
rlabel metal2 29900 3910 29900 3910 0 _027_
rlabel metal1 31326 4794 31326 4794 0 _028_
rlabel metal2 33074 2873 33074 2873 0 _029_
rlabel metal2 34730 3995 34730 3995 0 _030_
rlabel metal2 33166 2655 33166 2655 0 _031_
rlabel metal1 40020 3910 40020 3910 0 _032_
rlabel metal1 41538 7310 41538 7310 0 _033_
rlabel metal1 45586 4012 45586 4012 0 _034_
rlabel metal1 43792 3162 43792 3162 0 _035_
rlabel metal3 23598 10812 23598 10812 0 _036_
rlabel metal1 32430 6222 32430 6222 0 _037_
rlabel metal1 33074 5338 33074 5338 0 _038_
rlabel metal2 35098 6154 35098 6154 0 _039_
rlabel metal2 40802 2550 40802 2550 0 _040_
rlabel metal1 23828 4114 23828 4114 0 _041_
rlabel metal1 16422 4658 16422 4658 0 _042_
rlabel metal1 20838 8058 20838 8058 0 _043_
rlabel via2 32246 8619 32246 8619 0 _044_
rlabel metal2 14674 6460 14674 6460 0 _045_
rlabel metal1 19826 10438 19826 10438 0 _046_
rlabel metal1 19780 10506 19780 10506 0 _047_
rlabel metal1 26588 10642 26588 10642 0 _048_
rlabel metal1 22632 9486 22632 9486 0 _049_
rlabel metal2 21390 5185 21390 5185 0 _050_
rlabel metal2 22816 3978 22816 3978 0 _051_
rlabel metal1 18078 3978 18078 3978 0 _052_
rlabel metal1 35696 2482 35696 2482 0 _053_
rlabel metal1 39008 5542 39008 5542 0 _054_
rlabel metal2 21666 7650 21666 7650 0 _055_
rlabel metal1 20746 7344 20746 7344 0 _056_
rlabel metal2 21206 10353 21206 10353 0 _057_
rlabel metal1 21620 6086 21620 6086 0 _058_
rlabel metal1 22816 8942 22816 8942 0 _059_
rlabel metal1 23138 8942 23138 8942 0 _060_
rlabel metal1 20608 5542 20608 5542 0 _061_
rlabel metal2 22310 6222 22310 6222 0 _062_
rlabel metal2 20194 6630 20194 6630 0 _063_
rlabel metal1 23276 2618 23276 2618 0 _064_
rlabel metal1 26036 11526 26036 11526 0 _065_
rlabel metal1 24932 2822 24932 2822 0 _066_
rlabel metal2 24794 5627 24794 5627 0 _067_
rlabel metal2 25806 8092 25806 8092 0 _068_
rlabel metal1 25254 8058 25254 8058 0 _069_
rlabel metal1 27876 8466 27876 8466 0 _070_
rlabel metal1 28290 8466 28290 8466 0 _071_
rlabel metal1 27462 6358 27462 6358 0 _072_
rlabel metal2 35098 7072 35098 7072 0 _073_
rlabel metal1 27278 2618 27278 2618 0 _074_
rlabel metal2 30682 7514 30682 7514 0 _075_
rlabel metal1 32154 7480 32154 7480 0 _076_
rlabel metal1 33718 11730 33718 11730 0 _077_
rlabel metal2 27462 5763 27462 5763 0 _078_
rlabel metal2 30498 6596 30498 6596 0 _079_
rlabel metal1 29440 7922 29440 7922 0 _080_
rlabel metal1 32430 7276 32430 7276 0 _081_
rlabel metal1 32568 7378 32568 7378 0 _082_
rlabel metal1 33212 5270 33212 5270 0 _083_
rlabel metal2 35650 9690 35650 9690 0 _084_
rlabel metal1 33074 5236 33074 5236 0 _085_
rlabel metal1 35144 11050 35144 11050 0 _086_
rlabel metal2 36110 3264 36110 3264 0 _087_
rlabel metal1 39560 4454 39560 4454 0 _088_
rlabel metal2 37582 4352 37582 4352 0 _089_
rlabel metal2 36110 5491 36110 5491 0 _090_
rlabel metal1 35052 2482 35052 2482 0 _091_
rlabel metal1 36018 2618 36018 2618 0 _092_
rlabel metal4 32844 5372 32844 5372 0 _093_
rlabel via2 34454 5797 34454 5797 0 _094_
rlabel metal2 30958 6443 30958 6443 0 _095_
rlabel metal2 35466 6426 35466 6426 0 _096_
rlabel metal1 37306 5100 37306 5100 0 _097_
rlabel metal2 32890 5202 32890 5202 0 _098_
rlabel metal1 25392 5270 25392 5270 0 clknet_0_HCLK
rlabel metal2 13110 3196 13110 3196 0 clknet_2_0__leaf_HCLK
rlabel metal1 22264 7922 22264 7922 0 clknet_2_1__leaf_HCLK
rlabel metal1 38410 3094 38410 3094 0 clknet_2_2__leaf_HCLK
rlabel metal1 33856 5882 33856 5882 0 clknet_2_3__leaf_HCLK
rlabel metal1 59846 36754 59846 36754 0 gpio_oeb[0]
rlabel metal1 23138 37162 23138 37162 0 gpio_oeb[10]
rlabel metal1 19182 37230 19182 37230 0 gpio_oeb[11]
rlabel metal1 15594 37162 15594 37162 0 gpio_oeb[12]
rlabel metal1 11408 37230 11408 37230 0 gpio_oeb[13]
rlabel metal1 8372 37230 8372 37230 0 gpio_oeb[14]
rlabel metal1 4232 36822 4232 36822 0 gpio_oeb[15]
rlabel metal1 56442 37162 56442 37162 0 gpio_oeb[1]
rlabel metal1 52532 37230 52532 37230 0 gpio_oeb[2]
rlabel metal1 48806 37162 48806 37162 0 gpio_oeb[3]
rlabel metal1 44942 36686 44942 36686 0 gpio_oeb[4]
rlabel metal1 41492 37230 41492 37230 0 gpio_oeb[5]
rlabel metal1 37398 37230 37398 37230 0 gpio_oeb[6]
rlabel metal1 33810 37298 33810 37298 0 gpio_oeb[7]
rlabel metal1 30406 36754 30406 36754 0 gpio_oeb[8]
rlabel metal2 26174 38192 26174 38192 0 gpio_oeb[9]
rlabel metal1 58604 37162 58604 37162 0 gpio_out[0]
rlabel metal1 20792 37230 20792 37230 0 gpio_out[10]
rlabel metal1 17480 36822 17480 36822 0 gpio_out[11]
rlabel metal1 13432 37298 13432 37298 0 gpio_out[12]
rlabel metal1 9752 36822 9752 36822 0 gpio_out[13]
rlabel metal2 5934 38226 5934 38226 0 gpio_out[14]
rlabel metal1 2392 37298 2392 37298 0 gpio_out[15]
rlabel metal1 54280 37162 54280 37162 0 gpio_out[1]
rlabel metal1 50370 36686 50370 36686 0 gpio_out[2]
rlabel metal1 46920 37162 46920 37162 0 gpio_out[3]
rlabel metal1 43516 37162 43516 37162 0 gpio_out[4]
rlabel metal1 39330 37298 39330 37298 0 gpio_out[5]
rlabel metal2 35374 37954 35374 37954 0 gpio_out[6]
rlabel metal1 31740 37230 31740 37230 0 gpio_out[7]
rlabel metal1 28152 37230 28152 37230 0 gpio_out[8]
rlabel metal1 24472 36822 24472 36822 0 gpio_out[9]
rlabel metal2 9154 4420 9154 4420 0 last_HADDR\[0\]
rlabel metal1 33580 2890 33580 2890 0 last_HADDR\[10\]
rlabel metal1 36340 4250 36340 4250 0 last_HADDR\[11\]
rlabel metal2 40434 5406 40434 5406 0 last_HADDR\[12\]
rlabel metal1 41216 2414 41216 2414 0 last_HADDR\[13\]
rlabel metal2 42550 4182 42550 4182 0 last_HADDR\[14\]
rlabel metal1 45218 3162 45218 3162 0 last_HADDR\[15\]
rlabel metal2 9154 3434 9154 3434 0 last_HADDR\[1\]
rlabel metal2 18446 6698 18446 6698 0 last_HADDR\[2\]
rlabel metal1 20654 4114 20654 4114 0 last_HADDR\[3\]
rlabel metal1 16974 4998 16974 4998 0 last_HADDR\[4\]
rlabel metal1 25990 3434 25990 3434 0 last_HADDR\[5\]
rlabel metal1 27968 4454 27968 4454 0 last_HADDR\[6\]
rlabel metal1 16698 5100 16698 5100 0 last_HADDR\[7\]
rlabel via1 31786 4539 31786 4539 0 last_HADDR\[8\]
rlabel metal1 34040 3706 34040 3706 0 last_HADDR\[9\]
rlabel metal1 14122 7310 14122 7310 0 last_HSEL
rlabel metal1 15410 3502 15410 3502 0 last_HTRANS\[1\]
rlabel metal1 13294 2414 13294 2414 0 last_HWRITE
rlabel metal1 7314 2312 7314 2312 0 net1
rlabel metal2 17434 8772 17434 8772 0 net10
rlabel via2 37766 4029 37766 4029 0 net100
rlabel metal4 20148 8160 20148 8160 0 net101
rlabel metal1 21758 10676 21758 10676 0 net102
rlabel metal1 26588 4590 26588 4590 0 net1020
rlabel metal2 17894 4981 17894 4981 0 net103
rlabel metal2 7774 4930 7774 4930 0 net104
rlabel metal1 13524 5134 13524 5134 0 net1040
rlabel metal1 18308 10574 18308 10574 0 net1041
rlabel metal1 28658 5644 28658 5644 0 net105
rlabel metal1 19274 36720 19274 36720 0 net106
rlabel metal1 44390 36652 44390 36652 0 net107
rlabel metal2 21390 7242 21390 7242 0 net108
rlabel metal1 23414 2985 23414 2985 0 net109
rlabel metal1 16100 6290 16100 6290 0 net11
rlabel metal1 30314 11662 30314 11662 0 net110
rlabel metal1 12972 3162 12972 3162 0 net111
rlabel metal1 18906 6120 18906 6120 0 net112
rlabel metal1 10902 2346 10902 2346 0 net113
rlabel metal1 29762 11526 29762 11526 0 net114
rlabel metal2 49634 1656 49634 1656 0 net115
rlabel metal2 55430 1588 55430 1588 0 net116
rlabel metal2 59294 1792 59294 1792 0 net117
rlabel metal2 63158 1588 63158 1588 0 net118
rlabel metal2 72818 1622 72818 1622 0 net119
rlabel metal2 14858 3944 14858 3944 0 net12
rlabel metal1 10212 6630 10212 6630 0 net120
rlabel metal2 33166 9673 33166 9673 0 net121
rlabel metal1 18768 7922 18768 7922 0 net1218
rlabel metal2 16698 7582 16698 7582 0 net1219
rlabel metal1 22632 3162 22632 3162 0 net122
rlabel metal1 15088 4658 15088 4658 0 net1220
rlabel metal1 17296 6970 17296 6970 0 net1221
rlabel metal1 32660 3434 32660 3434 0 net123
rlabel metal1 12903 4658 12903 4658 0 net124
rlabel metal1 10350 3570 10350 3570 0 net125
rlabel metal1 15272 4454 15272 4454 0 net126
rlabel metal1 36432 10030 36432 10030 0 net127
rlabel metal2 34730 7259 34730 7259 0 net128
rlabel metal2 35650 3672 35650 3672 0 net129
rlabel metal2 17618 3587 17618 3587 0 net13
rlabel metal1 4784 2482 4784 2482 0 net130
rlabel metal1 11546 2618 11546 2618 0 net131
rlabel metal1 18170 3094 18170 3094 0 net132
rlabel metal1 47288 2618 47288 2618 0 net133
rlabel metal1 45402 2516 45402 2516 0 net134
rlabel metal1 41952 2958 41952 2958 0 net135
rlabel metal3 37283 9044 37283 9044 0 net136
rlabel metal1 39100 8398 39100 8398 0 net137
rlabel metal1 35190 2822 35190 2822 0 net138
rlabel metal1 50048 3434 50048 3434 0 net139
rlabel metal1 18446 6834 18446 6834 0 net1398
rlabel metal1 18584 7310 18584 7310 0 net1399
rlabel metal1 21896 5338 21896 5338 0 net14
rlabel metal1 47104 3706 47104 3706 0 net140
rlabel metal2 20286 8908 20286 8908 0 net1400
rlabel metal1 44261 3706 44261 3706 0 net141
rlabel metal2 3266 5644 3266 5644 0 net142
rlabel metal1 14582 7412 14582 7412 0 net143
rlabel metal1 13662 3672 13662 3672 0 net144
rlabel metal2 29302 8993 29302 8993 0 net145
rlabel metal1 24748 6834 24748 6834 0 net146
rlabel metal2 30038 6494 30038 6494 0 net147
rlabel metal2 12006 4641 12006 4641 0 net148
rlabel metal1 13294 4182 13294 4182 0 net149
rlabel via2 21114 2261 21114 2261 0 net15
rlabel metal2 24518 3893 24518 3893 0 net150
rlabel metal1 26864 9554 26864 9554 0 net151
rlabel metal1 26450 8908 26450 8908 0 net152
rlabel metal1 27140 3434 27140 3434 0 net153
rlabel metal2 30130 9537 30130 9537 0 net154
rlabel metal1 32292 10030 32292 10030 0 net155
rlabel metal1 32384 3094 32384 3094 0 net156
rlabel metal2 15410 5253 15410 5253 0 net157
rlabel metal1 19642 8500 19642 8500 0 net1578
rlabel metal1 15042 5270 15042 5270 0 net1579
rlabel via2 8234 3179 8234 3179 0 net158
rlabel metal1 19964 2958 19964 2958 0 net159
rlabel via3 34293 9724 34293 9724 0 net16
rlabel metal1 50140 2958 50140 2958 0 net160
rlabel metal1 46276 4794 46276 4794 0 net161
rlabel metal1 43700 3094 43700 3094 0 net162
rlabel metal2 40158 6205 40158 6205 0 net163
rlabel metal2 46506 5984 46506 5984 0 net164
rlabel metal2 38686 3774 38686 3774 0 net165
rlabel metal1 3358 2414 3358 2414 0 net166
rlabel metal2 14122 7106 14122 7106 0 net167
rlabel metal1 12282 2992 12282 2992 0 net168
rlabel metal2 6394 5474 6394 5474 0 net169
rlabel metal1 6302 3162 6302 3162 0 net17
rlabel metal1 8740 5338 8740 5338 0 net170
rlabel metal1 7084 3502 7084 3502 0 net171
rlabel metal2 11914 5831 11914 5831 0 net172
rlabel metal2 10626 7412 10626 7412 0 net173
rlabel metal2 13478 6528 13478 6528 0 net174
rlabel metal1 18078 6222 18078 6222 0 net175
rlabel metal2 19964 5542 19964 5542 0 net176
rlabel metal1 24518 6698 24518 6698 0 net177
rlabel metal2 17894 5882 17894 5882 0 net178
rlabel metal1 27094 8500 27094 8500 0 net179
rlabel metal2 8326 4828 8326 4828 0 net18
rlabel metal1 26808 6970 26808 6970 0 net180
rlabel metal2 10902 4284 10902 4284 0 net181
rlabel metal1 17572 6426 17572 6426 0 net182
rlabel metal1 24334 4046 24334 4046 0 net183
rlabel metal1 47058 3570 47058 3570 0 net184
rlabel metal1 35098 4590 35098 4590 0 net185
rlabel metal1 38042 4658 38042 4658 0 net186
rlabel metal1 17112 4182 17112 4182 0 net187
rlabel metal1 32568 6154 32568 6154 0 net188
rlabel metal2 32430 8092 32430 8092 0 net189
rlabel metal2 15318 7361 15318 7361 0 net19
rlabel metal1 22172 4046 22172 4046 0 net190
rlabel metal1 36018 6290 36018 6290 0 net191
rlabel metal1 35328 8058 35328 8058 0 net192
rlabel metal1 25990 11118 25990 11118 0 net193
rlabel metal2 29486 8908 29486 8908 0 net194
rlabel metal1 29762 8058 29762 8058 0 net195
rlabel metal1 7038 2618 7038 2618 0 net196
rlabel metal1 18124 6630 18124 6630 0 net197
rlabel metal2 24242 8670 24242 8670 0 net198
rlabel metal2 9154 6324 9154 6324 0 net199
rlabel metal2 34914 8313 34914 8313 0 net2
rlabel metal1 16238 7786 16238 7786 0 net20
rlabel metal1 15088 6426 15088 6426 0 net200
rlabel metal2 19274 9299 19274 9299 0 net201
rlabel metal2 7130 4114 7130 4114 0 net202
rlabel metal2 20378 8517 20378 8517 0 net203
rlabel metal1 22448 7786 22448 7786 0 net204
rlabel metal1 48300 3570 48300 3570 0 net205
rlabel metal1 43240 4794 43240 4794 0 net206
rlabel metal1 38272 6358 38272 6358 0 net207
rlabel via2 15778 3893 15778 3893 0 net208
rlabel metal1 28980 7786 28980 7786 0 net209
rlabel metal1 29670 2618 29670 2618 0 net21
rlabel metal1 25852 5746 25852 5746 0 net210
rlabel metal1 30314 5270 30314 5270 0 net211
rlabel metal1 48990 4250 48990 4250 0 net212
rlabel metal2 38686 7378 38686 7378 0 net213
rlabel metal2 30406 4862 30406 4862 0 net214
rlabel metal1 32706 5746 32706 5746 0 net215
rlabel metal2 31142 9741 31142 9741 0 net216
rlabel metal2 25162 5950 25162 5950 0 net217
rlabel metal1 28888 7310 28888 7310 0 net218
rlabel metal1 29440 7446 29440 7446 0 net219
rlabel metal1 37536 3910 37536 3910 0 net22
rlabel metal2 50830 3332 50830 3332 0 net220
rlabel metal1 39238 5100 39238 5100 0 net221
rlabel metal1 35972 5270 35972 5270 0 net222
rlabel metal1 37851 6970 37851 6970 0 net223
rlabel metal1 8648 5202 8648 5202 0 net224
rlabel metal2 15318 7684 15318 7684 0 net225
rlabel metal1 13800 6290 13800 6290 0 net226
rlabel metal1 21160 6290 21160 6290 0 net227
rlabel metal2 21022 9894 21022 9894 0 net228
rlabel metal1 14904 5202 14904 5202 0 net229
rlabel metal1 40158 3944 40158 3944 0 net23
rlabel metal1 14444 4114 14444 4114 0 net230
rlabel metal1 14536 2414 14536 2414 0 net231
rlabel metal2 39790 8636 39790 8636 0 net232
rlabel metal1 40342 4692 40342 4692 0 net233
rlabel metal1 37352 6834 37352 6834 0 net234
rlabel metal2 35926 7650 35926 7650 0 net235
rlabel via2 20838 9877 20838 9877 0 net236
rlabel metal1 15410 6222 15410 6222 0 net237
rlabel metal1 18814 5542 18814 5542 0 net238
rlabel metal2 36294 4301 36294 4301 0 net239
rlabel metal1 43470 2278 43470 2278 0 net24
rlabel metal2 45218 3230 45218 3230 0 net240
rlabel metal2 16698 5440 16698 5440 0 net241
rlabel metal2 19550 4301 19550 4301 0 net242
rlabel metal2 29670 4930 29670 4930 0 net243
rlabel metal1 20608 4658 20608 4658 0 net244
rlabel metal1 18446 5134 18446 5134 0 net245
rlabel metal2 23874 6647 23874 6647 0 net246
rlabel metal2 30222 8942 30222 8942 0 net247
rlabel metal1 30360 2414 30360 2414 0 net248
rlabel metal2 29578 7888 29578 7888 0 net249
rlabel metal1 47886 2278 47886 2278 0 net25
rlabel metal1 26312 7514 26312 7514 0 net250
rlabel metal2 29118 3774 29118 3774 0 net251
rlabel metal2 36938 5916 36938 5916 0 net252
rlabel metal2 39146 5610 39146 5610 0 net253
rlabel metal2 38594 3842 38594 3842 0 net254
rlabel metal2 28658 9316 28658 9316 0 net255
rlabel metal1 15456 4726 15456 4726 0 net256
rlabel metal2 26910 3536 26910 3536 0 net257
rlabel metal1 35328 5202 35328 5202 0 net258
rlabel metal1 35466 9418 35466 9418 0 net259
rlabel metal1 47794 4012 47794 4012 0 net26
rlabel metal1 36892 2414 36892 2414 0 net260
rlabel metal2 22034 8092 22034 8092 0 net261
rlabel metal2 18998 7140 18998 7140 0 net262
rlabel metal1 22862 3434 22862 3434 0 net263
rlabel metal2 33258 7514 33258 7514 0 net264
rlabel metal1 33948 9554 33948 9554 0 net265
rlabel metal2 35282 3230 35282 3230 0 net266
rlabel metal2 22586 6188 22586 6188 0 net267
rlabel via1 11546 4131 11546 4131 0 net268
rlabel metal1 18998 3672 18998 3672 0 net269
rlabel metal3 19757 8364 19757 8364 0 net27
rlabel metal1 41492 5678 41492 5678 0 net270
rlabel metal2 41998 4250 41998 4250 0 net271
rlabel metal1 43194 2414 43194 2414 0 net272
rlabel metal1 41147 4658 41147 4658 0 net273
rlabel metal2 40618 5338 40618 5338 0 net274
rlabel metal2 39422 2924 39422 2924 0 net275
rlabel metal2 19182 6103 19182 6103 0 net276
rlabel metal2 18906 8772 18906 8772 0 net277
rlabel metal1 19734 2482 19734 2482 0 net278
rlabel metal1 40388 5134 40388 5134 0 net279
rlabel metal1 14490 5678 14490 5678 0 net28
rlabel metal1 45908 2414 45908 2414 0 net280
rlabel metal2 46782 2754 46782 2754 0 net281
rlabel metal2 21298 8534 21298 8534 0 net282
rlabel metal3 15295 7004 15295 7004 0 net283
rlabel metal1 17204 2482 17204 2482 0 net284
rlabel metal1 27462 4182 27462 4182 0 net285
rlabel metal2 69506 3740 69506 3740 0 net289
rlabel metal1 22862 10098 22862 10098 0 net29
rlabel metal2 77050 3808 77050 3808 0 net290
rlabel metal4 33396 5848 33396 5848 0 net291
rlabel metal1 58144 3502 58144 3502 0 net293
rlabel metal1 62100 3502 62100 3502 0 net295
rlabel metal1 77326 2924 77326 2924 0 net296
rlabel metal1 76590 2482 76590 2482 0 net297
rlabel metal1 7314 4250 7314 4250 0 net298
rlabel metal1 9384 4794 9384 4794 0 net299
rlabel metal2 33258 2074 33258 2074 0 net3
rlabel metal1 17480 5338 17480 5338 0 net30
rlabel metal2 12650 3145 12650 3145 0 net300
rlabel metal2 6486 4284 6486 4284 0 net301
rlabel metal2 28106 4828 28106 4828 0 net302
rlabel metal1 67620 3502 67620 3502 0 net304
rlabel metal2 54050 3740 54050 3740 0 net306
rlabel metal1 57178 3060 57178 3060 0 net307
rlabel metal1 58788 3162 58788 3162 0 net308
rlabel metal1 58512 2482 58512 2482 0 net309
rlabel metal1 27416 8942 27416 8942 0 net31
rlabel metal2 27922 4488 27922 4488 0 net310
rlabel metal1 52164 3502 52164 3502 0 net312
rlabel metal1 72404 3502 72404 3502 0 net314
rlabel metal2 65458 3604 65458 3604 0 net316
rlabel metal2 65550 2754 65550 2754 0 net317
rlabel metal4 17940 6460 17940 6460 0 net318
rlabel metal1 65412 3502 65412 3502 0 net319
rlabel metal1 20332 4250 20332 4250 0 net32
rlabel metal2 53222 3876 53222 3876 0 net324
rlabel metal2 52118 2754 52118 2754 0 net325
rlabel metal2 14306 6188 14306 6188 0 net326
rlabel metal1 20102 2482 20102 2482 0 net33
rlabel metal2 56074 3196 56074 3196 0 net332
rlabel metal2 54050 2754 54050 2754 0 net333
rlabel metal2 41262 3706 41262 3706 0 net334
rlabel metal1 25530 3162 25530 3162 0 net34
rlabel metal2 68678 3876 68678 3876 0 net340
rlabel metal2 67666 2754 67666 2754 0 net341
rlabel metal1 40986 3536 40986 3536 0 net342
rlabel metal1 62560 3162 62560 3162 0 net348
rlabel metal2 61778 2754 61778 2754 0 net349
rlabel metal2 32062 4318 32062 4318 0 net35
rlabel metal2 12742 6528 12742 6528 0 net350
rlabel metal2 23414 4063 23414 4063 0 net351
rlabel metal2 71530 3196 71530 3196 0 net357
rlabel metal2 69506 2754 69506 2754 0 net358
rlabel metal2 41538 5168 41538 5168 0 net359
rlabel metal1 13018 5338 13018 5338 0 net36
rlabel metal2 73738 3740 73738 3740 0 net365
rlabel metal2 72634 2754 72634 2754 0 net366
rlabel metal1 4370 2924 4370 2924 0 net367
rlabel metal1 14950 9690 14950 9690 0 net368
rlabel metal1 18262 2448 18262 2448 0 net369
rlabel metal2 14858 7038 14858 7038 0 net37
rlabel metal2 10810 4437 10810 4437 0 net370
rlabel metal2 41078 4012 41078 4012 0 net371
rlabel metal1 35926 3536 35926 3536 0 net377
rlabel metal1 49634 4454 49634 4454 0 net378
rlabel metal1 49634 2482 49634 2482 0 net379
rlabel metal2 31970 6035 31970 6035 0 net38
rlabel metal1 32706 5882 32706 5882 0 net380
rlabel metal2 36938 7837 36938 7837 0 net381
rlabel metal1 24380 5882 24380 5882 0 net382
rlabel metal1 31901 10642 31901 10642 0 net383
rlabel metal2 30958 3995 30958 3995 0 net384
rlabel metal2 18906 3298 18906 3298 0 net385
rlabel metal1 18768 7514 18768 7514 0 net386
rlabel metal2 30314 7344 30314 7344 0 net387
rlabel metal3 27531 11084 27531 11084 0 net388
rlabel metal1 23092 5678 23092 5678 0 net389
rlabel metal1 37260 6426 37260 6426 0 net39
rlabel metal2 31694 3893 31694 3893 0 net390
rlabel metal2 3818 3604 3818 3604 0 net391
rlabel metal2 12466 5916 12466 5916 0 net392
rlabel metal1 8786 5134 8786 5134 0 net393
rlabel metal2 12650 2176 12650 2176 0 net394
rlabel metal1 8418 3502 8418 3502 0 net395
rlabel metal1 12006 3570 12006 3570 0 net396
rlabel metal1 24242 6766 24242 6766 0 net397
rlabel metal1 21068 3706 21068 3706 0 net398
rlabel metal2 16606 5865 16606 5865 0 net399
rlabel metal1 35834 2550 35834 2550 0 net4
rlabel metal1 36202 3502 36202 3502 0 net40
rlabel metal1 25392 10438 25392 10438 0 net400
rlabel metal1 16330 3910 16330 3910 0 net401
rlabel metal1 29026 6834 29026 6834 0 net402
rlabel metal1 29256 9146 29256 9146 0 net403
rlabel metal1 18170 4454 18170 4454 0 net404
rlabel metal1 28704 4114 28704 4114 0 net405
rlabel metal2 27370 8704 27370 8704 0 net406
rlabel metal1 27968 9554 27968 9554 0 net407
rlabel via2 13570 4675 13570 4675 0 net408
rlabel metal3 17940 4420 17940 4420 0 net409
rlabel metal1 42918 6222 42918 6222 0 net41
rlabel metal1 39192 7310 39192 7310 0 net410
rlabel metal2 35190 5814 35190 5814 0 net411
rlabel metal1 23828 8466 23828 8466 0 net412
rlabel metal1 18906 7888 18906 7888 0 net413
rlabel metal1 17940 5814 17940 5814 0 net414
rlabel metal1 22195 3502 22195 3502 0 net415
rlabel metal2 36570 7004 36570 7004 0 net416
rlabel metal1 33350 5066 33350 5066 0 net417
rlabel metal1 28336 5134 28336 5134 0 net418
rlabel metal1 36800 3502 36800 3502 0 net419
rlabel metal2 33258 4318 33258 4318 0 net42
rlabel metal1 34316 7514 34316 7514 0 net420
rlabel metal1 30406 3060 30406 3060 0 net421
rlabel metal1 34868 9690 34868 9690 0 net422
rlabel metal2 34086 6732 34086 6732 0 net423
rlabel metal1 40940 6222 40940 6222 0 net424
rlabel metal1 42136 5338 42136 5338 0 net425
rlabel metal1 37260 4726 37260 4726 0 net426
rlabel metal2 41354 4471 41354 4471 0 net427
rlabel metal1 19964 6290 19964 6290 0 net428
rlabel metal2 18170 5865 18170 5865 0 net429
rlabel metal2 42734 4811 42734 4811 0 net43
rlabel via2 18170 8347 18170 8347 0 net430
rlabel metal1 19918 8806 19918 8806 0 net431
rlabel metal1 40204 5678 40204 5678 0 net432
rlabel metal2 34178 4318 34178 4318 0 net433
rlabel metal2 21206 7684 21206 7684 0 net434
rlabel metal2 10442 7293 10442 7293 0 net435
rlabel metal2 16606 7718 16606 7718 0 net436
rlabel metal1 15318 2482 15318 2482 0 net437
rlabel metal2 34822 9401 34822 9401 0 net438
rlabel metal1 23000 3026 23000 3026 0 net439
rlabel metal2 48346 4454 48346 4454 0 net44
rlabel metal1 21896 3026 21896 3026 0 net440
rlabel metal2 30866 3264 30866 3264 0 net441
rlabel metal2 12834 4828 12834 4828 0 net444
rlabel metal4 14260 7412 14260 7412 0 net445
rlabel metal2 12282 4199 12282 4199 0 net446
rlabel metal2 10994 3417 10994 3417 0 net447
rlabel metal1 52394 3162 52394 3162 0 net45
rlabel metal2 21482 6239 21482 6239 0 net450
rlabel metal2 21666 5372 21666 5372 0 net451
rlabel metal2 29578 10268 29578 10268 0 net452
rlabel metal1 30084 4046 30084 4046 0 net453
rlabel metal1 25438 5202 25438 5202 0 net456
rlabel via2 35926 9877 35926 9877 0 net457
rlabel metal1 36064 9486 36064 9486 0 net458
rlabel metal2 35190 3774 35190 3774 0 net459
rlabel metal2 53866 3604 53866 3604 0 net46
rlabel metal2 40066 8500 40066 8500 0 net462
rlabel metal1 32407 2414 32407 2414 0 net463
rlabel metal2 37398 5304 37398 5304 0 net464
rlabel metal1 37168 4114 37168 4114 0 net465
rlabel metal1 14467 8942 14467 8942 0 net468
rlabel metal1 3864 2618 3864 2618 0 net469
rlabel metal1 10074 4114 10074 4114 0 net47
rlabel metal1 8050 2482 8050 2482 0 net470
rlabel metal1 17066 2414 17066 2414 0 net471
rlabel metal2 48898 4828 48898 4828 0 net474
rlabel metal1 49726 3366 49726 3366 0 net475
rlabel metal2 47978 4284 47978 4284 0 net476
rlabel metal1 43838 4046 43838 4046 0 net477
rlabel metal2 57362 3298 57362 3298 0 net48
rlabel metal2 4002 5406 4002 5406 0 net480
rlabel metal3 19711 9724 19711 9724 0 net481
rlabel metal3 18377 8772 18377 8772 0 net482
rlabel metal1 19872 4522 19872 4522 0 net483
rlabel metal2 8602 2689 8602 2689 0 net486
rlabel metal2 12650 8194 12650 8194 0 net487
rlabel viali 12742 4113 12742 4113 0 net488
rlabel metal1 23966 4590 23966 4590 0 net489
rlabel metal2 60950 3298 60950 3298 0 net49
rlabel metal2 47978 2244 47978 2244 0 net492
rlabel metal2 42274 3298 42274 3298 0 net493
rlabel metal1 39054 2482 39054 2482 0 net494
rlabel metal1 43125 2482 43125 2482 0 net495
rlabel metal2 41446 8126 41446 8126 0 net498
rlabel metal2 38410 2176 38410 2176 0 net499
rlabel metal2 42090 3604 42090 3604 0 net5
rlabel metal2 64538 3332 64538 3332 0 net50
rlabel metal1 33902 4114 33902 4114 0 net500
rlabel metal2 40526 3859 40526 3859 0 net501
rlabel metal1 28106 10778 28106 10778 0 net504
rlabel metal1 27738 9622 27738 9622 0 net505
rlabel metal1 17388 3162 17388 3162 0 net506
rlabel metal1 28290 4658 28290 4658 0 net507
rlabel metal1 67850 3162 67850 3162 0 net51
rlabel metal1 30176 9554 30176 9554 0 net510
rlabel metal1 21390 2414 21390 2414 0 net511
rlabel metal1 24518 5780 24518 5780 0 net512
rlabel metal2 31878 7276 31878 7276 0 net513
rlabel metal2 11546 6018 11546 6018 0 net516
rlabel via2 20470 10013 20470 10013 0 net517
rlabel metal2 7590 5134 7590 5134 0 net518
rlabel via2 21390 4029 21390 4029 0 net519
rlabel metal2 69322 3604 69322 3604 0 net52
rlabel metal1 6716 3570 6716 3570 0 net522
rlabel metal1 6670 2414 6670 2414 0 net523
rlabel metal2 5658 4556 5658 4556 0 net524
rlabel metal1 14398 3502 14398 3502 0 net525
rlabel metal2 47058 5372 47058 5372 0 net528
rlabel metal1 48346 3060 48346 3060 0 net529
rlabel metal1 71944 2618 71944 2618 0 net53
rlabel metal2 47242 4828 47242 4828 0 net530
rlabel metal1 42872 3162 42872 3162 0 net531
rlabel metal2 76958 4964 76958 4964 0 net536
rlabel metal2 75486 2958 75486 2958 0 net537
rlabel metal1 11270 5814 11270 5814 0 net538
rlabel metal1 18400 7990 18400 7990 0 net539
rlabel metal1 9154 3026 9154 3026 0 net54
rlabel metal2 15962 8262 15962 8262 0 net540
rlabel metal1 15042 3366 15042 3366 0 net541
rlabel metal1 14398 6766 14398 6766 0 net542
rlabel metal1 8027 2890 8027 2890 0 net543
rlabel metal1 14122 5644 14122 5644 0 net544
rlabel metal2 11546 3553 11546 3553 0 net545
rlabel metal2 19642 7616 19642 7616 0 net546
rlabel metal2 24702 4981 24702 4981 0 net547
rlabel metal1 15410 5338 15410 5338 0 net548
rlabel metal1 17572 6222 17572 6222 0 net549
rlabel metal2 74474 3332 74474 3332 0 net55
rlabel metal1 15916 4590 15916 4590 0 net550
rlabel metal1 21206 6358 21206 6358 0 net551
rlabel viali 27002 10028 27002 10028 0 net552
rlabel metal1 20102 5848 20102 5848 0 net553
rlabel metal1 26404 9010 26404 9010 0 net554
rlabel metal1 27508 6426 27508 6426 0 net555
rlabel metal1 35190 2278 35190 2278 0 net556
rlabel metal1 45264 3638 45264 3638 0 net557
rlabel metal1 36478 4114 36478 4114 0 net558
rlabel metal1 36984 4454 36984 4454 0 net559
rlabel metal1 75302 4080 75302 4080 0 net56
rlabel metal1 13892 6222 13892 6222 0 net560
rlabel metal1 9108 3162 9108 3162 0 net561
rlabel metal1 16192 5882 16192 5882 0 net562
rlabel metal2 20838 8364 20838 8364 0 net563
rlabel metal3 27715 10812 27715 10812 0 net564
rlabel metal4 20700 7956 20700 7956 0 net565
rlabel metal1 22816 5338 22816 5338 0 net566
rlabel metal1 27876 7446 27876 7446 0 net567
rlabel metal2 17526 3417 17526 3417 0 net568
rlabel metal1 32292 3502 32292 3502 0 net569
rlabel metal1 15686 5780 15686 5780 0 net57
rlabel metal2 30314 5848 30314 5848 0 net570
rlabel metal1 33212 6834 33212 6834 0 net571
rlabel via2 36662 10013 36662 10013 0 net572
rlabel metal1 30682 2482 30682 2482 0 net573
rlabel metal1 29670 5338 29670 5338 0 net574
rlabel metal1 33350 5236 33350 5236 0 net575
rlabel metal1 9798 3570 9798 3570 0 net576
rlabel metal1 5980 2278 5980 2278 0 net577
rlabel metal2 18722 8976 18722 8976 0 net578
rlabel metal2 22586 8772 22586 8772 0 net579
rlabel metal1 21666 3366 21666 3366 0 net58
rlabel metal1 45724 4658 45724 4658 0 net580
rlabel metal1 45770 2482 45770 2482 0 net581
rlabel metal1 41952 3706 41952 3706 0 net582
rlabel metal1 36616 5202 36616 5202 0 net583
rlabel metal2 74566 3196 74566 3196 0 net586
rlabel metal2 76222 2618 76222 2618 0 net587
rlabel metal2 76682 2822 76682 2822 0 net588
rlabel metal2 15134 3825 15134 3825 0 net589
rlabel metal2 26634 10540 26634 10540 0 net59
rlabel metal1 32637 10506 32637 10506 0 net590
rlabel metal1 26864 5882 26864 5882 0 net591
rlabel metal1 21390 4250 21390 4250 0 net592
rlabel metal2 20286 3587 20286 3587 0 net593
rlabel metal1 21390 2618 21390 2618 0 net594
rlabel metal2 48530 4318 48530 4318 0 net595
rlabel metal1 48392 2414 48392 2414 0 net596
rlabel metal2 45678 4828 45678 4828 0 net597
rlabel metal1 39192 8942 39192 8942 0 net598
rlabel metal1 38502 4148 38502 4148 0 net599
rlabel metal2 45586 4420 45586 4420 0 net6
rlabel metal1 17480 4590 17480 4590 0 net60
rlabel metal1 33534 4794 33534 4794 0 net600
rlabel metal1 53130 3570 53130 3570 0 net604
rlabel metal2 52854 3162 52854 3162 0 net605
rlabel metal1 54648 3502 54648 3502 0 net609
rlabel metal1 29900 9010 29900 9010 0 net61
rlabel metal2 55338 2618 55338 2618 0 net610
rlabel metal2 57454 3196 57454 3196 0 net614
rlabel metal2 58650 2890 58650 2890 0 net615
rlabel metal2 64906 3196 64906 3196 0 net619
rlabel metal2 32522 8313 32522 8313 0 net62
rlabel metal2 66286 3162 66286 3162 0 net620
rlabel metal2 61134 3196 61134 3196 0 net624
rlabel metal2 62790 2890 62790 2890 0 net625
rlabel metal1 70104 3502 70104 3502 0 net629
rlabel metal1 34178 9452 34178 9452 0 net63
rlabel metal2 70518 2618 70518 2618 0 net630
rlabel metal1 68540 3570 68540 3570 0 net634
rlabel metal2 68310 3162 68310 3162 0 net635
rlabel metal2 71714 3876 71714 3876 0 net639
rlabel metal1 59018 36618 59018 36618 0 net64
rlabel metal1 73186 2414 73186 2414 0 net640
rlabel metal2 51382 3468 51382 3468 0 net641
rlabel metal1 48852 3706 48852 3706 0 net642
rlabel metal1 45586 4250 45586 4250 0 net643
rlabel metal2 8602 6052 8602 6052 0 net644
rlabel metal1 6210 3026 6210 3026 0 net645
rlabel metal1 6256 3706 6256 3706 0 net646
rlabel metal2 22494 37060 22494 37060 0 net65
rlabel metal2 44206 4624 44206 4624 0 net650
rlabel metal1 19228 7854 19228 7854 0 net651
rlabel metal1 16330 4794 16330 4794 0 net652
rlabel metal1 19228 9146 19228 9146 0 net653
rlabel metal2 21758 11237 21758 11237 0 net654
rlabel metal2 17342 2227 17342 2227 0 net655
rlabel metal2 35282 6188 35282 6188 0 net656
rlabel metal1 36938 4658 36938 4658 0 net657
rlabel metal1 44068 4658 44068 4658 0 net658
rlabel metal1 41584 4794 41584 4794 0 net659
rlabel metal1 18906 36890 18906 36890 0 net66
rlabel metal1 41630 6290 41630 6290 0 net660
rlabel metal2 41170 5916 41170 5916 0 net661
rlabel metal1 40848 5202 40848 5202 0 net662
rlabel metal2 39330 6188 39330 6188 0 net663
rlabel metal1 39744 5202 39744 5202 0 net664
rlabel metal1 39330 5100 39330 5100 0 net665
rlabel metal1 32016 5746 32016 5746 0 net666
rlabel metal1 32890 5168 32890 5168 0 net667
rlabel metal1 35190 6834 35190 6834 0 net668
rlabel metal1 32407 4114 32407 4114 0 net669
rlabel metal2 15134 37060 15134 37060 0 net67
rlabel metal2 77602 4148 77602 4148 0 net672
rlabel metal2 76682 4250 76682 4250 0 net673
rlabel metal2 74658 3366 74658 3366 0 net674
rlabel metal2 37306 7854 37306 7854 0 net675
rlabel metal2 25162 9724 25162 9724 0 net676
rlabel metal1 30590 6834 30590 6834 0 net677
rlabel metal1 25622 7922 25622 7922 0 net678
rlabel metal1 33764 7310 33764 7310 0 net679
rlabel metal2 11914 37060 11914 37060 0 net68
rlabel metal2 31786 8126 31786 8126 0 net680
rlabel metal1 26864 7922 26864 7922 0 net681
rlabel metal1 21902 7378 21902 7378 0 net682
rlabel metal1 24058 5678 24058 5678 0 net683
rlabel metal2 32706 8806 32706 8806 0 net684
rlabel metal2 7774 37060 7774 37060 0 net69
rlabel metal1 47564 3162 47564 3162 0 net7
rlabel metal2 11822 36686 11822 36686 0 net70
rlabel metal2 55614 37060 55614 37060 0 net71
rlabel metal2 51934 37060 51934 37060 0 net72
rlabel metal2 48254 37060 48254 37060 0 net73
rlabel metal1 44574 36686 44574 36686 0 net74
rlabel metal2 40894 37060 40894 37060 0 net75
rlabel metal2 37030 37060 37030 37060 0 net76
rlabel metal2 33810 37060 33810 37060 0 net77
rlabel metal1 29854 36686 29854 36686 0 net78
rlabel metal1 26128 36890 26128 36890 0 net79
rlabel metal2 13570 7072 13570 7072 0 net8
rlabel metal2 58834 25840 58834 25840 0 net80
rlabel metal2 21942 30702 21942 30702 0 net81
rlabel metal2 18814 31858 18814 31858 0 net82
rlabel via3 14605 36516 14605 36516 0 net83
rlabel metal2 10994 33167 10994 33167 0 net84
rlabel metal2 7130 34833 7130 34833 0 net85
rlabel metal2 20010 8262 20010 8262 0 net853
rlabel metal1 18768 7378 18768 7378 0 net854
rlabel metal2 38318 7548 38318 7548 0 net855
rlabel metal1 37306 6188 37306 6188 0 net856
rlabel metal2 35834 5406 35834 5406 0 net857
rlabel metal2 3542 30668 3542 30668 0 net86
rlabel metal1 39422 29614 39422 29614 0 net87
rlabel metal2 27140 16560 27140 16560 0 net88
rlabel metal2 26312 16560 26312 16560 0 net89
rlabel metal1 19366 9554 19366 9554 0 net9
rlabel metal2 43378 25874 43378 25874 0 net90
rlabel metal2 39146 29308 39146 29308 0 net91
rlabel metal1 26818 2448 26818 2448 0 net92
rlabel metal3 32131 36380 32131 36380 0 net93
rlabel metal1 29486 37196 29486 37196 0 net94
rlabel metal2 25806 36550 25806 36550 0 net95
rlabel metal1 22816 11322 22816 11322 0 net96
rlabel metal2 33442 5100 33442 5100 0 net97
rlabel metal1 34776 7446 34776 7446 0 net98
rlabel metal1 9614 5644 9614 5644 0 net99
<< properties >>
string FIXED_BBOX 0 0 80000 40000
<< end >>
