VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ahb_counter
  CLASS BLOCK ;
  FOREIGN ahb_counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 200.000 ;
  PIN HADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END HADDR[0]
  PIN HADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END HADDR[10]
  PIN HADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END HADDR[11]
  PIN HADDR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END HADDR[12]
  PIN HADDR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END HADDR[13]
  PIN HADDR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END HADDR[14]
  PIN HADDR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END HADDR[15]
  PIN HADDR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END HADDR[16]
  PIN HADDR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END HADDR[17]
  PIN HADDR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END HADDR[18]
  PIN HADDR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END HADDR[19]
  PIN HADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END HADDR[1]
  PIN HADDR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END HADDR[20]
  PIN HADDR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END HADDR[21]
  PIN HADDR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END HADDR[22]
  PIN HADDR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END HADDR[23]
  PIN HADDR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END HADDR[24]
  PIN HADDR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END HADDR[25]
  PIN HADDR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END HADDR[26]
  PIN HADDR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END HADDR[27]
  PIN HADDR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END HADDR[28]
  PIN HADDR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END HADDR[29]
  PIN HADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END HADDR[2]
  PIN HADDR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END HADDR[30]
  PIN HADDR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END HADDR[31]
  PIN HADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END HADDR[3]
  PIN HADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END HADDR[4]
  PIN HADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END HADDR[5]
  PIN HADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END HADDR[6]
  PIN HADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END HADDR[7]
  PIN HADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END HADDR[8]
  PIN HADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END HADDR[9]
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END HCLK
  PIN HRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END HRDATA[0]
  PIN HRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END HRDATA[10]
  PIN HRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END HRDATA[11]
  PIN HRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END HRDATA[12]
  PIN HRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END HRDATA[13]
  PIN HRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END HRDATA[14]
  PIN HRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END HRDATA[15]
  PIN HRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END HRDATA[16]
  PIN HRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END HRDATA[17]
  PIN HRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END HRDATA[18]
  PIN HRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END HRDATA[19]
  PIN HRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END HRDATA[1]
  PIN HRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END HRDATA[20]
  PIN HRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END HRDATA[21]
  PIN HRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END HRDATA[22]
  PIN HRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END HRDATA[23]
  PIN HRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END HRDATA[24]
  PIN HRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END HRDATA[25]
  PIN HRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END HRDATA[26]
  PIN HRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END HRDATA[27]
  PIN HRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END HRDATA[28]
  PIN HRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END HRDATA[29]
  PIN HRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END HRDATA[2]
  PIN HRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END HRDATA[30]
  PIN HRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END HRDATA[31]
  PIN HRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END HRDATA[3]
  PIN HRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END HRDATA[4]
  PIN HRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END HRDATA[5]
  PIN HRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END HRDATA[6]
  PIN HRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END HRDATA[7]
  PIN HRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END HRDATA[8]
  PIN HRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END HRDATA[9]
  PIN HREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END HREADY
  PIN HREADYOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END HREADYOUT
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END HRESETn
  PIN HSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END HSEL
  PIN HSIZE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END HSIZE[0]
  PIN HSIZE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END HSIZE[1]
  PIN HSIZE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END HSIZE[2]
  PIN HTRANS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END HTRANS[0]
  PIN HTRANS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END HTRANS[1]
  PIN HWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END HWDATA[0]
  PIN HWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END HWDATA[10]
  PIN HWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END HWDATA[11]
  PIN HWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END HWDATA[12]
  PIN HWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END HWDATA[13]
  PIN HWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END HWDATA[14]
  PIN HWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END HWDATA[15]
  PIN HWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END HWDATA[16]
  PIN HWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END HWDATA[17]
  PIN HWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END HWDATA[18]
  PIN HWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END HWDATA[19]
  PIN HWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END HWDATA[1]
  PIN HWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END HWDATA[20]
  PIN HWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END HWDATA[21]
  PIN HWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END HWDATA[22]
  PIN HWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END HWDATA[23]
  PIN HWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END HWDATA[24]
  PIN HWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END HWDATA[25]
  PIN HWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END HWDATA[26]
  PIN HWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END HWDATA[27]
  PIN HWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END HWDATA[28]
  PIN HWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END HWDATA[29]
  PIN HWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END HWDATA[2]
  PIN HWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END HWDATA[30]
  PIN HWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END HWDATA[31]
  PIN HWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END HWDATA[3]
  PIN HWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END HWDATA[4]
  PIN HWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END HWDATA[5]
  PIN HWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END HWDATA[6]
  PIN HWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END HWDATA[7]
  PIN HWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END HWDATA[8]
  PIN HWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END HWDATA[9]
  PIN HWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END HWRITE
  PIN gpio_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 296.330 196.000 296.610 200.000 ;
    END
  END gpio_oeb[0]
  PIN gpio_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 112.330 196.000 112.610 200.000 ;
    END
  END gpio_oeb[10]
  PIN gpio_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 93.930 196.000 94.210 200.000 ;
    END
  END gpio_oeb[11]
  PIN gpio_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 75.530 196.000 75.810 200.000 ;
    END
  END gpio_oeb[12]
  PIN gpio_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 57.130 196.000 57.410 200.000 ;
    END
  END gpio_oeb[13]
  PIN gpio_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 196.000 39.010 200.000 ;
    END
  END gpio_oeb[14]
  PIN gpio_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 20.330 196.000 20.610 200.000 ;
    END
  END gpio_oeb[15]
  PIN gpio_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 277.930 196.000 278.210 200.000 ;
    END
  END gpio_oeb[1]
  PIN gpio_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 259.530 196.000 259.810 200.000 ;
    END
  END gpio_oeb[2]
  PIN gpio_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 241.130 196.000 241.410 200.000 ;
    END
  END gpio_oeb[3]
  PIN gpio_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 222.730 196.000 223.010 200.000 ;
    END
  END gpio_oeb[4]
  PIN gpio_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 204.330 196.000 204.610 200.000 ;
    END
  END gpio_oeb[5]
  PIN gpio_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 185.930 196.000 186.210 200.000 ;
    END
  END gpio_oeb[6]
  PIN gpio_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 167.530 196.000 167.810 200.000 ;
    END
  END gpio_oeb[7]
  PIN gpio_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 149.130 196.000 149.410 200.000 ;
    END
  END gpio_oeb[8]
  PIN gpio_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 130.730 196.000 131.010 200.000 ;
    END
  END gpio_oeb[9]
  PIN gpio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 287.130 196.000 287.410 200.000 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 196.000 103.410 200.000 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 84.730 196.000 85.010 200.000 ;
    END
  END gpio_out[11]
  PIN gpio_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 66.330 196.000 66.610 200.000 ;
    END
  END gpio_out[12]
  PIN gpio_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 47.930 196.000 48.210 200.000 ;
    END
  END gpio_out[13]
  PIN gpio_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 29.530 196.000 29.810 200.000 ;
    END
  END gpio_out[14]
  PIN gpio_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 11.130 196.000 11.410 200.000 ;
    END
  END gpio_out[15]
  PIN gpio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 268.730 196.000 269.010 200.000 ;
    END
  END gpio_out[1]
  PIN gpio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 250.330 196.000 250.610 200.000 ;
    END
  END gpio_out[2]
  PIN gpio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 231.930 196.000 232.210 200.000 ;
    END
  END gpio_out[3]
  PIN gpio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 213.530 196.000 213.810 200.000 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 195.130 196.000 195.410 200.000 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 176.730 196.000 177.010 200.000 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 158.330 196.000 158.610 200.000 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 139.930 196.000 140.210 200.000 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 121.530 196.000 121.810 200.000 ;
    END
  END gpio_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.640 10.640 27.240 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 179.240 10.640 180.840 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.840 10.640 334.440 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.940 10.640 30.540 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 182.540 10.640 184.140 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 336.140 10.640 337.740 187.920 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 9.930 10.795 389.810 187.870 ;
      LAYER li1 ;
        RECT 10.120 10.795 389.620 187.765 ;
      LAYER met1 ;
        RECT 10.120 0.380 389.620 187.920 ;
      LAYER met2 ;
        RECT 11.690 195.720 20.050 196.000 ;
        RECT 20.890 195.720 29.250 196.000 ;
        RECT 30.090 195.720 38.450 196.000 ;
        RECT 39.290 195.720 47.650 196.000 ;
        RECT 48.490 195.720 56.850 196.000 ;
        RECT 57.690 195.720 66.050 196.000 ;
        RECT 66.890 195.720 75.250 196.000 ;
        RECT 76.090 195.720 84.450 196.000 ;
        RECT 85.290 195.720 93.650 196.000 ;
        RECT 94.490 195.720 102.850 196.000 ;
        RECT 103.690 195.720 112.050 196.000 ;
        RECT 112.890 195.720 121.250 196.000 ;
        RECT 122.090 195.720 130.450 196.000 ;
        RECT 131.290 195.720 139.650 196.000 ;
        RECT 140.490 195.720 148.850 196.000 ;
        RECT 149.690 195.720 158.050 196.000 ;
        RECT 158.890 195.720 167.250 196.000 ;
        RECT 168.090 195.720 176.450 196.000 ;
        RECT 177.290 195.720 185.650 196.000 ;
        RECT 186.490 195.720 194.850 196.000 ;
        RECT 195.690 195.720 204.050 196.000 ;
        RECT 204.890 195.720 213.250 196.000 ;
        RECT 214.090 195.720 222.450 196.000 ;
        RECT 223.290 195.720 231.650 196.000 ;
        RECT 232.490 195.720 240.850 196.000 ;
        RECT 241.690 195.720 250.050 196.000 ;
        RECT 250.890 195.720 259.250 196.000 ;
        RECT 260.090 195.720 268.450 196.000 ;
        RECT 269.290 195.720 277.650 196.000 ;
        RECT 278.490 195.720 286.850 196.000 ;
        RECT 287.690 195.720 296.050 196.000 ;
        RECT 296.890 195.720 388.140 196.000 ;
        RECT 11.140 4.280 388.140 195.720 ;
        RECT 11.140 0.350 44.890 4.280 ;
        RECT 45.730 0.350 48.110 4.280 ;
        RECT 48.950 0.350 51.330 4.280 ;
        RECT 52.170 0.350 54.550 4.280 ;
        RECT 55.390 0.350 57.770 4.280 ;
        RECT 58.610 0.350 60.990 4.280 ;
        RECT 61.830 0.350 64.210 4.280 ;
        RECT 65.050 0.350 67.430 4.280 ;
        RECT 68.270 0.350 70.650 4.280 ;
        RECT 71.490 0.350 73.870 4.280 ;
        RECT 74.710 0.350 77.090 4.280 ;
        RECT 77.930 0.350 80.310 4.280 ;
        RECT 81.150 0.350 83.530 4.280 ;
        RECT 84.370 0.350 86.750 4.280 ;
        RECT 87.590 0.350 89.970 4.280 ;
        RECT 90.810 0.350 93.190 4.280 ;
        RECT 94.030 0.350 96.410 4.280 ;
        RECT 97.250 0.350 99.630 4.280 ;
        RECT 100.470 0.350 102.850 4.280 ;
        RECT 103.690 0.350 106.070 4.280 ;
        RECT 106.910 0.350 109.290 4.280 ;
        RECT 110.130 0.350 112.510 4.280 ;
        RECT 113.350 0.350 115.730 4.280 ;
        RECT 116.570 0.350 118.950 4.280 ;
        RECT 119.790 0.350 122.170 4.280 ;
        RECT 123.010 0.350 125.390 4.280 ;
        RECT 126.230 0.350 128.610 4.280 ;
        RECT 129.450 0.350 131.830 4.280 ;
        RECT 132.670 0.350 135.050 4.280 ;
        RECT 135.890 0.350 138.270 4.280 ;
        RECT 139.110 0.350 141.490 4.280 ;
        RECT 142.330 0.350 144.710 4.280 ;
        RECT 145.550 0.350 147.930 4.280 ;
        RECT 148.770 0.350 151.150 4.280 ;
        RECT 151.990 0.350 154.370 4.280 ;
        RECT 155.210 0.350 157.590 4.280 ;
        RECT 158.430 0.350 160.810 4.280 ;
        RECT 161.650 0.350 164.030 4.280 ;
        RECT 164.870 0.350 167.250 4.280 ;
        RECT 168.090 0.350 170.470 4.280 ;
        RECT 171.310 0.350 173.690 4.280 ;
        RECT 174.530 0.350 176.910 4.280 ;
        RECT 177.750 0.350 180.130 4.280 ;
        RECT 180.970 0.350 183.350 4.280 ;
        RECT 184.190 0.350 186.570 4.280 ;
        RECT 187.410 0.350 189.790 4.280 ;
        RECT 190.630 0.350 193.010 4.280 ;
        RECT 193.850 0.350 196.230 4.280 ;
        RECT 197.070 0.350 199.450 4.280 ;
        RECT 200.290 0.350 202.670 4.280 ;
        RECT 203.510 0.350 205.890 4.280 ;
        RECT 206.730 0.350 209.110 4.280 ;
        RECT 209.950 0.350 212.330 4.280 ;
        RECT 213.170 0.350 215.550 4.280 ;
        RECT 216.390 0.350 218.770 4.280 ;
        RECT 219.610 0.350 221.990 4.280 ;
        RECT 222.830 0.350 225.210 4.280 ;
        RECT 226.050 0.350 228.430 4.280 ;
        RECT 229.270 0.350 231.650 4.280 ;
        RECT 232.490 0.350 234.870 4.280 ;
        RECT 235.710 0.350 238.090 4.280 ;
        RECT 238.930 0.350 241.310 4.280 ;
        RECT 242.150 0.350 244.530 4.280 ;
        RECT 245.370 0.350 247.750 4.280 ;
        RECT 248.590 0.350 250.970 4.280 ;
        RECT 251.810 0.350 254.190 4.280 ;
        RECT 255.030 0.350 257.410 4.280 ;
        RECT 258.250 0.350 260.630 4.280 ;
        RECT 261.470 0.350 263.850 4.280 ;
        RECT 264.690 0.350 267.070 4.280 ;
        RECT 267.910 0.350 270.290 4.280 ;
        RECT 271.130 0.350 273.510 4.280 ;
        RECT 274.350 0.350 276.730 4.280 ;
        RECT 277.570 0.350 279.950 4.280 ;
        RECT 280.790 0.350 283.170 4.280 ;
        RECT 284.010 0.350 286.390 4.280 ;
        RECT 287.230 0.350 289.610 4.280 ;
        RECT 290.450 0.350 292.830 4.280 ;
        RECT 293.670 0.350 296.050 4.280 ;
        RECT 296.890 0.350 299.270 4.280 ;
        RECT 300.110 0.350 302.490 4.280 ;
        RECT 303.330 0.350 305.710 4.280 ;
        RECT 306.550 0.350 308.930 4.280 ;
        RECT 309.770 0.350 312.150 4.280 ;
        RECT 312.990 0.350 315.370 4.280 ;
        RECT 316.210 0.350 318.590 4.280 ;
        RECT 319.430 0.350 321.810 4.280 ;
        RECT 322.650 0.350 325.030 4.280 ;
        RECT 325.870 0.350 328.250 4.280 ;
        RECT 329.090 0.350 331.470 4.280 ;
        RECT 332.310 0.350 334.690 4.280 ;
        RECT 335.530 0.350 337.910 4.280 ;
        RECT 338.750 0.350 341.130 4.280 ;
        RECT 341.970 0.350 344.350 4.280 ;
        RECT 345.190 0.350 347.570 4.280 ;
        RECT 348.410 0.350 350.790 4.280 ;
        RECT 351.630 0.350 354.010 4.280 ;
        RECT 354.850 0.350 357.230 4.280 ;
        RECT 358.070 0.350 360.450 4.280 ;
        RECT 361.290 0.350 363.670 4.280 ;
        RECT 364.510 0.350 366.890 4.280 ;
        RECT 367.730 0.350 370.110 4.280 ;
        RECT 370.950 0.350 373.330 4.280 ;
        RECT 374.170 0.350 376.550 4.280 ;
        RECT 377.390 0.350 379.770 4.280 ;
        RECT 380.610 0.350 382.990 4.280 ;
        RECT 383.830 0.350 386.210 4.280 ;
        RECT 387.050 0.350 388.140 4.280 ;
      LAYER met3 ;
        RECT 17.545 4.935 370.920 187.845 ;
      LAYER met4 ;
        RECT 23.790 10.240 25.240 182.745 ;
        RECT 27.640 10.240 28.540 182.745 ;
        RECT 30.940 10.240 178.840 182.745 ;
        RECT 181.240 10.240 182.140 182.745 ;
        RECT 184.540 10.240 332.440 182.745 ;
        RECT 334.840 10.240 335.740 182.745 ;
        RECT 338.140 10.240 370.890 182.745 ;
        RECT 23.790 4.935 370.890 10.240 ;
      LAYER met5 ;
        RECT 23.580 11.100 371.100 53.500 ;
  END
END ahb_counter
END LIBRARY

