magic
tech sky130A
magscale 1 2
timestamp 1740783807
<< metal1 >>
rect 104618 3816 104624 3868
rect 104676 3856 104682 3868
rect 104802 3856 104808 3868
rect 104676 3828 104808 3856
rect 104676 3816 104682 3828
rect 104802 3816 104808 3828
rect 104860 3816 104866 3868
rect 147122 484 147128 536
rect 147180 524 147186 536
rect 163406 524 163412 536
rect 147180 496 163412 524
rect 147180 484 147186 496
rect 163406 484 163412 496
rect 163464 484 163470 536
rect 137554 416 137560 468
rect 137612 456 137618 468
rect 156322 456 156328 468
rect 137612 428 156328 456
rect 137612 416 137618 428
rect 156322 416 156328 428
rect 156380 416 156386 468
rect 121454 348 121460 400
rect 121512 388 121518 400
rect 154758 388 154764 400
rect 121512 360 154764 388
rect 121512 348 121518 360
rect 154758 348 154764 360
rect 154816 348 154822 400
rect 127342 280 127348 332
rect 127400 320 127406 332
rect 161014 320 161020 332
rect 127400 292 161020 320
rect 127400 280 127406 292
rect 161014 280 161020 292
rect 161072 280 161078 332
rect 111794 212 111800 264
rect 111852 252 111858 264
rect 153194 252 153200 264
rect 111852 224 153200 252
rect 111852 212 111858 224
rect 153194 212 153200 224
rect 153252 212 153258 264
rect 109034 144 109040 196
rect 109092 184 109098 196
rect 157886 184 157892 196
rect 109092 156 157892 184
rect 109092 144 109098 156
rect 157886 144 157892 156
rect 157944 144 157950 196
rect 108298 76 108304 128
rect 108356 116 108362 128
rect 212626 116 212632 128
rect 108356 88 212632 116
rect 108356 76 108362 88
rect 212626 76 212632 88
rect 212684 76 212690 128
rect 110414 8 110420 60
rect 110472 48 110478 60
rect 159450 48 159456 60
rect 110472 20 159456 48
rect 110472 8 110478 20
rect 159450 8 159456 20
rect 159508 8 159514 60
<< via1 >>
rect 104624 3816 104676 3868
rect 104808 3816 104860 3868
rect 147128 484 147180 536
rect 163412 484 163464 536
rect 137560 416 137612 468
rect 156328 416 156380 468
rect 121460 348 121512 400
rect 154764 348 154816 400
rect 127348 280 127400 332
rect 161020 280 161072 332
rect 111800 212 111852 264
rect 153200 212 153252 264
rect 109040 144 109092 196
rect 157892 144 157944 196
rect 108304 76 108356 128
rect 212632 76 212684 128
rect 110420 8 110472 60
rect 159456 8 159508 60
<< metal2 >>
rect 12530 459200 12586 460400
rect 14370 459200 14426 460400
rect 16210 459200 16266 460400
rect 18050 459200 18106 460400
rect 19890 459200 19946 460400
rect 21730 459200 21786 460400
rect 23570 459200 23626 460400
rect 25410 459200 25466 460400
rect 27250 459200 27306 460400
rect 29090 459200 29146 460400
rect 30930 459200 30986 460400
rect 32770 459200 32826 460400
rect 34610 459200 34666 460400
rect 36450 459200 36506 460400
rect 38290 459200 38346 460400
rect 40130 459200 40186 460400
rect 41970 459200 42026 460400
rect 43810 459200 43866 460400
rect 45650 459200 45706 460400
rect 47490 459200 47546 460400
rect 49330 459200 49386 460400
rect 51170 459200 51226 460400
rect 53010 459200 53066 460400
rect 54850 459200 54906 460400
rect 489090 459200 489146 460400
rect 490930 459200 490986 460400
rect 492770 459200 492826 460400
rect 494610 459200 494666 460400
rect 496450 459200 496506 460400
rect 498290 459200 498346 460400
rect 500130 459200 500186 460400
rect 501970 459200 502026 460400
rect 503810 459200 503866 460400
rect 505650 459200 505706 460400
rect 507490 459200 507546 460400
rect 509330 459200 509386 460400
rect 511170 459200 511226 460400
rect 513010 459200 513066 460400
rect 514850 459200 514906 460400
rect 516690 459200 516746 460400
rect 518530 459200 518586 460400
rect 520370 459200 520426 460400
rect 522210 459200 522266 460400
rect 524050 459200 524106 460400
rect 525890 459200 525946 460400
rect 527730 459200 527786 460400
rect 529570 459200 529626 460400
rect 531410 459200 531466 460400
rect 123482 285424 123538 285433
rect 123482 285359 123538 285368
rect 121642 280800 121698 280809
rect 121642 280735 121698 280744
rect 93122 276176 93178 276185
rect 93122 276111 93178 276120
rect 110 266656 166 266665
rect 110 266591 166 266600
rect 124 59401 152 266591
rect 294 252784 350 252793
rect 294 252719 350 252728
rect 308 59537 336 252719
rect 3422 248432 3478 248441
rect 3422 248367 3478 248376
rect 478 235512 534 235521
rect 478 235447 534 235456
rect 492 59673 520 235447
rect 846 225176 902 225185
rect 846 225111 902 225120
rect 860 219434 888 225111
rect 676 219406 888 219434
rect 676 59809 704 219406
rect 846 211304 902 211313
rect 846 211239 902 211248
rect 860 59945 888 211239
rect 1030 197568 1086 197577
rect 1030 197503 1086 197512
rect 1044 60081 1072 197503
rect 1214 179072 1270 179081
rect 1214 179007 1270 179016
rect 1228 60217 1256 179007
rect 3436 62801 3464 248367
rect 14462 234560 14518 234569
rect 14462 234495 14518 234504
rect 14476 162081 14504 234495
rect 92202 183696 92258 183705
rect 92202 183631 92258 183640
rect 14462 162072 14518 162081
rect 14462 162007 14518 162016
rect 3422 62792 3478 62801
rect 3422 62727 3478 62736
rect 1214 60208 1270 60217
rect 1214 60143 1270 60152
rect 1030 60072 1086 60081
rect 1030 60007 1086 60016
rect 846 59936 902 59945
rect 92216 59908 92244 183631
rect 93136 61441 93164 276111
rect 115202 262304 115258 262313
rect 115202 262239 115258 262248
rect 104162 220688 104218 220697
rect 104162 220623 104218 220632
rect 101402 206816 101458 206825
rect 101402 206751 101458 206760
rect 97722 192944 97778 192953
rect 97722 192879 97778 192888
rect 93122 61432 93178 61441
rect 93122 61367 93178 61376
rect 94042 60208 94098 60217
rect 94042 60143 94098 60152
rect 94056 59908 94084 60143
rect 95514 60072 95570 60081
rect 95514 60007 95570 60016
rect 95528 59922 95556 60007
rect 95528 59894 95910 59922
rect 97736 59908 97764 192879
rect 99562 59936 99618 59945
rect 846 59871 902 59880
rect 101416 59908 101444 206751
rect 104176 62121 104204 220623
rect 108762 162072 108818 162081
rect 108762 162007 108818 162016
rect 104162 62112 104218 62121
rect 104162 62047 104218 62056
rect 105082 62112 105138 62121
rect 105082 62047 105138 62056
rect 105096 59908 105124 62047
rect 108776 59908 108804 162007
rect 112442 62792 112498 62801
rect 112442 62727 112498 62736
rect 112456 59908 112484 62727
rect 115216 59945 115244 262239
rect 119802 61432 119858 61441
rect 119802 61367 119858 61376
rect 117962 60208 118018 60217
rect 117962 60143 118018 60152
rect 115202 59936 115258 59945
rect 99562 59871 99618 59880
rect 115202 59871 115258 59880
rect 116122 59936 116178 59945
rect 117976 59908 118004 60143
rect 119816 59908 119844 61367
rect 121656 59908 121684 280735
rect 123496 59908 123524 285359
rect 127162 271552 127218 271561
rect 127162 271487 127218 271496
rect 125322 266928 125378 266937
rect 125322 266863 125378 266872
rect 125336 59908 125364 266863
rect 127176 59908 127204 271487
rect 130842 257680 130898 257689
rect 130842 257615 130898 257624
rect 129002 253056 129058 253065
rect 129002 252991 129058 253000
rect 129016 59908 129044 252991
rect 130856 59908 130884 257615
rect 543278 243536 543334 243545
rect 543278 243471 543334 243480
rect 132682 239184 132738 239193
rect 132682 239119 132738 239128
rect 132696 59908 132724 239119
rect 543094 229800 543150 229809
rect 543094 229735 543150 229744
rect 136362 225312 136418 225321
rect 136362 225247 136418 225256
rect 136376 59908 136404 225247
rect 141882 216064 141938 216073
rect 141882 215999 141938 216008
rect 140042 211440 140098 211449
rect 140042 211375 140098 211384
rect 140056 59908 140084 211375
rect 141896 59908 141924 215999
rect 145562 202192 145618 202201
rect 145562 202127 145618 202136
rect 143722 197568 143778 197577
rect 143722 197503 143778 197512
rect 143736 59908 143764 197503
rect 145576 59908 145604 202127
rect 149242 188320 149298 188329
rect 149242 188255 149298 188264
rect 147402 183696 147458 183705
rect 147402 183631 147458 183640
rect 147416 59908 147444 183631
rect 149256 59908 149284 188255
rect 116122 59871 116178 59880
rect 662 59800 718 59809
rect 662 59735 718 59744
rect 103242 59800 103298 59809
rect 103242 59735 103298 59744
rect 478 59664 534 59673
rect 478 59599 534 59608
rect 106922 59664 106978 59673
rect 106922 59599 106978 59608
rect 543108 59537 543136 229735
rect 294 59528 350 59537
rect 294 59463 350 59472
rect 110602 59528 110658 59537
rect 110602 59463 110658 59472
rect 138202 59528 138258 59537
rect 138202 59463 138258 59472
rect 543094 59528 543150 59537
rect 543094 59463 543150 59472
rect 543292 59401 543320 243471
rect 110 59392 166 59401
rect 110 59327 166 59336
rect 114282 59392 114338 59401
rect 114282 59327 114338 59336
rect 134522 59392 134578 59401
rect 134522 59327 134578 59336
rect 543278 59392 543334 59401
rect 543278 59327 543334 59336
rect 99070 19802 99098 20060
rect 99070 19774 99144 19802
rect 53102 18864 53158 18873
rect 53102 18799 53158 18808
rect 53116 1329 53144 18799
rect 64142 18728 64198 18737
rect 64142 18663 64198 18672
rect 59450 10568 59506 10577
rect 59450 10503 59506 10512
rect 57886 9208 57942 9217
rect 57886 9143 57942 9152
rect 56322 7848 56378 7857
rect 56322 7783 56378 7792
rect 53194 6488 53250 6497
rect 53194 6423 53250 6432
rect 51630 1320 51686 1329
rect 51630 1255 51686 1264
rect 53102 1320 53158 1329
rect 53102 1255 53158 1264
rect 46952 870 47072 898
rect 46952 800 46980 870
rect 46930 -400 46986 800
rect 47044 105 47072 870
rect 48516 870 48636 898
rect 48516 800 48544 870
rect 47030 96 47086 105
rect 47030 31 47086 40
rect 48494 -400 48550 800
rect 48608 241 48636 870
rect 50080 870 50200 898
rect 50080 800 50108 870
rect 48594 232 48650 241
rect 48594 167 48650 176
rect 50058 -400 50114 800
rect 50172 377 50200 870
rect 51644 800 51672 1255
rect 53208 800 53236 6423
rect 54758 2272 54814 2281
rect 54758 2207 54814 2216
rect 54772 800 54800 2207
rect 56336 800 56364 7783
rect 57900 800 57928 9143
rect 59464 800 59492 10503
rect 61014 5128 61070 5137
rect 61014 5063 61070 5072
rect 61028 800 61056 5063
rect 62578 2136 62634 2145
rect 62578 2071 62634 2080
rect 62592 800 62620 2071
rect 64156 800 64184 18663
rect 82910 18592 82966 18601
rect 82910 18527 82966 18536
rect 67270 17368 67326 17377
rect 67270 17303 67326 17312
rect 65706 11928 65762 11937
rect 65706 11863 65762 11872
rect 65720 800 65748 11863
rect 67284 800 67312 17303
rect 68834 16008 68890 16017
rect 68834 15943 68890 15952
rect 68848 800 68876 15943
rect 71962 14648 72018 14657
rect 71962 14583 72018 14592
rect 70398 3496 70454 3505
rect 70398 3431 70454 3440
rect 70412 800 70440 3431
rect 71976 800 72004 14583
rect 73526 13152 73582 13161
rect 73526 13087 73582 13096
rect 73540 800 73568 13087
rect 75090 11792 75146 11801
rect 75090 11727 75146 11736
rect 75104 800 75132 11727
rect 78218 10432 78274 10441
rect 78218 10367 78274 10376
rect 76654 4992 76710 5001
rect 76654 4927 76710 4936
rect 76668 800 76696 4927
rect 78232 800 78260 10367
rect 79782 9072 79838 9081
rect 79782 9007 79838 9016
rect 79796 800 79824 9007
rect 81346 7576 81402 7585
rect 81346 7511 81402 7520
rect 81360 800 81388 7511
rect 82924 800 82952 18527
rect 86038 17232 86094 17241
rect 86038 17167 86094 17176
rect 84474 6216 84530 6225
rect 84474 6151 84530 6160
rect 84488 800 84516 6151
rect 86052 800 86080 17167
rect 89166 15872 89222 15881
rect 89166 15807 89222 15816
rect 87602 3360 87658 3369
rect 87602 3295 87658 3304
rect 87616 800 87644 3295
rect 89180 800 89208 15807
rect 90730 14512 90786 14521
rect 90730 14447 90786 14456
rect 90744 800 90772 14447
rect 92294 13016 92350 13025
rect 92294 12951 92350 12960
rect 92308 800 92336 12951
rect 95422 11656 95478 11665
rect 95422 11591 95478 11600
rect 93858 2000 93914 2009
rect 93858 1935 93914 1944
rect 93872 800 93900 1935
rect 95436 800 95464 11591
rect 96986 10296 97042 10305
rect 96986 10231 97042 10240
rect 97000 800 97028 10231
rect 98550 4856 98606 4865
rect 98550 4791 98606 4800
rect 98564 800 98592 4791
rect 50158 368 50214 377
rect 50158 303 50214 312
rect 51622 -400 51678 800
rect 53186 -400 53242 800
rect 54750 -400 54806 800
rect 56314 -400 56370 800
rect 57878 -400 57934 800
rect 59442 -400 59498 800
rect 61006 -400 61062 800
rect 62570 -400 62626 800
rect 64134 -400 64190 800
rect 65698 -400 65754 800
rect 67262 -400 67318 800
rect 68826 -400 68882 800
rect 70390 -400 70446 800
rect 71954 -400 72010 800
rect 73518 -400 73574 800
rect 75082 -400 75138 800
rect 76646 -400 76702 800
rect 78210 -400 78266 800
rect 79774 -400 79830 800
rect 81338 -400 81394 800
rect 82902 -400 82958 800
rect 84466 -400 84522 800
rect 86030 -400 86086 800
rect 87594 -400 87650 800
rect 89158 -400 89214 800
rect 90722 -400 90778 800
rect 92286 -400 92342 800
rect 93850 -400 93906 800
rect 95414 -400 95470 800
rect 96978 -400 97034 800
rect 98542 -400 98598 800
rect 99116 105 99144 19774
rect 99668 6633 99696 20060
rect 100312 19417 100340 20060
rect 100298 19408 100354 19417
rect 100298 19343 100354 19352
rect 100114 8936 100170 8945
rect 100114 8871 100170 8880
rect 99654 6624 99710 6633
rect 99654 6559 99710 6568
rect 100128 800 100156 8871
rect 99102 96 99158 105
rect 99102 31 99158 40
rect 100106 -400 100162 800
rect 100956 241 100984 20060
rect 101600 6914 101628 20060
rect 101770 19680 101826 19689
rect 101770 19615 101826 19624
rect 101784 6914 101812 19615
rect 101416 6886 101628 6914
rect 101692 6886 101812 6914
rect 101416 377 101444 6886
rect 101692 800 101720 6886
rect 102244 1193 102272 20060
rect 102888 18873 102916 20060
rect 102874 18864 102930 18873
rect 102874 18799 102930 18808
rect 103242 16144 103298 16153
rect 103242 16079 103298 16088
rect 102230 1184 102286 1193
rect 102230 1119 102286 1128
rect 103256 800 103284 16079
rect 103532 6361 103560 20060
rect 103518 6352 103574 6361
rect 103518 6287 103574 6296
rect 104176 1329 104204 20060
rect 104714 18320 104770 18329
rect 104714 18255 104770 18264
rect 104624 3868 104676 3874
rect 104624 3810 104676 3816
rect 104162 1320 104218 1329
rect 104162 1255 104218 1264
rect 104636 921 104664 3810
rect 104728 3482 104756 18255
rect 104820 3874 104848 20060
rect 105464 19689 105492 20060
rect 105450 19680 105506 19689
rect 105450 19615 105506 19624
rect 106108 6497 106136 20060
rect 106370 19544 106426 19553
rect 106370 19479 106426 19488
rect 106094 6488 106150 6497
rect 106094 6423 106150 6432
rect 104808 3868 104860 3874
rect 104808 3810 104860 3816
rect 104728 3454 104848 3482
rect 104622 912 104678 921
rect 104622 847 104678 856
rect 104820 800 104848 3454
rect 106384 800 106412 19479
rect 106752 7721 106780 20060
rect 106738 7712 106794 7721
rect 106738 7647 106794 7656
rect 107396 921 107424 20060
rect 108040 19417 108068 20060
rect 108210 19816 108266 19825
rect 108210 19751 108266 19760
rect 108026 19408 108082 19417
rect 108026 19343 108082 19352
rect 107382 912 107438 921
rect 107382 847 107438 856
rect 107948 870 108068 898
rect 107948 800 107976 870
rect 101402 368 101458 377
rect 101402 303 101458 312
rect 100942 232 100998 241
rect 100942 167 100998 176
rect 101670 -400 101726 800
rect 103234 -400 103290 800
rect 104798 -400 104854 800
rect 106362 -400 106418 800
rect 107926 -400 107982 800
rect 108040 762 108068 870
rect 108224 762 108252 19751
rect 108684 16153 108712 20060
rect 108670 16144 108726 16153
rect 108670 16079 108726 16088
rect 109328 2281 109356 20060
rect 109498 17504 109554 17513
rect 109498 17439 109554 17448
rect 109314 2272 109370 2281
rect 109314 2207 109370 2216
rect 109038 1320 109094 1329
rect 109038 1255 109094 1264
rect 108302 1048 108358 1057
rect 108302 983 108358 992
rect 108040 734 108252 762
rect 108316 134 108344 983
rect 109052 202 109080 1255
rect 109512 800 109540 17439
rect 109972 3641 110000 20060
rect 109958 3632 110014 3641
rect 109958 3567 110014 3576
rect 110616 1329 110644 20060
rect 111260 18329 111288 20060
rect 111246 18320 111302 18329
rect 111246 18255 111302 18264
rect 111904 7857 111932 20060
rect 112548 14793 112576 20060
rect 113192 19553 113220 20060
rect 113178 19544 113234 19553
rect 113178 19479 113234 19488
rect 112534 14784 112590 14793
rect 112534 14719 112590 14728
rect 113836 9217 113864 20060
rect 114480 13297 114508 20060
rect 115124 19825 115152 20060
rect 115110 19816 115166 19825
rect 115110 19751 115166 19760
rect 114466 13288 114522 13297
rect 114466 13223 114522 13232
rect 115768 10577 115796 20060
rect 116412 18873 116440 20060
rect 116398 18864 116454 18873
rect 116398 18799 116454 18808
rect 117056 17513 117084 20060
rect 117042 17504 117098 17513
rect 117042 17439 117098 17448
rect 115754 10568 115810 10577
rect 115754 10503 115810 10512
rect 113822 9208 113878 9217
rect 113822 9143 113878 9152
rect 111890 7848 111946 7857
rect 111890 7783 111946 7792
rect 117700 5137 117728 20060
rect 118344 10577 118372 20060
rect 118988 16574 119016 20060
rect 118988 16546 119200 16574
rect 118330 10568 118386 10577
rect 118330 10503 118386 10512
rect 117686 5128 117742 5137
rect 117686 5063 117742 5072
rect 110602 1320 110658 1329
rect 110602 1255 110658 1264
rect 111798 1184 111854 1193
rect 111798 1119 111854 1128
rect 110418 912 110474 921
rect 110418 847 110474 856
rect 111076 870 111196 898
rect 109040 196 109092 202
rect 109040 138 109092 144
rect 108304 128 108356 134
rect 108304 70 108356 76
rect 109490 -400 109546 800
rect 110432 66 110460 847
rect 111076 800 111104 870
rect 110420 60 110472 66
rect 110420 2 110472 8
rect 111054 -400 111110 800
rect 111168 513 111196 870
rect 111154 504 111210 513
rect 111154 439 111210 448
rect 111812 270 111840 1119
rect 115754 1048 115810 1057
rect 115754 983 115810 992
rect 112640 870 112760 898
rect 112640 800 112668 870
rect 111800 264 111852 270
rect 111800 206 111852 212
rect 112618 -400 112674 800
rect 112732 105 112760 870
rect 114204 870 114324 898
rect 114204 800 114232 870
rect 112718 96 112774 105
rect 112718 31 112774 40
rect 114182 -400 114238 800
rect 114296 377 114324 870
rect 115768 800 115796 983
rect 118882 912 118938 921
rect 117332 870 117452 898
rect 117332 800 117360 870
rect 114282 368 114338 377
rect 114282 303 114338 312
rect 115746 -400 115802 800
rect 117310 -400 117366 800
rect 117424 241 117452 870
rect 118882 847 118938 856
rect 118896 800 118924 847
rect 117410 232 117466 241
rect 117410 167 117466 176
rect 118874 -400 118930 800
rect 119172 513 119200 16546
rect 119632 2145 119660 20060
rect 120276 16153 120304 20060
rect 120262 16144 120318 16153
rect 120262 16079 120318 16088
rect 119618 2136 119674 2145
rect 119618 2071 119674 2080
rect 120460 870 120580 898
rect 120460 800 120488 870
rect 119158 504 119214 513
rect 119158 439 119214 448
rect 120438 -400 120494 800
rect 120552 649 120580 870
rect 120538 640 120594 649
rect 120538 575 120594 584
rect 120920 105 120948 20060
rect 121564 18737 121592 20060
rect 121550 18728 121606 18737
rect 121550 18663 121606 18672
rect 122208 12073 122236 20060
rect 122194 12064 122250 12073
rect 122194 11999 122250 12008
rect 122010 1320 122066 1329
rect 122010 1255 122066 1264
rect 122024 800 122052 1255
rect 121458 776 121514 785
rect 121458 711 121514 720
rect 121472 406 121500 711
rect 121460 400 121512 406
rect 121460 342 121512 348
rect 120906 96 120962 105
rect 120906 31 120962 40
rect 122002 -400 122058 800
rect 122852 377 122880 20060
rect 123496 11937 123524 20060
rect 124140 17513 124168 20060
rect 124126 17504 124182 17513
rect 124126 17439 124182 17448
rect 123482 11928 123538 11937
rect 123482 11863 123538 11872
rect 124784 1057 124812 20060
rect 125428 17377 125456 20060
rect 125414 17368 125470 17377
rect 125414 17303 125470 17312
rect 126072 2145 126100 20060
rect 126716 6914 126744 20060
rect 127360 16017 127388 20060
rect 127346 16008 127402 16017
rect 127346 15943 127402 15952
rect 126440 6886 126744 6914
rect 126058 2136 126114 2145
rect 126058 2071 126114 2080
rect 124770 1048 124826 1057
rect 124770 983 124826 992
rect 123588 870 123708 898
rect 123588 800 123616 870
rect 122838 368 122894 377
rect 122838 303 122894 312
rect 123566 -400 123622 800
rect 123680 785 123708 870
rect 125152 870 125272 898
rect 125152 800 125180 870
rect 123666 776 123722 785
rect 123666 711 123722 720
rect 125130 -400 125186 800
rect 125244 649 125272 870
rect 125230 640 125286 649
rect 125230 575 125286 584
rect 126440 241 126468 6886
rect 128004 2281 128032 20060
rect 127990 2272 128046 2281
rect 127990 2207 128046 2216
rect 127346 1184 127402 1193
rect 127346 1119 127402 1128
rect 126716 870 126836 898
rect 126716 800 126744 870
rect 126426 232 126482 241
rect 126426 167 126482 176
rect 126694 -400 126750 800
rect 126808 105 126836 870
rect 127360 338 127388 1119
rect 128648 921 128676 20060
rect 129292 3505 129320 20060
rect 129936 18737 129964 20060
rect 129922 18728 129978 18737
rect 129922 18663 129978 18672
rect 129278 3496 129334 3505
rect 129278 3431 129334 3440
rect 128634 912 128690 921
rect 128188 870 128308 898
rect 128188 377 128216 870
rect 128280 800 128308 870
rect 128634 847 128690 856
rect 129844 870 129964 898
rect 129844 800 129872 870
rect 128174 368 128230 377
rect 127348 332 127400 338
rect 128174 303 128230 312
rect 127348 274 127400 280
rect 126794 96 126850 105
rect 126794 31 126850 40
rect 128258 -400 128314 800
rect 129822 -400 129878 800
rect 129936 241 129964 870
rect 130580 513 130608 20060
rect 131224 14657 131252 20060
rect 131868 17377 131896 20060
rect 131854 17368 131910 17377
rect 131854 17303 131910 17312
rect 131210 14648 131266 14657
rect 131210 14583 131266 14592
rect 132512 1329 132540 20060
rect 133156 13161 133184 20060
rect 133142 13152 133198 13161
rect 133142 13087 133198 13096
rect 133800 7857 133828 20060
rect 133786 7848 133842 7857
rect 133786 7783 133842 7792
rect 134444 6914 134472 20060
rect 135088 11801 135116 20060
rect 135074 11792 135130 11801
rect 135074 11727 135130 11736
rect 134168 6886 134472 6914
rect 132498 1320 132554 1329
rect 132498 1255 132554 1264
rect 131394 1048 131450 1057
rect 131394 983 131450 992
rect 131408 800 131436 983
rect 132972 870 133092 898
rect 132972 800 133000 870
rect 130566 504 130622 513
rect 130566 439 130622 448
rect 129922 232 129978 241
rect 129922 167 129978 176
rect 131386 -400 131442 800
rect 132950 -400 133006 800
rect 133064 513 133092 870
rect 134168 785 134196 6886
rect 135732 3505 135760 20060
rect 135718 3496 135774 3505
rect 135718 3431 135774 3440
rect 136376 921 136404 20060
rect 137020 5001 137048 20060
rect 137664 5001 137692 20060
rect 137006 4992 137062 5001
rect 137006 4927 137062 4936
rect 137650 4992 137706 5001
rect 137650 4927 137706 4936
rect 137558 1048 137614 1057
rect 137558 983 137614 992
rect 136362 912 136418 921
rect 134536 870 134656 898
rect 134536 800 134564 870
rect 134154 776 134210 785
rect 134154 711 134210 720
rect 133050 504 133106 513
rect 133050 439 133106 448
rect 134514 -400 134570 800
rect 134628 649 134656 870
rect 136100 870 136220 898
rect 136100 800 136128 870
rect 134614 640 134670 649
rect 134614 575 134670 584
rect 136078 -400 136134 800
rect 136192 785 136220 870
rect 136362 847 136418 856
rect 136178 776 136234 785
rect 136178 711 136234 720
rect 137572 474 137600 983
rect 137650 912 137706 921
rect 137650 847 137706 856
rect 137664 800 137692 847
rect 137560 468 137612 474
rect 137560 410 137612 416
rect 137642 -400 137698 800
rect 138308 105 138336 20060
rect 138952 10441 138980 20060
rect 139596 16017 139624 20060
rect 139582 16008 139638 16017
rect 139582 15943 139638 15952
rect 138938 10432 138994 10441
rect 138938 10367 138994 10376
rect 139582 912 139638 921
rect 139228 870 139348 898
rect 139228 800 139256 870
rect 138294 96 138350 105
rect 138294 31 138350 40
rect 139206 -400 139262 800
rect 139320 785 139348 870
rect 139582 847 139638 856
rect 139306 776 139362 785
rect 139306 711 139362 720
rect 139596 513 139624 847
rect 139582 504 139638 513
rect 139582 439 139638 448
rect 140240 377 140268 20060
rect 140884 9081 140912 20060
rect 141528 14657 141556 20060
rect 141514 14648 141570 14657
rect 141514 14583 141570 14592
rect 140870 9072 140926 9081
rect 140870 9007 140926 9016
rect 140792 870 140912 898
rect 140792 800 140820 870
rect 140226 368 140282 377
rect 140226 303 140282 312
rect 140770 -400 140826 800
rect 140884 513 140912 870
rect 140870 504 140926 513
rect 140870 439 140926 448
rect 142066 232 142122 241
rect 142172 218 142200 20060
rect 142816 7585 142844 20060
rect 143460 13161 143488 20060
rect 143446 13152 143502 13161
rect 143446 13087 143502 13096
rect 142802 7576 142858 7585
rect 142802 7511 142858 7520
rect 144104 1329 144132 20060
rect 144748 18601 144776 20060
rect 144734 18592 144790 18601
rect 144734 18527 144790 18536
rect 145392 11801 145420 20060
rect 145378 11792 145434 11801
rect 145378 11727 145434 11736
rect 144090 1320 144146 1329
rect 144090 1255 144146 1264
rect 146036 921 146064 20060
rect 146680 6225 146708 20060
rect 147324 6225 147352 20060
rect 146666 6216 146722 6225
rect 146666 6151 146722 6160
rect 147310 6216 147366 6225
rect 147310 6151 147366 6160
rect 146022 912 146078 921
rect 142356 870 142476 898
rect 142356 800 142384 870
rect 142122 190 142200 218
rect 142066 167 142122 176
rect 142334 -400 142390 800
rect 142448 105 142476 870
rect 143920 870 144040 898
rect 143920 800 143948 870
rect 142434 96 142490 105
rect 142434 31 142490 40
rect 143898 -400 143954 800
rect 144012 241 144040 870
rect 145484 870 145604 898
rect 145484 800 145512 870
rect 143998 232 144054 241
rect 143998 167 144054 176
rect 145462 -400 145518 800
rect 145576 377 145604 870
rect 146022 847 146078 856
rect 147048 870 147168 898
rect 147048 800 147076 870
rect 145562 368 145618 377
rect 145562 303 145618 312
rect 147026 -400 147082 800
rect 147140 542 147168 870
rect 147968 649 147996 20060
rect 148612 17241 148640 20060
rect 148598 17232 148654 17241
rect 148598 17167 148654 17176
rect 149256 10441 149284 20060
rect 149242 10432 149298 10441
rect 149242 10367 149298 10376
rect 149900 1057 149928 20060
rect 150544 3369 150572 20060
rect 151188 9081 151216 20060
rect 151832 19417 151860 20060
rect 151818 19408 151874 19417
rect 151818 19343 151874 19352
rect 152476 15881 152504 20060
rect 153120 18601 153148 20060
rect 153106 18592 153162 18601
rect 153106 18527 153162 18536
rect 152462 15872 152518 15881
rect 152462 15807 152518 15816
rect 151174 9072 151230 9081
rect 151174 9007 151230 9016
rect 151726 6624 151782 6633
rect 151726 6559 151782 6568
rect 150530 3360 150586 3369
rect 150530 3295 150586 3304
rect 149886 1048 149942 1057
rect 149886 983 149942 992
rect 150162 912 150218 921
rect 148612 870 148732 898
rect 148612 800 148640 870
rect 147954 640 148010 649
rect 147954 575 148010 584
rect 147128 536 147180 542
rect 147128 478 147180 484
rect 148590 -400 148646 800
rect 148704 649 148732 870
rect 150162 847 150218 856
rect 150176 800 150204 847
rect 151740 800 151768 6559
rect 153212 870 153332 898
rect 148690 640 148746 649
rect 148690 575 148746 584
rect 150154 -400 150210 800
rect 151718 -400 151774 800
rect 153212 270 153240 870
rect 153304 800 153332 870
rect 153200 264 153252 270
rect 153200 206 153252 212
rect 153282 -400 153338 800
rect 153764 785 153792 20060
rect 154408 14521 154436 20060
rect 155052 17241 155080 20060
rect 155038 17232 155094 17241
rect 155038 17167 155094 17176
rect 154394 14512 154450 14521
rect 154394 14447 154450 14456
rect 154776 870 154896 898
rect 153750 776 153806 785
rect 153750 711 153806 720
rect 154776 406 154804 870
rect 154868 800 154896 870
rect 154764 400 154816 406
rect 154764 342 154816 348
rect 154846 -400 154902 800
rect 155696 513 155724 20060
rect 156340 13025 156368 20060
rect 156984 15881 157012 20060
rect 156970 15872 157026 15881
rect 156970 15807 157026 15816
rect 156326 13016 156382 13025
rect 156326 12951 156382 12960
rect 156340 870 156460 898
rect 155682 504 155738 513
rect 156340 474 156368 870
rect 156432 800 156460 870
rect 155682 439 155738 448
rect 156328 468 156380 474
rect 156328 410 156380 416
rect 156410 -400 156466 800
rect 157628 105 157656 20060
rect 158272 2009 158300 20060
rect 158258 2000 158314 2009
rect 158258 1935 158314 1944
rect 157904 870 158024 898
rect 157904 202 157932 870
rect 157996 800 158024 870
rect 157892 196 157944 202
rect 157892 138 157944 144
rect 157614 96 157670 105
rect 157614 31 157670 40
rect 157974 -400 158030 800
rect 158916 105 158944 20060
rect 159560 16574 159588 20060
rect 159560 16546 159864 16574
rect 159468 870 159588 898
rect 158902 96 158958 105
rect 159468 66 159496 870
rect 159560 800 159588 870
rect 158902 31 158958 40
rect 159456 60 159508 66
rect 159456 2 159508 8
rect 159538 -400 159594 800
rect 159836 241 159864 16546
rect 160204 11665 160232 20060
rect 160190 11656 160246 11665
rect 160190 11591 160246 11600
rect 160848 241 160876 20060
rect 161032 870 161152 898
rect 161032 338 161060 870
rect 161124 800 161152 870
rect 161020 332 161072 338
rect 161020 274 161072 280
rect 159822 232 159878 241
rect 159822 167 159878 176
rect 160834 232 160890 241
rect 160834 167 160890 176
rect 161102 -400 161158 800
rect 161492 377 161520 20060
rect 162136 10305 162164 20060
rect 162122 10296 162178 10305
rect 162122 10231 162178 10240
rect 162674 6352 162730 6361
rect 162674 6287 162730 6296
rect 162688 800 162716 6287
rect 161478 368 161534 377
rect 161478 303 161534 312
rect 162666 -400 162722 800
rect 162780 354 162808 20060
rect 163424 542 163452 20060
rect 164068 4865 164096 20060
rect 164238 7712 164294 7721
rect 164238 7647 164294 7656
rect 164054 4856 164110 4865
rect 164054 4791 164110 4800
rect 164252 800 164280 7647
rect 163412 536 163464 542
rect 163412 478 163464 484
rect 162950 368 163006 377
rect 162780 326 162950 354
rect 162950 303 163006 312
rect 164230 -400 164286 800
rect 164712 513 164740 20060
rect 165356 649 165384 20060
rect 166000 8945 166028 20060
rect 165986 8936 166042 8945
rect 165986 8871 166042 8880
rect 165802 3632 165858 3641
rect 165802 3567 165858 3576
rect 165816 800 165844 3567
rect 165342 640 165398 649
rect 165342 575 165398 584
rect 164698 504 164754 513
rect 164698 439 164754 448
rect 165794 -400 165850 800
rect 166644 649 166672 20060
rect 167288 921 167316 20060
rect 170494 18864 170550 18873
rect 170494 18799 170550 18808
rect 167366 14784 167422 14793
rect 167366 14719 167422 14728
rect 167274 912 167330 921
rect 167274 847 167330 856
rect 167380 800 167408 14719
rect 168930 13288 168986 13297
rect 168930 13223 168986 13232
rect 168944 800 168972 13223
rect 170508 800 170536 18799
rect 181442 18728 181498 18737
rect 181442 18663 181498 18672
rect 176750 17504 176806 17513
rect 176750 17439 176806 17448
rect 173622 16144 173678 16153
rect 173622 16079 173678 16088
rect 172058 10568 172114 10577
rect 172058 10503 172114 10512
rect 172072 800 172100 10503
rect 173636 800 173664 16079
rect 175186 12064 175242 12073
rect 175186 11999 175242 12008
rect 175200 800 175228 11999
rect 176764 800 176792 17439
rect 179878 2272 179934 2281
rect 179878 2207 179934 2216
rect 178314 2136 178370 2145
rect 178314 2071 178370 2080
rect 178328 800 178356 2071
rect 179892 800 179920 2207
rect 181456 800 181484 18663
rect 200210 18592 200266 18601
rect 200210 18527 200266 18536
rect 183006 17368 183062 17377
rect 183006 17303 183062 17312
rect 183020 800 183048 17303
rect 189262 16008 189318 16017
rect 189262 15943 189318 15952
rect 184570 7848 184626 7857
rect 184570 7783 184626 7792
rect 184584 800 184612 7783
rect 187698 4992 187754 5001
rect 187698 4927 187754 4936
rect 186134 3496 186190 3505
rect 186134 3431 186190 3440
rect 186148 800 186176 3431
rect 187712 800 187740 4927
rect 189276 800 189304 15943
rect 190826 14648 190882 14657
rect 190826 14583 190882 14592
rect 190840 800 190868 14583
rect 192390 13152 192446 13161
rect 192390 13087 192446 13096
rect 192404 800 192432 13087
rect 193954 11792 194010 11801
rect 193954 11727 194010 11736
rect 193968 800 193996 11727
rect 197082 10432 197138 10441
rect 197082 10367 197138 10376
rect 195518 6216 195574 6225
rect 195518 6151 195574 6160
rect 195532 800 195560 6151
rect 197096 800 197124 10367
rect 198646 9072 198702 9081
rect 198646 9007 198702 9016
rect 198660 800 198688 9007
rect 200224 800 200252 18527
rect 201774 17232 201830 17241
rect 201774 17167 201830 17176
rect 201788 800 201816 17167
rect 203338 15872 203394 15881
rect 203338 15807 203394 15816
rect 203352 800 203380 15807
rect 204824 870 204944 898
rect 166630 640 166686 649
rect 166630 575 166686 584
rect 167358 -400 167414 800
rect 168922 -400 168978 800
rect 170486 -400 170542 800
rect 172050 -400 172106 800
rect 173614 -400 173670 800
rect 175178 -400 175234 800
rect 176742 -400 176798 800
rect 178306 -400 178362 800
rect 179870 -400 179926 800
rect 181434 -400 181490 800
rect 182998 -400 183054 800
rect 184562 -400 184618 800
rect 186126 -400 186182 800
rect 187690 -400 187746 800
rect 189254 -400 189310 800
rect 190818 -400 190874 800
rect 192382 -400 192438 800
rect 193946 -400 194002 800
rect 195510 -400 195566 800
rect 197074 -400 197130 800
rect 198638 -400 198694 800
rect 200202 -400 200258 800
rect 201766 -400 201822 800
rect 203330 -400 203386 800
rect 204824 105 204852 870
rect 204916 800 204944 870
rect 206388 870 206508 898
rect 204810 96 204866 105
rect 204810 31 204866 40
rect 204894 -400 204950 800
rect 206388 241 206416 870
rect 206480 800 206508 870
rect 207952 870 208072 898
rect 206374 232 206430 241
rect 206374 167 206430 176
rect 206458 -400 206514 800
rect 207952 377 207980 870
rect 208044 800 208072 870
rect 209516 870 209636 898
rect 207938 368 207994 377
rect 207938 303 207994 312
rect 208022 -400 208078 800
rect 209516 513 209544 870
rect 209608 800 209636 870
rect 211172 870 211292 898
rect 211172 800 211200 870
rect 209502 504 209558 513
rect 209502 439 209558 448
rect 209586 -400 209642 800
rect 211150 -400 211206 800
rect 211264 649 211292 870
rect 212644 870 212764 898
rect 211250 640 211306 649
rect 211250 575 211306 584
rect 212644 134 212672 870
rect 212736 800 212764 870
rect 212632 128 212684 134
rect 212632 70 212684 76
rect 212714 -400 212770 800
rect 214278 -400 214334 800
rect 215842 -400 215898 800
rect 217406 -400 217462 800
rect 218970 -400 219026 800
rect 220534 -400 220590 800
rect 222098 -400 222154 800
rect 223662 -400 223718 800
rect 225226 -400 225282 800
rect 226790 -400 226846 800
rect 228354 -400 228410 800
rect 229918 -400 229974 800
rect 231482 -400 231538 800
rect 233046 -400 233102 800
rect 234610 -400 234666 800
rect 236174 -400 236230 800
rect 237738 -400 237794 800
rect 489194 -400 489250 800
rect 490758 -400 490814 800
rect 492322 -400 492378 800
rect 493886 -400 493942 800
rect 495450 -400 495506 800
rect 497014 -400 497070 800
<< via2 >>
rect 123482 285368 123538 285424
rect 121642 280744 121698 280800
rect 93122 276120 93178 276176
rect 110 266600 166 266656
rect 294 252728 350 252784
rect 3422 248376 3478 248432
rect 478 235456 534 235512
rect 846 225120 902 225176
rect 846 211248 902 211304
rect 1030 197512 1086 197568
rect 1214 179016 1270 179072
rect 14462 234504 14518 234560
rect 92202 183640 92258 183696
rect 14462 162016 14518 162072
rect 3422 62736 3478 62792
rect 1214 60152 1270 60208
rect 1030 60016 1086 60072
rect 846 59880 902 59936
rect 115202 262248 115258 262304
rect 104162 220632 104218 220688
rect 101402 206760 101458 206816
rect 97722 192888 97778 192944
rect 93122 61376 93178 61432
rect 94042 60152 94098 60208
rect 95514 60016 95570 60072
rect 99562 59880 99618 59936
rect 108762 162016 108818 162072
rect 104162 62056 104218 62112
rect 105082 62056 105138 62112
rect 112442 62736 112498 62792
rect 119802 61376 119858 61432
rect 117962 60152 118018 60208
rect 115202 59880 115258 59936
rect 116122 59880 116178 59936
rect 127162 271496 127218 271552
rect 125322 266872 125378 266928
rect 130842 257624 130898 257680
rect 129002 253000 129058 253056
rect 543278 243480 543334 243536
rect 132682 239128 132738 239184
rect 543094 229744 543150 229800
rect 136362 225256 136418 225312
rect 141882 216008 141938 216064
rect 140042 211384 140098 211440
rect 145562 202136 145618 202192
rect 143722 197512 143778 197568
rect 149242 188264 149298 188320
rect 147402 183640 147458 183696
rect 662 59744 718 59800
rect 103242 59744 103298 59800
rect 478 59608 534 59664
rect 106922 59608 106978 59664
rect 294 59472 350 59528
rect 110602 59472 110658 59528
rect 138202 59472 138258 59528
rect 543094 59472 543150 59528
rect 110 59336 166 59392
rect 114282 59336 114338 59392
rect 134522 59336 134578 59392
rect 543278 59336 543334 59392
rect 53102 18808 53158 18864
rect 64142 18672 64198 18728
rect 59450 10512 59506 10568
rect 57886 9152 57942 9208
rect 56322 7792 56378 7848
rect 53194 6432 53250 6488
rect 51630 1264 51686 1320
rect 53102 1264 53158 1320
rect 47030 40 47086 96
rect 48594 176 48650 232
rect 54758 2216 54814 2272
rect 61014 5072 61070 5128
rect 62578 2080 62634 2136
rect 82910 18536 82966 18592
rect 67270 17312 67326 17368
rect 65706 11872 65762 11928
rect 68834 15952 68890 16008
rect 71962 14592 72018 14648
rect 70398 3440 70454 3496
rect 73526 13096 73582 13152
rect 75090 11736 75146 11792
rect 78218 10376 78274 10432
rect 76654 4936 76710 4992
rect 79782 9016 79838 9072
rect 81346 7520 81402 7576
rect 86038 17176 86094 17232
rect 84474 6160 84530 6216
rect 89166 15816 89222 15872
rect 87602 3304 87658 3360
rect 90730 14456 90786 14512
rect 92294 12960 92350 13016
rect 95422 11600 95478 11656
rect 93858 1944 93914 2000
rect 96986 10240 97042 10296
rect 98550 4800 98606 4856
rect 50158 312 50214 368
rect 100298 19352 100354 19408
rect 100114 8880 100170 8936
rect 99654 6568 99710 6624
rect 99102 40 99158 96
rect 101770 19624 101826 19680
rect 102874 18808 102930 18864
rect 103242 16088 103298 16144
rect 102230 1128 102286 1184
rect 103518 6296 103574 6352
rect 104714 18264 104770 18320
rect 104162 1264 104218 1320
rect 105450 19624 105506 19680
rect 106370 19488 106426 19544
rect 106094 6432 106150 6488
rect 104622 856 104678 912
rect 106738 7656 106794 7712
rect 108210 19760 108266 19816
rect 108026 19352 108082 19408
rect 107382 856 107438 912
rect 101402 312 101458 368
rect 100942 176 100998 232
rect 108670 16088 108726 16144
rect 109498 17448 109554 17504
rect 109314 2216 109370 2272
rect 109038 1264 109094 1320
rect 108302 992 108358 1048
rect 109958 3576 110014 3632
rect 111246 18264 111302 18320
rect 113178 19488 113234 19544
rect 112534 14728 112590 14784
rect 115110 19760 115166 19816
rect 114466 13232 114522 13288
rect 116398 18808 116454 18864
rect 117042 17448 117098 17504
rect 115754 10512 115810 10568
rect 113822 9152 113878 9208
rect 111890 7792 111946 7848
rect 118330 10512 118386 10568
rect 117686 5072 117742 5128
rect 110602 1264 110658 1320
rect 111798 1128 111854 1184
rect 110418 856 110474 912
rect 111154 448 111210 504
rect 115754 992 115810 1048
rect 112718 40 112774 96
rect 114282 312 114338 368
rect 118882 856 118938 912
rect 117410 176 117466 232
rect 120262 16088 120318 16144
rect 119618 2080 119674 2136
rect 119158 448 119214 504
rect 120538 584 120594 640
rect 121550 18672 121606 18728
rect 122194 12008 122250 12064
rect 122010 1264 122066 1320
rect 121458 720 121514 776
rect 120906 40 120962 96
rect 124126 17448 124182 17504
rect 123482 11872 123538 11928
rect 125414 17312 125470 17368
rect 127346 15952 127402 16008
rect 126058 2080 126114 2136
rect 124770 992 124826 1048
rect 122838 312 122894 368
rect 123666 720 123722 776
rect 125230 584 125286 640
rect 127990 2216 128046 2272
rect 127346 1128 127402 1184
rect 126426 176 126482 232
rect 129922 18672 129978 18728
rect 129278 3440 129334 3496
rect 128634 856 128690 912
rect 128174 312 128230 368
rect 126794 40 126850 96
rect 131854 17312 131910 17368
rect 131210 14592 131266 14648
rect 133142 13096 133198 13152
rect 133786 7792 133842 7848
rect 135074 11736 135130 11792
rect 132498 1264 132554 1320
rect 131394 992 131450 1048
rect 130566 448 130622 504
rect 129922 176 129978 232
rect 135718 3440 135774 3496
rect 137006 4936 137062 4992
rect 137650 4936 137706 4992
rect 137558 992 137614 1048
rect 134154 720 134210 776
rect 133050 448 133106 504
rect 134614 584 134670 640
rect 136362 856 136418 912
rect 136178 720 136234 776
rect 137650 856 137706 912
rect 139582 15952 139638 16008
rect 138938 10376 138994 10432
rect 138294 40 138350 96
rect 139582 856 139638 912
rect 139306 720 139362 776
rect 139582 448 139638 504
rect 141514 14592 141570 14648
rect 140870 9016 140926 9072
rect 140226 312 140282 368
rect 140870 448 140926 504
rect 142066 176 142122 232
rect 143446 13096 143502 13152
rect 142802 7520 142858 7576
rect 144734 18536 144790 18592
rect 145378 11736 145434 11792
rect 144090 1264 144146 1320
rect 146666 6160 146722 6216
rect 147310 6160 147366 6216
rect 142434 40 142490 96
rect 143998 176 144054 232
rect 146022 856 146078 912
rect 145562 312 145618 368
rect 148598 17176 148654 17232
rect 149242 10376 149298 10432
rect 151818 19352 151874 19408
rect 153106 18536 153162 18592
rect 152462 15816 152518 15872
rect 151174 9016 151230 9072
rect 151726 6568 151782 6624
rect 150530 3304 150586 3360
rect 149886 992 149942 1048
rect 147954 584 148010 640
rect 150162 856 150218 912
rect 148690 584 148746 640
rect 155038 17176 155094 17232
rect 154394 14456 154450 14512
rect 153750 720 153806 776
rect 156970 15816 157026 15872
rect 156326 12960 156382 13016
rect 155682 448 155738 504
rect 158258 1944 158314 2000
rect 157614 40 157670 96
rect 158902 40 158958 96
rect 160190 11600 160246 11656
rect 159822 176 159878 232
rect 160834 176 160890 232
rect 162122 10240 162178 10296
rect 162674 6296 162730 6352
rect 161478 312 161534 368
rect 164238 7656 164294 7712
rect 164054 4800 164110 4856
rect 162950 312 163006 368
rect 165986 8880 166042 8936
rect 165802 3576 165858 3632
rect 165342 584 165398 640
rect 164698 448 164754 504
rect 170494 18808 170550 18864
rect 167366 14728 167422 14784
rect 167274 856 167330 912
rect 168930 13232 168986 13288
rect 181442 18672 181498 18728
rect 176750 17448 176806 17504
rect 173622 16088 173678 16144
rect 172058 10512 172114 10568
rect 175186 12008 175242 12064
rect 179878 2216 179934 2272
rect 178314 2080 178370 2136
rect 200210 18536 200266 18592
rect 183006 17312 183062 17368
rect 189262 15952 189318 16008
rect 184570 7792 184626 7848
rect 187698 4936 187754 4992
rect 186134 3440 186190 3496
rect 190826 14592 190882 14648
rect 192390 13096 192446 13152
rect 193954 11736 194010 11792
rect 197082 10376 197138 10432
rect 195518 6160 195574 6216
rect 198646 9016 198702 9072
rect 201774 17176 201830 17232
rect 203338 15816 203394 15872
rect 166630 584 166686 640
rect 204810 40 204866 96
rect 206374 176 206430 232
rect 207938 312 207994 368
rect 209502 448 209558 504
rect 211250 584 211306 640
<< metal3 >>
rect -400 456824 800 456944
rect 543200 456424 544400 456544
rect -400 452200 800 452320
rect 543200 451800 544400 451920
rect -400 447576 800 447696
rect 543200 447176 544400 447296
rect -400 442952 800 443072
rect 543200 442552 544400 442672
rect -400 438328 800 438448
rect 543200 437928 544400 438048
rect -400 433704 800 433824
rect 543200 433304 544400 433424
rect -400 429080 800 429200
rect 543200 428680 544400 428800
rect -400 424456 800 424576
rect 543200 424056 544400 424176
rect -400 419832 800 419952
rect 543200 419432 544400 419552
rect -400 415208 800 415328
rect 543200 414808 544400 414928
rect -400 410584 800 410704
rect 543200 410184 544400 410304
rect -400 405960 800 406080
rect 543200 405560 544400 405680
rect 0 380308 644 385088
rect 543356 378550 544000 383330
rect 0 370329 644 375109
rect 543356 368571 544000 373351
rect 0 357308 644 362088
rect 543356 354551 544000 359331
rect 0 347329 644 352109
rect 543356 344572 544000 349352
rect -400 340824 800 340944
rect 543200 340824 544400 340944
rect -400 336200 800 336320
rect 543200 336200 544400 336320
rect -400 331576 800 331696
rect 543200 331576 544400 331696
rect -400 326952 800 327072
rect 543200 326952 544400 327072
rect -400 322328 800 322448
rect 543200 322328 544400 322448
rect -400 317704 800 317824
rect 543200 317704 544400 317824
rect -400 313080 800 313200
rect 543200 313080 544400 313200
rect -400 308456 800 308576
rect 543200 308456 544400 308576
rect -400 303832 800 303952
rect 543200 303832 544400 303952
rect -400 299208 800 299328
rect 543200 299208 544400 299328
rect -400 294584 800 294704
rect 543200 294584 544400 294704
rect -400 289960 800 290080
rect 543200 289960 544400 290080
rect -400 285336 800 285456
rect 123477 285426 123543 285429
rect 543200 285426 544400 285456
rect 123477 285424 544400 285426
rect 123477 285368 123482 285424
rect 123538 285368 544400 285424
rect 123477 285366 544400 285368
rect 123477 285363 123543 285366
rect 543200 285336 544400 285366
rect -400 280802 800 280832
rect 121637 280802 121703 280805
rect 543200 280802 544400 280832
rect -400 280742 1042 280802
rect -400 280712 800 280742
rect 54 280468 60 280532
rect 124 280530 130 280532
rect 982 280530 1042 280742
rect 121637 280800 544400 280802
rect 121637 280744 121642 280800
rect 121698 280744 544400 280800
rect 121637 280742 544400 280744
rect 121637 280739 121703 280742
rect 543200 280712 544400 280742
rect 124 280470 1042 280530
rect 124 280468 130 280470
rect -400 276178 800 276208
rect 93117 276178 93183 276181
rect -400 276176 93183 276178
rect -400 276120 93122 276176
rect 93178 276120 93183 276176
rect -400 276118 93183 276120
rect -400 276088 800 276118
rect 93117 276115 93183 276118
rect 543200 276088 544400 276208
rect -400 271464 800 271584
rect 127157 271554 127223 271557
rect 543200 271554 544400 271584
rect 127157 271552 544400 271554
rect 127157 271496 127162 271552
rect 127218 271496 544400 271552
rect 127157 271494 544400 271496
rect 127157 271491 127223 271494
rect 543200 271464 544400 271494
rect -400 266930 800 266960
rect 125317 266930 125383 266933
rect 543200 266930 544400 266960
rect -400 266870 1042 266930
rect -400 266840 800 266870
rect 105 266658 171 266661
rect 982 266658 1042 266870
rect 125317 266928 544400 266930
rect 125317 266872 125322 266928
rect 125378 266872 544400 266928
rect 125317 266870 544400 266872
rect 125317 266867 125383 266870
rect 543200 266840 544400 266870
rect 105 266656 1042 266658
rect 105 266600 110 266656
rect 166 266600 1042 266656
rect 105 266598 1042 266600
rect 105 266595 171 266598
rect -400 262306 800 262336
rect 115197 262306 115263 262309
rect -400 262304 115263 262306
rect -400 262248 115202 262304
rect 115258 262248 115263 262304
rect -400 262246 115263 262248
rect -400 262216 800 262246
rect 115197 262243 115263 262246
rect 543200 262216 544400 262336
rect -400 257592 800 257712
rect 130837 257682 130903 257685
rect 543200 257682 544400 257712
rect 130837 257680 544400 257682
rect 130837 257624 130842 257680
rect 130898 257624 544400 257680
rect 130837 257622 544400 257624
rect 130837 257619 130903 257622
rect 543200 257592 544400 257622
rect -400 253058 800 253088
rect 128997 253058 129063 253061
rect 543200 253058 544400 253088
rect -400 252998 1042 253058
rect -400 252968 800 252998
rect 289 252786 355 252789
rect 982 252786 1042 252998
rect 128997 253056 544400 253058
rect 128997 253000 129002 253056
rect 129058 253000 544400 253056
rect 128997 252998 544400 253000
rect 128997 252995 129063 252998
rect 543200 252968 544400 252998
rect 289 252784 1042 252786
rect 289 252728 294 252784
rect 350 252728 1042 252784
rect 289 252726 1042 252728
rect 289 252723 355 252726
rect -400 248434 800 248464
rect 3417 248434 3483 248437
rect -400 248432 3483 248434
rect -400 248376 3422 248432
rect 3478 248376 3483 248432
rect -400 248374 3483 248376
rect -400 248344 800 248374
rect 3417 248371 3483 248374
rect 543200 248344 544400 248464
rect -400 243720 800 243840
rect 543200 243810 544400 243840
rect 543046 243750 544400 243810
rect 543046 243538 543106 243750
rect 543200 243720 544400 243750
rect 543273 243538 543339 243541
rect 543046 243536 543339 243538
rect 543046 243480 543278 243536
rect 543334 243480 543339 243536
rect 543046 243478 543339 243480
rect 543273 243475 543339 243478
rect -400 239188 800 239216
rect -400 239124 796 239188
rect 860 239124 866 239188
rect 132677 239186 132743 239189
rect 543200 239186 544400 239216
rect 132677 239184 544400 239186
rect 132677 239128 132682 239184
rect 132738 239128 544400 239184
rect 132677 239126 544400 239128
rect -400 239096 800 239124
rect 132677 239123 132743 239126
rect 543200 239096 544400 239126
rect 473 235514 539 235517
rect 790 235514 796 235516
rect 473 235512 796 235514
rect 473 235456 478 235512
rect 534 235456 796 235512
rect 473 235454 796 235456
rect 473 235451 539 235454
rect 790 235452 796 235454
rect 860 235452 866 235516
rect -400 234562 800 234592
rect 14457 234562 14523 234565
rect -400 234560 14523 234562
rect -400 234504 14462 234560
rect 14518 234504 14523 234560
rect -400 234502 14523 234504
rect -400 234472 800 234502
rect 14457 234499 14523 234502
rect 543200 234472 544400 234592
rect -400 229848 800 229968
rect 543200 229938 544400 229968
rect 543046 229878 544400 229938
rect 543046 229805 543106 229878
rect 543200 229848 544400 229878
rect 543046 229800 543155 229805
rect 543046 229744 543094 229800
rect 543150 229744 543155 229800
rect 543046 229742 543155 229744
rect 543089 229739 543155 229742
rect -400 225314 800 225344
rect 136357 225314 136423 225317
rect 543200 225314 544400 225344
rect -400 225224 858 225314
rect 136357 225312 544400 225314
rect 136357 225256 136362 225312
rect 136418 225256 544400 225312
rect 136357 225254 544400 225256
rect 136357 225251 136423 225254
rect 543200 225224 544400 225254
rect 798 225181 858 225224
rect 798 225176 907 225181
rect 798 225120 846 225176
rect 902 225120 907 225176
rect 798 225118 907 225120
rect 841 225115 907 225118
rect -400 220690 800 220720
rect 104157 220690 104223 220693
rect -400 220688 104223 220690
rect -400 220632 104162 220688
rect 104218 220632 104223 220688
rect -400 220630 104223 220632
rect -400 220600 800 220630
rect 104157 220627 104223 220630
rect 543200 220600 544400 220720
rect -400 215976 800 216096
rect 141877 216066 141943 216069
rect 543200 216066 544400 216096
rect 141877 216064 544400 216066
rect 141877 216008 141882 216064
rect 141938 216008 544400 216064
rect 141877 216006 544400 216008
rect 141877 216003 141943 216006
rect 543200 215976 544400 216006
rect -400 211442 800 211472
rect 140037 211442 140103 211445
rect 543200 211442 544400 211472
rect -400 211352 858 211442
rect 140037 211440 544400 211442
rect 140037 211384 140042 211440
rect 140098 211384 544400 211440
rect 140037 211382 544400 211384
rect 140037 211379 140103 211382
rect 543200 211352 544400 211382
rect 798 211309 858 211352
rect 798 211304 907 211309
rect 798 211248 846 211304
rect 902 211248 907 211304
rect 798 211246 907 211248
rect 841 211243 907 211246
rect -400 206818 800 206848
rect 101397 206818 101463 206821
rect -400 206816 101463 206818
rect -400 206760 101402 206816
rect 101458 206760 101463 206816
rect -400 206758 101463 206760
rect -400 206728 800 206758
rect 101397 206755 101463 206758
rect 543200 206728 544400 206848
rect -400 202104 800 202224
rect 145557 202194 145623 202197
rect 543200 202194 544400 202224
rect 145557 202192 544400 202194
rect 145557 202136 145562 202192
rect 145618 202136 544400 202192
rect 145557 202134 544400 202136
rect 145557 202131 145623 202134
rect 543200 202104 544400 202134
rect -400 197570 800 197600
rect 1025 197570 1091 197573
rect -400 197568 1091 197570
rect -400 197512 1030 197568
rect 1086 197512 1091 197568
rect -400 197510 1091 197512
rect -400 197480 800 197510
rect 1025 197507 1091 197510
rect 143717 197570 143783 197573
rect 543200 197570 544400 197600
rect 143717 197568 544400 197570
rect 143717 197512 143722 197568
rect 143778 197512 544400 197568
rect 143717 197510 544400 197512
rect 143717 197507 143783 197510
rect 543200 197480 544400 197510
rect -400 192946 800 192976
rect 97717 192946 97783 192949
rect -400 192944 97783 192946
rect -400 192888 97722 192944
rect 97778 192888 97783 192944
rect -400 192886 97783 192888
rect -400 192856 800 192886
rect 97717 192883 97783 192886
rect 543200 192856 544400 192976
rect -400 188232 800 188352
rect 149237 188322 149303 188325
rect 543200 188322 544400 188352
rect 149237 188320 544400 188322
rect 149237 188264 149242 188320
rect 149298 188264 544400 188320
rect 149237 188262 544400 188264
rect 149237 188259 149303 188262
rect 543200 188232 544400 188262
rect -400 183698 800 183728
rect 92197 183698 92263 183701
rect -400 183696 92263 183698
rect -400 183640 92202 183696
rect 92258 183640 92263 183696
rect -400 183638 92263 183640
rect -400 183608 800 183638
rect 92197 183635 92263 183638
rect 147397 183698 147463 183701
rect 543200 183698 544400 183728
rect 147397 183696 544400 183698
rect 147397 183640 147402 183696
rect 147458 183640 544400 183696
rect 147397 183638 544400 183640
rect 147397 183635 147463 183638
rect 543200 183608 544400 183638
rect -400 179074 800 179104
rect 1209 179074 1275 179077
rect -400 179072 1275 179074
rect -400 179016 1214 179072
rect 1270 179016 1275 179072
rect -400 179014 1275 179016
rect -400 178984 800 179014
rect 1209 179011 1275 179014
rect 543200 178984 544400 179104
rect -400 174064 800 174184
rect -400 169440 800 169560
rect -400 164816 800 164936
rect 14457 162074 14523 162077
rect 108757 162074 108823 162077
rect 14457 162072 108823 162074
rect 14457 162016 14462 162072
rect 14518 162016 108762 162072
rect 108818 162016 108823 162072
rect 14457 162014 108823 162016
rect 14457 162011 14523 162014
rect 108757 162011 108823 162014
rect -400 160192 800 160312
rect -400 155568 800 155688
rect -400 150944 800 151064
rect -400 146320 800 146440
rect 543200 125770 544400 125890
rect -400 123496 800 123616
rect 543200 121146 544400 121266
rect -400 118872 800 118992
rect 543200 116522 544400 116642
rect -400 114248 800 114368
rect 543200 111898 544400 112018
rect -400 109624 800 109744
rect 543200 107274 544400 107394
rect -400 105000 800 105120
rect 543200 102650 544400 102770
rect -400 100376 800 100496
rect 543200 98026 544400 98146
rect -400 95752 800 95872
rect 543200 93402 544400 93522
rect -400 91128 800 91248
rect 543200 88778 544400 88898
rect -400 86504 800 86624
rect 543200 84154 544400 84274
rect -400 81880 800 82000
rect 543200 79530 544400 79650
rect -400 77256 800 77376
rect 543200 74906 544400 75026
rect -400 72632 800 72752
rect 543200 70282 544400 70402
rect -400 68008 800 68128
rect 543200 65658 544400 65778
rect -400 63384 800 63504
rect 3417 62794 3483 62797
rect 112437 62794 112503 62797
rect 3417 62792 112503 62794
rect 3417 62736 3422 62792
rect 3478 62736 112442 62792
rect 112498 62736 112503 62792
rect 3417 62734 112503 62736
rect 3417 62731 3483 62734
rect 112437 62731 112503 62734
rect 104157 62114 104223 62117
rect 105077 62114 105143 62117
rect 104157 62112 105143 62114
rect 104157 62056 104162 62112
rect 104218 62056 105082 62112
rect 105138 62056 105143 62112
rect 104157 62054 105143 62056
rect 104157 62051 104223 62054
rect 105077 62051 105143 62054
rect 93117 61434 93183 61437
rect 119797 61434 119863 61437
rect 93117 61432 119863 61434
rect 93117 61376 93122 61432
rect 93178 61376 119802 61432
rect 119858 61376 119863 61432
rect 93117 61374 119863 61376
rect 93117 61371 93183 61374
rect 119797 61371 119863 61374
rect 543200 61034 544400 61154
rect 1209 60210 1275 60213
rect 94037 60210 94103 60213
rect 1209 60208 94103 60210
rect 1209 60152 1214 60208
rect 1270 60152 94042 60208
rect 94098 60152 94103 60208
rect 1209 60150 94103 60152
rect 1209 60147 1275 60150
rect 94037 60147 94103 60150
rect 117814 60148 117820 60212
rect 117884 60210 117890 60212
rect 117957 60210 118023 60213
rect 117884 60208 118023 60210
rect 117884 60152 117962 60208
rect 118018 60152 118023 60208
rect 117884 60150 118023 60152
rect 117884 60148 117890 60150
rect 117957 60147 118023 60150
rect 1025 60074 1091 60077
rect 95509 60074 95575 60077
rect 1025 60072 95575 60074
rect 1025 60016 1030 60072
rect 1086 60016 95514 60072
rect 95570 60016 95575 60072
rect 1025 60014 95575 60016
rect 1025 60011 1091 60014
rect 95509 60011 95575 60014
rect 841 59938 907 59941
rect 99557 59938 99623 59941
rect 841 59936 99623 59938
rect 841 59880 846 59936
rect 902 59880 99562 59936
rect 99618 59880 99623 59936
rect 841 59878 99623 59880
rect 841 59875 907 59878
rect 99557 59875 99623 59878
rect 115197 59938 115263 59941
rect 116117 59938 116183 59941
rect 115197 59936 116183 59938
rect 115197 59880 115202 59936
rect 115258 59880 116122 59936
rect 116178 59880 116183 59936
rect 115197 59878 116183 59880
rect 115197 59875 115263 59878
rect 116117 59875 116183 59878
rect 657 59802 723 59805
rect 103237 59802 103303 59805
rect 657 59800 103303 59802
rect 657 59744 662 59800
rect 718 59744 103242 59800
rect 103298 59744 103303 59800
rect 657 59742 103303 59744
rect 657 59739 723 59742
rect 103237 59739 103303 59742
rect 473 59666 539 59669
rect 106917 59666 106983 59669
rect 473 59664 106983 59666
rect 473 59608 478 59664
rect 534 59608 106922 59664
rect 106978 59608 106983 59664
rect 473 59606 106983 59608
rect 473 59603 539 59606
rect 106917 59603 106983 59606
rect 289 59530 355 59533
rect 110597 59530 110663 59533
rect 289 59528 110663 59530
rect 289 59472 294 59528
rect 350 59472 110602 59528
rect 110658 59472 110663 59528
rect 289 59470 110663 59472
rect 289 59467 355 59470
rect 110597 59467 110663 59470
rect 138197 59530 138263 59533
rect 543089 59530 543155 59533
rect 138197 59528 543155 59530
rect 138197 59472 138202 59528
rect 138258 59472 543094 59528
rect 543150 59472 543155 59528
rect 138197 59470 543155 59472
rect 138197 59467 138263 59470
rect 543089 59467 543155 59470
rect 105 59394 171 59397
rect 114277 59394 114343 59397
rect 105 59392 114343 59394
rect 105 59336 110 59392
rect 166 59336 114282 59392
rect 114338 59336 114343 59392
rect 105 59334 114343 59336
rect 105 59331 171 59334
rect 114277 59331 114343 59334
rect 134517 59394 134583 59397
rect 543273 59394 543339 59397
rect 134517 59392 543339 59394
rect 134517 59336 134522 59392
rect 134578 59336 543278 59392
rect 543334 59336 543339 59392
rect 134517 59334 543339 59336
rect 134517 59331 134583 59334
rect 543273 59331 543339 59334
rect -400 58760 800 58880
rect 543200 56410 544400 56530
rect -400 54136 800 54256
rect 543200 51786 544400 51906
rect -400 49512 800 49632
rect 543200 47162 544400 47282
rect 543200 42538 544400 42658
rect 543200 37914 544400 38034
rect 543200 33290 544400 33410
rect 543200 28666 544400 28786
rect 543200 24042 544400 24162
rect 108205 19818 108271 19821
rect 115105 19818 115171 19821
rect 108205 19816 115171 19818
rect 108205 19760 108210 19816
rect 108266 19760 115110 19816
rect 115166 19760 115171 19816
rect 108205 19758 115171 19760
rect 108205 19755 108271 19758
rect 115105 19755 115171 19758
rect 101765 19682 101831 19685
rect 105445 19682 105511 19685
rect 101765 19680 105511 19682
rect 101765 19624 101770 19680
rect 101826 19624 105450 19680
rect 105506 19624 105511 19680
rect 101765 19622 105511 19624
rect 101765 19619 101831 19622
rect 105445 19619 105511 19622
rect 106365 19546 106431 19549
rect 113173 19546 113239 19549
rect 106365 19544 113239 19546
rect 106365 19488 106370 19544
rect 106426 19488 113178 19544
rect 113234 19488 113239 19544
rect 106365 19486 113239 19488
rect 106365 19483 106431 19486
rect 113173 19483 113239 19486
rect 543200 19418 544400 19538
rect 100293 19412 100359 19413
rect 100293 19408 100340 19412
rect 100404 19410 100410 19412
rect 108021 19410 108087 19413
rect 151813 19412 151879 19413
rect 108430 19410 108436 19412
rect 100293 19352 100298 19408
rect 100293 19348 100340 19352
rect 100404 19350 100450 19410
rect 108021 19408 108436 19410
rect 108021 19352 108026 19408
rect 108082 19352 108436 19408
rect 108021 19350 108436 19352
rect 100404 19348 100410 19350
rect 100293 19347 100359 19348
rect 108021 19347 108087 19350
rect 108430 19348 108436 19350
rect 108500 19348 108506 19412
rect 151813 19408 151860 19412
rect 151924 19410 151930 19412
rect 151813 19352 151818 19408
rect 151813 19348 151860 19352
rect 151924 19350 151970 19410
rect 151924 19348 151930 19350
rect 151813 19347 151879 19348
rect 53097 18866 53163 18869
rect 102869 18866 102935 18869
rect 53097 18864 102935 18866
rect 53097 18808 53102 18864
rect 53158 18808 102874 18864
rect 102930 18808 102935 18864
rect 53097 18806 102935 18808
rect 53097 18803 53163 18806
rect 102869 18803 102935 18806
rect 116393 18866 116459 18869
rect 170489 18866 170555 18869
rect 116393 18864 170555 18866
rect 116393 18808 116398 18864
rect 116454 18808 170494 18864
rect 170550 18808 170555 18864
rect 116393 18806 170555 18808
rect 116393 18803 116459 18806
rect 170489 18803 170555 18806
rect 64137 18730 64203 18733
rect 121545 18730 121611 18733
rect 64137 18728 121611 18730
rect 64137 18672 64142 18728
rect 64198 18672 121550 18728
rect 121606 18672 121611 18728
rect 64137 18670 121611 18672
rect 64137 18667 64203 18670
rect 121545 18667 121611 18670
rect 129917 18730 129983 18733
rect 181437 18730 181503 18733
rect 129917 18728 181503 18730
rect 129917 18672 129922 18728
rect 129978 18672 181442 18728
rect 181498 18672 181503 18728
rect 129917 18670 181503 18672
rect 129917 18667 129983 18670
rect 181437 18667 181503 18670
rect 82905 18594 82971 18597
rect 144729 18594 144795 18597
rect 82905 18592 144795 18594
rect 82905 18536 82910 18592
rect 82966 18536 144734 18592
rect 144790 18536 144795 18592
rect 82905 18534 144795 18536
rect 82905 18531 82971 18534
rect 144729 18531 144795 18534
rect 153101 18594 153167 18597
rect 200205 18594 200271 18597
rect 153101 18592 200271 18594
rect 153101 18536 153106 18592
rect 153162 18536 200210 18592
rect 200266 18536 200271 18592
rect 153101 18534 200271 18536
rect 153101 18531 153167 18534
rect 200205 18531 200271 18534
rect 104709 18322 104775 18325
rect 111241 18322 111307 18325
rect 104709 18320 111307 18322
rect 104709 18264 104714 18320
rect 104770 18264 111246 18320
rect 111302 18264 111307 18320
rect 104709 18262 111307 18264
rect 104709 18259 104775 18262
rect 111241 18259 111307 18262
rect 109493 17506 109559 17509
rect 117037 17506 117103 17509
rect 109493 17504 117103 17506
rect 109493 17448 109498 17504
rect 109554 17448 117042 17504
rect 117098 17448 117103 17504
rect 109493 17446 117103 17448
rect 109493 17443 109559 17446
rect 117037 17443 117103 17446
rect 124121 17506 124187 17509
rect 176745 17506 176811 17509
rect 124121 17504 176811 17506
rect 124121 17448 124126 17504
rect 124182 17448 176750 17504
rect 176806 17448 176811 17504
rect 124121 17446 176811 17448
rect 124121 17443 124187 17446
rect 176745 17443 176811 17446
rect 67265 17370 67331 17373
rect 125409 17370 125475 17373
rect 67265 17368 125475 17370
rect 67265 17312 67270 17368
rect 67326 17312 125414 17368
rect 125470 17312 125475 17368
rect 67265 17310 125475 17312
rect 67265 17307 67331 17310
rect 125409 17307 125475 17310
rect 131849 17370 131915 17373
rect 183001 17370 183067 17373
rect 131849 17368 183067 17370
rect 131849 17312 131854 17368
rect 131910 17312 183006 17368
rect 183062 17312 183067 17368
rect 131849 17310 183067 17312
rect 131849 17307 131915 17310
rect 183001 17307 183067 17310
rect 86033 17234 86099 17237
rect 148593 17234 148659 17237
rect 86033 17232 148659 17234
rect 86033 17176 86038 17232
rect 86094 17176 148598 17232
rect 148654 17176 148659 17232
rect 86033 17174 148659 17176
rect 86033 17171 86099 17174
rect 148593 17171 148659 17174
rect 155033 17234 155099 17237
rect 201769 17234 201835 17237
rect 155033 17232 201835 17234
rect 155033 17176 155038 17232
rect 155094 17176 201774 17232
rect 201830 17176 201835 17232
rect 155033 17174 201835 17176
rect 155033 17171 155099 17174
rect 201769 17171 201835 17174
rect 103237 16146 103303 16149
rect 108665 16146 108731 16149
rect 103237 16144 108731 16146
rect 103237 16088 103242 16144
rect 103298 16088 108670 16144
rect 108726 16088 108731 16144
rect 103237 16086 108731 16088
rect 103237 16083 103303 16086
rect 108665 16083 108731 16086
rect 120257 16146 120323 16149
rect 173617 16146 173683 16149
rect 120257 16144 173683 16146
rect 120257 16088 120262 16144
rect 120318 16088 173622 16144
rect 173678 16088 173683 16144
rect 120257 16086 173683 16088
rect 120257 16083 120323 16086
rect 173617 16083 173683 16086
rect 68829 16010 68895 16013
rect 127341 16010 127407 16013
rect 68829 16008 127407 16010
rect 68829 15952 68834 16008
rect 68890 15952 127346 16008
rect 127402 15952 127407 16008
rect 68829 15950 127407 15952
rect 68829 15947 68895 15950
rect 127341 15947 127407 15950
rect 139577 16010 139643 16013
rect 189257 16010 189323 16013
rect 139577 16008 189323 16010
rect 139577 15952 139582 16008
rect 139638 15952 189262 16008
rect 189318 15952 189323 16008
rect 139577 15950 189323 15952
rect 139577 15947 139643 15950
rect 189257 15947 189323 15950
rect 89161 15874 89227 15877
rect 152457 15874 152523 15877
rect 89161 15872 152523 15874
rect 89161 15816 89166 15872
rect 89222 15816 152462 15872
rect 152518 15816 152523 15872
rect 89161 15814 152523 15816
rect 89161 15811 89227 15814
rect 152457 15811 152523 15814
rect 156965 15874 157031 15877
rect 203333 15874 203399 15877
rect 156965 15872 203399 15874
rect 156965 15816 156970 15872
rect 157026 15816 203338 15872
rect 203394 15816 203399 15872
rect 156965 15814 203399 15816
rect 156965 15811 157031 15814
rect 203333 15811 203399 15814
rect 112529 14786 112595 14789
rect 167361 14786 167427 14789
rect 112529 14784 167427 14786
rect 112529 14728 112534 14784
rect 112590 14728 167366 14784
rect 167422 14728 167427 14784
rect 112529 14726 167427 14728
rect 112529 14723 112595 14726
rect 167361 14723 167427 14726
rect 71957 14650 72023 14653
rect 131205 14650 131271 14653
rect 71957 14648 131271 14650
rect 71957 14592 71962 14648
rect 72018 14592 131210 14648
rect 131266 14592 131271 14648
rect 71957 14590 131271 14592
rect 71957 14587 72023 14590
rect 131205 14587 131271 14590
rect 141509 14650 141575 14653
rect 190821 14650 190887 14653
rect 141509 14648 190887 14650
rect 141509 14592 141514 14648
rect 141570 14592 190826 14648
rect 190882 14592 190887 14648
rect 141509 14590 190887 14592
rect 141509 14587 141575 14590
rect 190821 14587 190887 14590
rect 90725 14514 90791 14517
rect 154389 14514 154455 14517
rect 90725 14512 154455 14514
rect 90725 14456 90730 14512
rect 90786 14456 154394 14512
rect 154450 14456 154455 14512
rect 90725 14454 154455 14456
rect 90725 14451 90791 14454
rect 154389 14451 154455 14454
rect 114461 13290 114527 13293
rect 168925 13290 168991 13293
rect 114461 13288 168991 13290
rect 114461 13232 114466 13288
rect 114522 13232 168930 13288
rect 168986 13232 168991 13288
rect 114461 13230 168991 13232
rect 114461 13227 114527 13230
rect 168925 13227 168991 13230
rect 73521 13154 73587 13157
rect 133137 13154 133203 13157
rect 73521 13152 133203 13154
rect 73521 13096 73526 13152
rect 73582 13096 133142 13152
rect 133198 13096 133203 13152
rect 73521 13094 133203 13096
rect 73521 13091 73587 13094
rect 133137 13091 133203 13094
rect 143441 13154 143507 13157
rect 192385 13154 192451 13157
rect 143441 13152 192451 13154
rect 143441 13096 143446 13152
rect 143502 13096 192390 13152
rect 192446 13096 192451 13152
rect 143441 13094 192451 13096
rect 143441 13091 143507 13094
rect 192385 13091 192451 13094
rect 92289 13018 92355 13021
rect 156321 13018 156387 13021
rect 92289 13016 156387 13018
rect 92289 12960 92294 13016
rect 92350 12960 156326 13016
rect 156382 12960 156387 13016
rect 92289 12958 156387 12960
rect 92289 12955 92355 12958
rect 156321 12955 156387 12958
rect 122189 12066 122255 12069
rect 175181 12066 175247 12069
rect 122189 12064 175247 12066
rect 122189 12008 122194 12064
rect 122250 12008 175186 12064
rect 175242 12008 175247 12064
rect 122189 12006 175247 12008
rect 122189 12003 122255 12006
rect 175181 12003 175247 12006
rect 65701 11930 65767 11933
rect 123477 11930 123543 11933
rect 65701 11928 123543 11930
rect 65701 11872 65706 11928
rect 65762 11872 123482 11928
rect 123538 11872 123543 11928
rect 65701 11870 123543 11872
rect 65701 11867 65767 11870
rect 123477 11867 123543 11870
rect 75085 11794 75151 11797
rect 135069 11794 135135 11797
rect 75085 11792 135135 11794
rect 75085 11736 75090 11792
rect 75146 11736 135074 11792
rect 135130 11736 135135 11792
rect 75085 11734 135135 11736
rect 75085 11731 75151 11734
rect 135069 11731 135135 11734
rect 145373 11794 145439 11797
rect 193949 11794 194015 11797
rect 145373 11792 194015 11794
rect 145373 11736 145378 11792
rect 145434 11736 193954 11792
rect 194010 11736 194015 11792
rect 145373 11734 194015 11736
rect 145373 11731 145439 11734
rect 193949 11731 194015 11734
rect 95417 11658 95483 11661
rect 160185 11658 160251 11661
rect 95417 11656 160251 11658
rect 95417 11600 95422 11656
rect 95478 11600 160190 11656
rect 160246 11600 160251 11656
rect 95417 11598 160251 11600
rect 95417 11595 95483 11598
rect 160185 11595 160251 11598
rect 59445 10570 59511 10573
rect 115749 10570 115815 10573
rect 59445 10568 115815 10570
rect 59445 10512 59450 10568
rect 59506 10512 115754 10568
rect 115810 10512 115815 10568
rect 59445 10510 115815 10512
rect 59445 10507 59511 10510
rect 115749 10507 115815 10510
rect 118325 10570 118391 10573
rect 172053 10570 172119 10573
rect 118325 10568 172119 10570
rect 118325 10512 118330 10568
rect 118386 10512 172058 10568
rect 172114 10512 172119 10568
rect 118325 10510 172119 10512
rect 118325 10507 118391 10510
rect 172053 10507 172119 10510
rect 78213 10434 78279 10437
rect 138933 10434 138999 10437
rect 78213 10432 138999 10434
rect 78213 10376 78218 10432
rect 78274 10376 138938 10432
rect 138994 10376 138999 10432
rect 78213 10374 138999 10376
rect 78213 10371 78279 10374
rect 138933 10371 138999 10374
rect 149237 10434 149303 10437
rect 197077 10434 197143 10437
rect 149237 10432 197143 10434
rect 149237 10376 149242 10432
rect 149298 10376 197082 10432
rect 197138 10376 197143 10432
rect 149237 10374 197143 10376
rect 149237 10371 149303 10374
rect 197077 10371 197143 10374
rect 96981 10298 97047 10301
rect 162117 10298 162183 10301
rect 96981 10296 162183 10298
rect 96981 10240 96986 10296
rect 97042 10240 162122 10296
rect 162178 10240 162183 10296
rect 96981 10238 162183 10240
rect 96981 10235 97047 10238
rect 162117 10235 162183 10238
rect 57881 9210 57947 9213
rect 113817 9210 113883 9213
rect 57881 9208 113883 9210
rect 57881 9152 57886 9208
rect 57942 9152 113822 9208
rect 113878 9152 113883 9208
rect 57881 9150 113883 9152
rect 57881 9147 57947 9150
rect 113817 9147 113883 9150
rect 79777 9074 79843 9077
rect 140865 9074 140931 9077
rect 79777 9072 140931 9074
rect 79777 9016 79782 9072
rect 79838 9016 140870 9072
rect 140926 9016 140931 9072
rect 79777 9014 140931 9016
rect 79777 9011 79843 9014
rect 140865 9011 140931 9014
rect 151169 9074 151235 9077
rect 198641 9074 198707 9077
rect 151169 9072 198707 9074
rect 151169 9016 151174 9072
rect 151230 9016 198646 9072
rect 198702 9016 198707 9072
rect 151169 9014 198707 9016
rect 151169 9011 151235 9014
rect 198641 9011 198707 9014
rect 100109 8938 100175 8941
rect 165981 8938 166047 8941
rect 100109 8936 166047 8938
rect 100109 8880 100114 8936
rect 100170 8880 165986 8936
rect 166042 8880 166047 8936
rect 100109 8878 166047 8880
rect 100109 8875 100175 8878
rect 165981 8875 166047 8878
rect 56317 7850 56383 7853
rect 111885 7850 111951 7853
rect 56317 7848 111951 7850
rect 56317 7792 56322 7848
rect 56378 7792 111890 7848
rect 111946 7792 111951 7848
rect 56317 7790 111951 7792
rect 56317 7787 56383 7790
rect 111885 7787 111951 7790
rect 133781 7850 133847 7853
rect 184565 7850 184631 7853
rect 133781 7848 184631 7850
rect 133781 7792 133786 7848
rect 133842 7792 184570 7848
rect 184626 7792 184631 7848
rect 133781 7790 184631 7792
rect 133781 7787 133847 7790
rect 184565 7787 184631 7790
rect 106733 7714 106799 7717
rect 164233 7714 164299 7717
rect 106733 7712 164299 7714
rect 106733 7656 106738 7712
rect 106794 7656 164238 7712
rect 164294 7656 164299 7712
rect 106733 7654 164299 7656
rect 106733 7651 106799 7654
rect 164233 7651 164299 7654
rect 81341 7578 81407 7581
rect 142797 7578 142863 7581
rect 81341 7576 142863 7578
rect 81341 7520 81346 7576
rect 81402 7520 142802 7576
rect 142858 7520 142863 7576
rect 81341 7518 142863 7520
rect 81341 7515 81407 7518
rect 142797 7515 142863 7518
rect 99649 6626 99715 6629
rect 151721 6626 151787 6629
rect 99649 6624 151787 6626
rect 99649 6568 99654 6624
rect 99710 6568 151726 6624
rect 151782 6568 151787 6624
rect 99649 6566 151787 6568
rect 99649 6563 99715 6566
rect 151721 6563 151787 6566
rect 53189 6490 53255 6493
rect 106089 6490 106155 6493
rect 53189 6488 106155 6490
rect 53189 6432 53194 6488
rect 53250 6432 106094 6488
rect 106150 6432 106155 6488
rect 53189 6430 106155 6432
rect 53189 6427 53255 6430
rect 106089 6427 106155 6430
rect 103513 6354 103579 6357
rect 162669 6354 162735 6357
rect 103513 6352 162735 6354
rect 103513 6296 103518 6352
rect 103574 6296 162674 6352
rect 162730 6296 162735 6352
rect 103513 6294 162735 6296
rect 103513 6291 103579 6294
rect 162669 6291 162735 6294
rect 84469 6218 84535 6221
rect 146661 6218 146727 6221
rect 84469 6216 146727 6218
rect 84469 6160 84474 6216
rect 84530 6160 146666 6216
rect 146722 6160 146727 6216
rect 84469 6158 146727 6160
rect 84469 6155 84535 6158
rect 146661 6155 146727 6158
rect 147305 6218 147371 6221
rect 195513 6218 195579 6221
rect 147305 6216 195579 6218
rect 147305 6160 147310 6216
rect 147366 6160 195518 6216
rect 195574 6160 195579 6216
rect 147305 6158 195579 6160
rect 147305 6155 147371 6158
rect 195513 6155 195579 6158
rect 61009 5130 61075 5133
rect 117681 5130 117747 5133
rect 61009 5128 117747 5130
rect 61009 5072 61014 5128
rect 61070 5072 117686 5128
rect 117742 5072 117747 5128
rect 61009 5070 117747 5072
rect 61009 5067 61075 5070
rect 117681 5067 117747 5070
rect 76649 4994 76715 4997
rect 137001 4994 137067 4997
rect 76649 4992 137067 4994
rect 76649 4936 76654 4992
rect 76710 4936 137006 4992
rect 137062 4936 137067 4992
rect 76649 4934 137067 4936
rect 76649 4931 76715 4934
rect 137001 4931 137067 4934
rect 137645 4994 137711 4997
rect 187693 4994 187759 4997
rect 137645 4992 187759 4994
rect 137645 4936 137650 4992
rect 137706 4936 187698 4992
rect 187754 4936 187759 4992
rect 137645 4934 187759 4936
rect 137645 4931 137711 4934
rect 187693 4931 187759 4934
rect 98545 4858 98611 4861
rect 164049 4858 164115 4861
rect 98545 4856 164115 4858
rect 98545 4800 98550 4856
rect 98606 4800 164054 4856
rect 164110 4800 164115 4856
rect 98545 4798 164115 4800
rect 98545 4795 98611 4798
rect 164049 4795 164115 4798
rect 109953 3634 110019 3637
rect 165797 3634 165863 3637
rect 109953 3632 165863 3634
rect 109953 3576 109958 3632
rect 110014 3576 165802 3632
rect 165858 3576 165863 3632
rect 109953 3574 165863 3576
rect 109953 3571 110019 3574
rect 165797 3571 165863 3574
rect 70393 3498 70459 3501
rect 129273 3498 129339 3501
rect 70393 3496 129339 3498
rect 70393 3440 70398 3496
rect 70454 3440 129278 3496
rect 129334 3440 129339 3496
rect 70393 3438 129339 3440
rect 70393 3435 70459 3438
rect 129273 3435 129339 3438
rect 135713 3498 135779 3501
rect 186129 3498 186195 3501
rect 135713 3496 186195 3498
rect 135713 3440 135718 3496
rect 135774 3440 186134 3496
rect 186190 3440 186195 3496
rect 135713 3438 186195 3440
rect 135713 3435 135779 3438
rect 186129 3435 186195 3438
rect 87597 3362 87663 3365
rect 150525 3362 150591 3365
rect 87597 3360 150591 3362
rect 87597 3304 87602 3360
rect 87658 3304 150530 3360
rect 150586 3304 150591 3360
rect 87597 3302 150591 3304
rect 87597 3299 87663 3302
rect 150525 3299 150591 3302
rect 54753 2274 54819 2277
rect 109309 2274 109375 2277
rect 54753 2272 109375 2274
rect 54753 2216 54758 2272
rect 54814 2216 109314 2272
rect 109370 2216 109375 2272
rect 54753 2214 109375 2216
rect 54753 2211 54819 2214
rect 109309 2211 109375 2214
rect 127985 2274 128051 2277
rect 179873 2274 179939 2277
rect 127985 2272 179939 2274
rect 127985 2216 127990 2272
rect 128046 2216 179878 2272
rect 179934 2216 179939 2272
rect 127985 2214 179939 2216
rect 127985 2211 128051 2214
rect 179873 2211 179939 2214
rect 62573 2138 62639 2141
rect 119613 2138 119679 2141
rect 62573 2136 119679 2138
rect 62573 2080 62578 2136
rect 62634 2080 119618 2136
rect 119674 2080 119679 2136
rect 62573 2078 119679 2080
rect 62573 2075 62639 2078
rect 119613 2075 119679 2078
rect 126053 2138 126119 2141
rect 178309 2138 178375 2141
rect 126053 2136 178375 2138
rect 126053 2080 126058 2136
rect 126114 2080 178314 2136
rect 178370 2080 178375 2136
rect 126053 2078 178375 2080
rect 126053 2075 126119 2078
rect 178309 2075 178375 2078
rect 93853 2002 93919 2005
rect 158253 2002 158319 2005
rect 93853 2000 158319 2002
rect 93853 1944 93858 2000
rect 93914 1944 158258 2000
rect 158314 1944 158319 2000
rect 93853 1942 158319 1944
rect 93853 1939 93919 1942
rect 158253 1939 158319 1942
rect 51625 1322 51691 1325
rect 53097 1322 53163 1325
rect 51625 1320 53163 1322
rect 51625 1264 51630 1320
rect 51686 1264 53102 1320
rect 53158 1264 53163 1320
rect 51625 1262 53163 1264
rect 51625 1259 51691 1262
rect 53097 1259 53163 1262
rect 104157 1322 104223 1325
rect 109033 1322 109099 1325
rect 104157 1320 109099 1322
rect 104157 1264 104162 1320
rect 104218 1264 109038 1320
rect 109094 1264 109099 1320
rect 104157 1262 109099 1264
rect 104157 1259 104223 1262
rect 109033 1259 109099 1262
rect 110597 1322 110663 1325
rect 122005 1322 122071 1325
rect 132493 1322 132559 1325
rect 144085 1322 144151 1325
rect 110597 1320 113190 1322
rect 110597 1264 110602 1320
rect 110658 1264 113190 1320
rect 110597 1262 113190 1264
rect 110597 1259 110663 1262
rect 102225 1186 102291 1189
rect 111793 1186 111859 1189
rect 102225 1184 111859 1186
rect 102225 1128 102230 1184
rect 102286 1128 111798 1184
rect 111854 1128 111859 1184
rect 102225 1126 111859 1128
rect 113130 1186 113190 1262
rect 122005 1320 132559 1322
rect 122005 1264 122010 1320
rect 122066 1264 132498 1320
rect 132554 1264 132559 1320
rect 122005 1262 132559 1264
rect 122005 1259 122071 1262
rect 132493 1259 132559 1262
rect 137326 1320 144151 1322
rect 137326 1264 144090 1320
rect 144146 1264 144151 1320
rect 137326 1262 144151 1264
rect 127341 1186 127407 1189
rect 113130 1184 127407 1186
rect 113130 1128 127346 1184
rect 127402 1128 127407 1184
rect 113130 1126 127407 1128
rect 102225 1123 102291 1126
rect 111793 1123 111859 1126
rect 127341 1123 127407 1126
rect 108297 1052 108363 1053
rect 108246 1050 108252 1052
rect 108206 990 108252 1050
rect 108316 1048 108363 1052
rect 108358 992 108363 1048
rect 108246 988 108252 990
rect 108316 988 108363 992
rect 108297 987 108363 988
rect 115749 1050 115815 1053
rect 124765 1050 124831 1053
rect 115749 1048 124831 1050
rect 115749 992 115754 1048
rect 115810 992 124770 1048
rect 124826 992 124831 1048
rect 115749 990 124831 992
rect 115749 987 115815 990
rect 124765 987 124831 990
rect 131389 1050 131455 1053
rect 137326 1050 137386 1262
rect 144085 1259 144151 1262
rect 137553 1052 137619 1053
rect 131389 1048 137386 1050
rect 131389 992 131394 1048
rect 131450 992 137386 1048
rect 131389 990 137386 992
rect 131389 987 131455 990
rect 137502 988 137508 1052
rect 137572 1050 137619 1052
rect 149881 1050 149947 1053
rect 137572 1048 137664 1050
rect 137614 992 137664 1048
rect 137572 990 137664 992
rect 139166 1048 149947 1050
rect 139166 992 149886 1048
rect 149942 992 149947 1048
rect 139166 990 149947 992
rect 137572 988 137619 990
rect 137553 987 137619 988
rect 104617 914 104683 917
rect 107377 914 107443 917
rect 110413 914 110479 917
rect 104617 912 104818 914
rect 104617 856 104622 912
rect 104678 856 104818 912
rect 104617 854 104818 856
rect 104617 851 104683 854
rect 104758 778 104818 854
rect 107377 912 110479 914
rect 107377 856 107382 912
rect 107438 856 110418 912
rect 110474 856 110479 912
rect 107377 854 110479 856
rect 107377 851 107443 854
rect 110413 851 110479 854
rect 118877 914 118943 917
rect 128629 914 128695 917
rect 136357 914 136423 917
rect 118877 912 128695 914
rect 118877 856 118882 912
rect 118938 856 128634 912
rect 128690 856 128695 912
rect 118877 854 128695 856
rect 118877 851 118943 854
rect 128629 851 128695 854
rect 134382 912 136423 914
rect 134382 856 136362 912
rect 136418 856 136423 912
rect 134382 854 136423 856
rect 121453 778 121519 781
rect 104758 776 121519 778
rect 104758 720 121458 776
rect 121514 720 121519 776
rect 104758 718 121519 720
rect 121453 715 121519 718
rect 123661 778 123727 781
rect 134149 778 134215 781
rect 123661 776 134215 778
rect 123661 720 123666 776
rect 123722 720 134154 776
rect 134210 720 134215 776
rect 123661 718 134215 720
rect 123661 715 123727 718
rect 134149 715 134215 718
rect 120533 642 120599 645
rect 125225 642 125291 645
rect 134382 642 134442 854
rect 136357 851 136423 854
rect 137645 914 137711 917
rect 137870 914 137876 916
rect 137645 912 137876 914
rect 137645 856 137650 912
rect 137706 856 137876 912
rect 137645 854 137876 856
rect 137645 851 137711 854
rect 137870 852 137876 854
rect 137940 852 137946 916
rect 136173 778 136239 781
rect 139166 778 139226 990
rect 149881 987 149947 990
rect 139577 914 139643 917
rect 146017 914 146083 917
rect 139577 912 146083 914
rect 139577 856 139582 912
rect 139638 856 146022 912
rect 146078 856 146083 912
rect 139577 854 146083 856
rect 139577 851 139643 854
rect 146017 851 146083 854
rect 150157 914 150223 917
rect 167269 914 167335 917
rect 150157 912 167335 914
rect 150157 856 150162 912
rect 150218 856 167274 912
rect 167330 856 167335 912
rect 150157 854 167335 856
rect 150157 851 150223 854
rect 167269 851 167335 854
rect 136173 776 139226 778
rect 136173 720 136178 776
rect 136234 720 139226 776
rect 136173 718 139226 720
rect 139301 778 139367 781
rect 153745 778 153811 781
rect 139301 776 153811 778
rect 139301 720 139306 776
rect 139362 720 153750 776
rect 153806 720 153811 776
rect 139301 718 153811 720
rect 136173 715 136239 718
rect 139301 715 139367 718
rect 153745 715 153811 718
rect 120533 640 122850 642
rect 120533 584 120538 640
rect 120594 584 122850 640
rect 120533 582 122850 584
rect 120533 579 120599 582
rect 111149 506 111215 509
rect 119153 506 119219 509
rect 111149 504 119219 506
rect 111149 448 111154 504
rect 111210 448 119158 504
rect 119214 448 119219 504
rect 111149 446 119219 448
rect 122790 506 122850 582
rect 125225 640 134442 642
rect 125225 584 125230 640
rect 125286 584 134442 640
rect 125225 582 134442 584
rect 134609 642 134675 645
rect 147949 642 148015 645
rect 134609 640 148015 642
rect 134609 584 134614 640
rect 134670 584 147954 640
rect 148010 584 148015 640
rect 134609 582 148015 584
rect 125225 579 125291 582
rect 134609 579 134675 582
rect 147949 579 148015 582
rect 148685 642 148751 645
rect 165337 642 165403 645
rect 148685 640 165403 642
rect 148685 584 148690 640
rect 148746 584 165342 640
rect 165398 584 165403 640
rect 148685 582 165403 584
rect 148685 579 148751 582
rect 165337 579 165403 582
rect 166625 642 166691 645
rect 211245 642 211311 645
rect 166625 640 211311 642
rect 166625 584 166630 640
rect 166686 584 211250 640
rect 211306 584 211311 640
rect 166625 582 211311 584
rect 166625 579 166691 582
rect 211245 579 211311 582
rect 130561 506 130627 509
rect 122790 504 130627 506
rect 122790 448 130566 504
rect 130622 448 130627 504
rect 122790 446 130627 448
rect 111149 443 111215 446
rect 119153 443 119219 446
rect 130561 443 130627 446
rect 133045 506 133111 509
rect 139577 506 139643 509
rect 133045 504 139643 506
rect 133045 448 133050 504
rect 133106 448 139582 504
rect 139638 448 139643 504
rect 133045 446 139643 448
rect 133045 443 133111 446
rect 139577 443 139643 446
rect 140865 506 140931 509
rect 155677 506 155743 509
rect 140865 504 155743 506
rect 140865 448 140870 504
rect 140926 448 155682 504
rect 155738 448 155743 504
rect 140865 446 155743 448
rect 140865 443 140931 446
rect 155677 443 155743 446
rect 164693 506 164759 509
rect 209497 506 209563 509
rect 164693 504 209563 506
rect 164693 448 164698 504
rect 164754 448 209502 504
rect 209558 448 209563 504
rect 164693 446 209563 448
rect 164693 443 164759 446
rect 209497 443 209563 446
rect 50153 370 50219 373
rect 101397 370 101463 373
rect 50153 368 101463 370
rect 50153 312 50158 368
rect 50214 312 101402 368
rect 101458 312 101463 368
rect 50153 310 101463 312
rect 50153 307 50219 310
rect 101397 307 101463 310
rect 114277 370 114343 373
rect 122833 370 122899 373
rect 114277 368 122899 370
rect 114277 312 114282 368
rect 114338 312 122838 368
rect 122894 312 122899 368
rect 114277 310 122899 312
rect 114277 307 114343 310
rect 122833 307 122899 310
rect 128169 370 128235 373
rect 140221 370 140287 373
rect 128169 368 140287 370
rect 128169 312 128174 368
rect 128230 312 140226 368
rect 140282 312 140287 368
rect 128169 310 140287 312
rect 128169 307 128235 310
rect 140221 307 140287 310
rect 145557 370 145623 373
rect 161473 370 161539 373
rect 145557 368 161539 370
rect 145557 312 145562 368
rect 145618 312 161478 368
rect 161534 312 161539 368
rect 145557 310 161539 312
rect 145557 307 145623 310
rect 161473 307 161539 310
rect 162945 370 163011 373
rect 207933 370 207999 373
rect 162945 368 207999 370
rect 162945 312 162950 368
rect 163006 312 207938 368
rect 207994 312 207999 368
rect 162945 310 207999 312
rect 162945 307 163011 310
rect 207933 307 207999 310
rect 48589 234 48655 237
rect 100937 234 101003 237
rect 48589 232 101003 234
rect 48589 176 48594 232
rect 48650 176 100942 232
rect 100998 176 101003 232
rect 48589 174 101003 176
rect 48589 171 48655 174
rect 100937 171 101003 174
rect 117405 234 117471 237
rect 126421 234 126487 237
rect 117405 232 126487 234
rect 117405 176 117410 232
rect 117466 176 126426 232
rect 126482 176 126487 232
rect 117405 174 126487 176
rect 117405 171 117471 174
rect 126421 171 126487 174
rect 129917 234 129983 237
rect 142061 234 142127 237
rect 129917 232 142127 234
rect 129917 176 129922 232
rect 129978 176 142066 232
rect 142122 176 142127 232
rect 129917 174 142127 176
rect 129917 171 129983 174
rect 142061 171 142127 174
rect 143993 234 144059 237
rect 159817 234 159883 237
rect 143993 232 159883 234
rect 143993 176 143998 232
rect 144054 176 159822 232
rect 159878 176 159883 232
rect 143993 174 159883 176
rect 143993 171 144059 174
rect 159817 171 159883 174
rect 160829 234 160895 237
rect 206369 234 206435 237
rect 160829 232 206435 234
rect 160829 176 160834 232
rect 160890 176 206374 232
rect 206430 176 206435 232
rect 160829 174 206435 176
rect 160829 171 160895 174
rect 206369 171 206435 174
rect 47025 98 47091 101
rect 99097 98 99163 101
rect 47025 96 99163 98
rect 47025 40 47030 96
rect 47086 40 99102 96
rect 99158 40 99163 96
rect 47025 38 99163 40
rect 47025 35 47091 38
rect 99097 35 99163 38
rect 112713 98 112779 101
rect 120901 98 120967 101
rect 112713 96 120967 98
rect 112713 40 112718 96
rect 112774 40 120906 96
rect 120962 40 120967 96
rect 112713 38 120967 40
rect 112713 35 112779 38
rect 120901 35 120967 38
rect 126789 98 126855 101
rect 138289 98 138355 101
rect 126789 96 138355 98
rect 126789 40 126794 96
rect 126850 40 138294 96
rect 138350 40 138355 96
rect 126789 38 138355 40
rect 126789 35 126855 38
rect 138289 35 138355 38
rect 142429 98 142495 101
rect 157609 98 157675 101
rect 142429 96 157675 98
rect 142429 40 142434 96
rect 142490 40 157614 96
rect 157670 40 157675 96
rect 142429 38 157675 40
rect 142429 35 142495 38
rect 157609 35 157675 38
rect 158897 98 158963 101
rect 204805 98 204871 101
rect 158897 96 204871 98
rect 158897 40 158902 96
rect 158958 40 204810 96
rect 204866 40 204871 96
rect 158897 38 204871 40
rect 158897 35 158963 38
rect 204805 35 204871 38
<< via3 >>
rect 60 280468 124 280532
rect 796 239124 860 239188
rect 796 235452 860 235516
rect 117820 60148 117884 60212
rect 100340 19408 100404 19412
rect 100340 19352 100354 19408
rect 100354 19352 100404 19408
rect 100340 19348 100404 19352
rect 108436 19348 108500 19412
rect 151860 19408 151924 19412
rect 151860 19352 151874 19408
rect 151874 19352 151924 19408
rect 151860 19348 151924 19352
rect 108252 1048 108316 1052
rect 108252 992 108302 1048
rect 108302 992 108316 1048
rect 108252 988 108316 992
rect 137508 1048 137572 1052
rect 137508 992 137558 1048
rect 137558 992 137572 1048
rect 137508 988 137572 992
rect 137876 852 137940 916
<< metal4 >>
rect -4476 463972 -3856 464004
rect -4476 463736 -4444 463972
rect -4208 463736 -4124 463972
rect -3888 463736 -3856 463972
rect -4476 463652 -3856 463736
rect -4476 463416 -4444 463652
rect -4208 463416 -4124 463652
rect -3888 463416 -3856 463652
rect -4476 448614 -3856 463416
rect -4476 448378 -4444 448614
rect -4208 448378 -4124 448614
rect -3888 448378 -3856 448614
rect -4476 448294 -3856 448378
rect -4476 448058 -4444 448294
rect -4208 448058 -4124 448294
rect -3888 448058 -3856 448294
rect -4476 430614 -3856 448058
rect -4476 430378 -4444 430614
rect -4208 430378 -4124 430614
rect -3888 430378 -3856 430614
rect -4476 430294 -3856 430378
rect -4476 430058 -4444 430294
rect -4208 430058 -4124 430294
rect -3888 430058 -3856 430294
rect -4476 412614 -3856 430058
rect -4476 412378 -4444 412614
rect -4208 412378 -4124 412614
rect -3888 412378 -3856 412614
rect -4476 412294 -3856 412378
rect -4476 412058 -4444 412294
rect -4208 412058 -4124 412294
rect -3888 412058 -3856 412294
rect -4476 394614 -3856 412058
rect -4476 394378 -4444 394614
rect -4208 394378 -4124 394614
rect -3888 394378 -3856 394614
rect -4476 394294 -3856 394378
rect -4476 394058 -4444 394294
rect -4208 394058 -4124 394294
rect -3888 394058 -3856 394294
rect -4476 376614 -3856 394058
rect -4476 376378 -4444 376614
rect -4208 376378 -4124 376614
rect -3888 376378 -3856 376614
rect -4476 376294 -3856 376378
rect -4476 376058 -4444 376294
rect -4208 376058 -4124 376294
rect -3888 376058 -3856 376294
rect -4476 358614 -3856 376058
rect -4476 358378 -4444 358614
rect -4208 358378 -4124 358614
rect -3888 358378 -3856 358614
rect -4476 358294 -3856 358378
rect -4476 358058 -4444 358294
rect -4208 358058 -4124 358294
rect -3888 358058 -3856 358294
rect -4476 340614 -3856 358058
rect -4476 340378 -4444 340614
rect -4208 340378 -4124 340614
rect -3888 340378 -3856 340614
rect -4476 340294 -3856 340378
rect -4476 340058 -4444 340294
rect -4208 340058 -4124 340294
rect -3888 340058 -3856 340294
rect -4476 322614 -3856 340058
rect -4476 322378 -4444 322614
rect -4208 322378 -4124 322614
rect -3888 322378 -3856 322614
rect -4476 322294 -3856 322378
rect -4476 322058 -4444 322294
rect -4208 322058 -4124 322294
rect -3888 322058 -3856 322294
rect -4476 304614 -3856 322058
rect -4476 304378 -4444 304614
rect -4208 304378 -4124 304614
rect -3888 304378 -3856 304614
rect -4476 304294 -3856 304378
rect -4476 304058 -4444 304294
rect -4208 304058 -4124 304294
rect -3888 304058 -3856 304294
rect -4476 286614 -3856 304058
rect -4476 286378 -4444 286614
rect -4208 286378 -4124 286614
rect -3888 286378 -3856 286614
rect -4476 286294 -3856 286378
rect -4476 286058 -4444 286294
rect -4208 286058 -4124 286294
rect -3888 286058 -3856 286294
rect -4476 268614 -3856 286058
rect -4476 268378 -4444 268614
rect -4208 268378 -4124 268614
rect -3888 268378 -3856 268614
rect -4476 268294 -3856 268378
rect -4476 268058 -4444 268294
rect -4208 268058 -4124 268294
rect -3888 268058 -3856 268294
rect -4476 250614 -3856 268058
rect -4476 250378 -4444 250614
rect -4208 250378 -4124 250614
rect -3888 250378 -3856 250614
rect -4476 250294 -3856 250378
rect -4476 250058 -4444 250294
rect -4208 250058 -4124 250294
rect -3888 250058 -3856 250294
rect -4476 232614 -3856 250058
rect -4476 232378 -4444 232614
rect -4208 232378 -4124 232614
rect -3888 232378 -3856 232614
rect -4476 232294 -3856 232378
rect -4476 232058 -4444 232294
rect -4208 232058 -4124 232294
rect -3888 232058 -3856 232294
rect -4476 214614 -3856 232058
rect -4476 214378 -4444 214614
rect -4208 214378 -4124 214614
rect -3888 214378 -3856 214614
rect -4476 214294 -3856 214378
rect -4476 214058 -4444 214294
rect -4208 214058 -4124 214294
rect -3888 214058 -3856 214294
rect -4476 196614 -3856 214058
rect -4476 196378 -4444 196614
rect -4208 196378 -4124 196614
rect -3888 196378 -3856 196614
rect -4476 196294 -3856 196378
rect -4476 196058 -4444 196294
rect -4208 196058 -4124 196294
rect -3888 196058 -3856 196294
rect -4476 178614 -3856 196058
rect -4476 178378 -4444 178614
rect -4208 178378 -4124 178614
rect -3888 178378 -3856 178614
rect -4476 178294 -3856 178378
rect -4476 178058 -4444 178294
rect -4208 178058 -4124 178294
rect -3888 178058 -3856 178294
rect -4476 160614 -3856 178058
rect -4476 160378 -4444 160614
rect -4208 160378 -4124 160614
rect -3888 160378 -3856 160614
rect -4476 160294 -3856 160378
rect -4476 160058 -4444 160294
rect -4208 160058 -4124 160294
rect -3888 160058 -3856 160294
rect -4476 142614 -3856 160058
rect -4476 142378 -4444 142614
rect -4208 142378 -4124 142614
rect -3888 142378 -3856 142614
rect -4476 142294 -3856 142378
rect -4476 142058 -4444 142294
rect -4208 142058 -4124 142294
rect -3888 142058 -3856 142294
rect -4476 124614 -3856 142058
rect -4476 124378 -4444 124614
rect -4208 124378 -4124 124614
rect -3888 124378 -3856 124614
rect -4476 124294 -3856 124378
rect -4476 124058 -4444 124294
rect -4208 124058 -4124 124294
rect -3888 124058 -3856 124294
rect -4476 106614 -3856 124058
rect -4476 106378 -4444 106614
rect -4208 106378 -4124 106614
rect -3888 106378 -3856 106614
rect -4476 106294 -3856 106378
rect -4476 106058 -4444 106294
rect -4208 106058 -4124 106294
rect -3888 106058 -3856 106294
rect -4476 88614 -3856 106058
rect -4476 88378 -4444 88614
rect -4208 88378 -4124 88614
rect -3888 88378 -3856 88614
rect -4476 88294 -3856 88378
rect -4476 88058 -4444 88294
rect -4208 88058 -4124 88294
rect -3888 88058 -3856 88294
rect -4476 70614 -3856 88058
rect -4476 70378 -4444 70614
rect -4208 70378 -4124 70614
rect -3888 70378 -3856 70614
rect -4476 70294 -3856 70378
rect -4476 70058 -4444 70294
rect -4208 70058 -4124 70294
rect -3888 70058 -3856 70294
rect -4476 52614 -3856 70058
rect -4476 52378 -4444 52614
rect -4208 52378 -4124 52614
rect -3888 52378 -3856 52614
rect -4476 52294 -3856 52378
rect -4476 52058 -4444 52294
rect -4208 52058 -4124 52294
rect -3888 52058 -3856 52294
rect -4476 34614 -3856 52058
rect -4476 34378 -4444 34614
rect -4208 34378 -4124 34614
rect -3888 34378 -3856 34614
rect -4476 34294 -3856 34378
rect -4476 34058 -4444 34294
rect -4208 34058 -4124 34294
rect -3888 34058 -3856 34294
rect -4476 16614 -3856 34058
rect -4476 16378 -4444 16614
rect -4208 16378 -4124 16614
rect -3888 16378 -3856 16614
rect -4476 16294 -3856 16378
rect -4476 16058 -4444 16294
rect -4208 16058 -4124 16294
rect -3888 16058 -3856 16294
rect -4476 -3736 -3856 16058
rect -3516 463012 -2896 463044
rect -3516 462776 -3484 463012
rect -3248 462776 -3164 463012
rect -2928 462776 -2896 463012
rect -3516 462692 -2896 462776
rect -3516 462456 -3484 462692
rect -3248 462456 -3164 462692
rect -2928 462456 -2896 462692
rect -3516 444894 -2896 462456
rect -3516 444658 -3484 444894
rect -3248 444658 -3164 444894
rect -2928 444658 -2896 444894
rect -3516 444574 -2896 444658
rect -3516 444338 -3484 444574
rect -3248 444338 -3164 444574
rect -2928 444338 -2896 444574
rect -3516 426894 -2896 444338
rect -3516 426658 -3484 426894
rect -3248 426658 -3164 426894
rect -2928 426658 -2896 426894
rect -3516 426574 -2896 426658
rect -3516 426338 -3484 426574
rect -3248 426338 -3164 426574
rect -2928 426338 -2896 426574
rect -3516 408894 -2896 426338
rect -3516 408658 -3484 408894
rect -3248 408658 -3164 408894
rect -2928 408658 -2896 408894
rect -3516 408574 -2896 408658
rect -3516 408338 -3484 408574
rect -3248 408338 -3164 408574
rect -2928 408338 -2896 408574
rect -3516 390894 -2896 408338
rect -3516 390658 -3484 390894
rect -3248 390658 -3164 390894
rect -2928 390658 -2896 390894
rect -3516 390574 -2896 390658
rect -3516 390338 -3484 390574
rect -3248 390338 -3164 390574
rect -2928 390338 -2896 390574
rect -3516 372894 -2896 390338
rect -3516 372658 -3484 372894
rect -3248 372658 -3164 372894
rect -2928 372658 -2896 372894
rect -3516 372574 -2896 372658
rect -3516 372338 -3484 372574
rect -3248 372338 -3164 372574
rect -2928 372338 -2896 372574
rect -3516 354894 -2896 372338
rect -3516 354658 -3484 354894
rect -3248 354658 -3164 354894
rect -2928 354658 -2896 354894
rect -3516 354574 -2896 354658
rect -3516 354338 -3484 354574
rect -3248 354338 -3164 354574
rect -2928 354338 -2896 354574
rect -3516 336894 -2896 354338
rect -3516 336658 -3484 336894
rect -3248 336658 -3164 336894
rect -2928 336658 -2896 336894
rect -3516 336574 -2896 336658
rect -3516 336338 -3484 336574
rect -3248 336338 -3164 336574
rect -2928 336338 -2896 336574
rect -3516 318894 -2896 336338
rect -3516 318658 -3484 318894
rect -3248 318658 -3164 318894
rect -2928 318658 -2896 318894
rect -3516 318574 -2896 318658
rect -3516 318338 -3484 318574
rect -3248 318338 -3164 318574
rect -2928 318338 -2896 318574
rect -3516 300894 -2896 318338
rect -3516 300658 -3484 300894
rect -3248 300658 -3164 300894
rect -2928 300658 -2896 300894
rect -3516 300574 -2896 300658
rect -3516 300338 -3484 300574
rect -3248 300338 -3164 300574
rect -2928 300338 -2896 300574
rect -3516 282894 -2896 300338
rect -3516 282658 -3484 282894
rect -3248 282658 -3164 282894
rect -2928 282658 -2896 282894
rect -3516 282574 -2896 282658
rect -3516 282338 -3484 282574
rect -3248 282338 -3164 282574
rect -2928 282338 -2896 282574
rect -3516 264894 -2896 282338
rect -3516 264658 -3484 264894
rect -3248 264658 -3164 264894
rect -2928 264658 -2896 264894
rect -3516 264574 -2896 264658
rect -3516 264338 -3484 264574
rect -3248 264338 -3164 264574
rect -2928 264338 -2896 264574
rect -3516 246894 -2896 264338
rect -3516 246658 -3484 246894
rect -3248 246658 -3164 246894
rect -2928 246658 -2896 246894
rect -3516 246574 -2896 246658
rect -3516 246338 -3484 246574
rect -3248 246338 -3164 246574
rect -2928 246338 -2896 246574
rect -3516 228894 -2896 246338
rect -3516 228658 -3484 228894
rect -3248 228658 -3164 228894
rect -2928 228658 -2896 228894
rect -3516 228574 -2896 228658
rect -3516 228338 -3484 228574
rect -3248 228338 -3164 228574
rect -2928 228338 -2896 228574
rect -3516 210894 -2896 228338
rect -3516 210658 -3484 210894
rect -3248 210658 -3164 210894
rect -2928 210658 -2896 210894
rect -3516 210574 -2896 210658
rect -3516 210338 -3484 210574
rect -3248 210338 -3164 210574
rect -2928 210338 -2896 210574
rect -3516 192894 -2896 210338
rect -3516 192658 -3484 192894
rect -3248 192658 -3164 192894
rect -2928 192658 -2896 192894
rect -3516 192574 -2896 192658
rect -3516 192338 -3484 192574
rect -3248 192338 -3164 192574
rect -2928 192338 -2896 192574
rect -3516 174894 -2896 192338
rect -3516 174658 -3484 174894
rect -3248 174658 -3164 174894
rect -2928 174658 -2896 174894
rect -3516 174574 -2896 174658
rect -3516 174338 -3484 174574
rect -3248 174338 -3164 174574
rect -2928 174338 -2896 174574
rect -3516 156894 -2896 174338
rect -3516 156658 -3484 156894
rect -3248 156658 -3164 156894
rect -2928 156658 -2896 156894
rect -3516 156574 -2896 156658
rect -3516 156338 -3484 156574
rect -3248 156338 -3164 156574
rect -2928 156338 -2896 156574
rect -3516 138894 -2896 156338
rect -3516 138658 -3484 138894
rect -3248 138658 -3164 138894
rect -2928 138658 -2896 138894
rect -3516 138574 -2896 138658
rect -3516 138338 -3484 138574
rect -3248 138338 -3164 138574
rect -2928 138338 -2896 138574
rect -3516 120894 -2896 138338
rect -3516 120658 -3484 120894
rect -3248 120658 -3164 120894
rect -2928 120658 -2896 120894
rect -3516 120574 -2896 120658
rect -3516 120338 -3484 120574
rect -3248 120338 -3164 120574
rect -2928 120338 -2896 120574
rect -3516 102894 -2896 120338
rect -3516 102658 -3484 102894
rect -3248 102658 -3164 102894
rect -2928 102658 -2896 102894
rect -3516 102574 -2896 102658
rect -3516 102338 -3484 102574
rect -3248 102338 -3164 102574
rect -2928 102338 -2896 102574
rect -3516 84894 -2896 102338
rect -3516 84658 -3484 84894
rect -3248 84658 -3164 84894
rect -2928 84658 -2896 84894
rect -3516 84574 -2896 84658
rect -3516 84338 -3484 84574
rect -3248 84338 -3164 84574
rect -2928 84338 -2896 84574
rect -3516 66894 -2896 84338
rect -3516 66658 -3484 66894
rect -3248 66658 -3164 66894
rect -2928 66658 -2896 66894
rect -3516 66574 -2896 66658
rect -3516 66338 -3484 66574
rect -3248 66338 -3164 66574
rect -2928 66338 -2896 66574
rect -3516 48894 -2896 66338
rect -3516 48658 -3484 48894
rect -3248 48658 -3164 48894
rect -2928 48658 -2896 48894
rect -3516 48574 -2896 48658
rect -3516 48338 -3484 48574
rect -3248 48338 -3164 48574
rect -2928 48338 -2896 48574
rect -3516 30894 -2896 48338
rect -3516 30658 -3484 30894
rect -3248 30658 -3164 30894
rect -2928 30658 -2896 30894
rect -3516 30574 -2896 30658
rect -3516 30338 -3484 30574
rect -3248 30338 -3164 30574
rect -2928 30338 -2896 30574
rect -3516 12894 -2896 30338
rect -3516 12658 -3484 12894
rect -3248 12658 -3164 12894
rect -2928 12658 -2896 12894
rect -3516 12574 -2896 12658
rect -3516 12338 -3484 12574
rect -3248 12338 -3164 12574
rect -2928 12338 -2896 12574
rect -3516 -2776 -2896 12338
rect -2556 462052 -1936 462084
rect -2556 461816 -2524 462052
rect -2288 461816 -2204 462052
rect -1968 461816 -1936 462052
rect -2556 461732 -1936 461816
rect -2556 461496 -2524 461732
rect -2288 461496 -2204 461732
rect -1968 461496 -1936 461732
rect -2556 441174 -1936 461496
rect -2556 440938 -2524 441174
rect -2288 440938 -2204 441174
rect -1968 440938 -1936 441174
rect -2556 440854 -1936 440938
rect -2556 440618 -2524 440854
rect -2288 440618 -2204 440854
rect -1968 440618 -1936 440854
rect -2556 423174 -1936 440618
rect -2556 422938 -2524 423174
rect -2288 422938 -2204 423174
rect -1968 422938 -1936 423174
rect -2556 422854 -1936 422938
rect -2556 422618 -2524 422854
rect -2288 422618 -2204 422854
rect -1968 422618 -1936 422854
rect -2556 405174 -1936 422618
rect -2556 404938 -2524 405174
rect -2288 404938 -2204 405174
rect -1968 404938 -1936 405174
rect -2556 404854 -1936 404938
rect -2556 404618 -2524 404854
rect -2288 404618 -2204 404854
rect -1968 404618 -1936 404854
rect -2556 387174 -1936 404618
rect -2556 386938 -2524 387174
rect -2288 386938 -2204 387174
rect -1968 386938 -1936 387174
rect -2556 386854 -1936 386938
rect -2556 386618 -2524 386854
rect -2288 386618 -2204 386854
rect -1968 386618 -1936 386854
rect -2556 369174 -1936 386618
rect -2556 368938 -2524 369174
rect -2288 368938 -2204 369174
rect -1968 368938 -1936 369174
rect -2556 368854 -1936 368938
rect -2556 368618 -2524 368854
rect -2288 368618 -2204 368854
rect -1968 368618 -1936 368854
rect -2556 351174 -1936 368618
rect -2556 350938 -2524 351174
rect -2288 350938 -2204 351174
rect -1968 350938 -1936 351174
rect -2556 350854 -1936 350938
rect -2556 350618 -2524 350854
rect -2288 350618 -2204 350854
rect -1968 350618 -1936 350854
rect -2556 333174 -1936 350618
rect -2556 332938 -2524 333174
rect -2288 332938 -2204 333174
rect -1968 332938 -1936 333174
rect -2556 332854 -1936 332938
rect -2556 332618 -2524 332854
rect -2288 332618 -2204 332854
rect -1968 332618 -1936 332854
rect -2556 315174 -1936 332618
rect -2556 314938 -2524 315174
rect -2288 314938 -2204 315174
rect -1968 314938 -1936 315174
rect -2556 314854 -1936 314938
rect -2556 314618 -2524 314854
rect -2288 314618 -2204 314854
rect -1968 314618 -1936 314854
rect -2556 297174 -1936 314618
rect -2556 296938 -2524 297174
rect -2288 296938 -2204 297174
rect -1968 296938 -1936 297174
rect -2556 296854 -1936 296938
rect -2556 296618 -2524 296854
rect -2288 296618 -2204 296854
rect -1968 296618 -1936 296854
rect -2556 279174 -1936 296618
rect -2556 278938 -2524 279174
rect -2288 278938 -2204 279174
rect -1968 278938 -1936 279174
rect -2556 278854 -1936 278938
rect -2556 278618 -2524 278854
rect -2288 278618 -2204 278854
rect -1968 278618 -1936 278854
rect -2556 261174 -1936 278618
rect -2556 260938 -2524 261174
rect -2288 260938 -2204 261174
rect -1968 260938 -1936 261174
rect -2556 260854 -1936 260938
rect -2556 260618 -2524 260854
rect -2288 260618 -2204 260854
rect -1968 260618 -1936 260854
rect -2556 243174 -1936 260618
rect -2556 242938 -2524 243174
rect -2288 242938 -2204 243174
rect -1968 242938 -1936 243174
rect -2556 242854 -1936 242938
rect -2556 242618 -2524 242854
rect -2288 242618 -2204 242854
rect -1968 242618 -1936 242854
rect -2556 225174 -1936 242618
rect -2556 224938 -2524 225174
rect -2288 224938 -2204 225174
rect -1968 224938 -1936 225174
rect -2556 224854 -1936 224938
rect -2556 224618 -2524 224854
rect -2288 224618 -2204 224854
rect -1968 224618 -1936 224854
rect -2556 207174 -1936 224618
rect -2556 206938 -2524 207174
rect -2288 206938 -2204 207174
rect -1968 206938 -1936 207174
rect -2556 206854 -1936 206938
rect -2556 206618 -2524 206854
rect -2288 206618 -2204 206854
rect -1968 206618 -1936 206854
rect -2556 189174 -1936 206618
rect -2556 188938 -2524 189174
rect -2288 188938 -2204 189174
rect -1968 188938 -1936 189174
rect -2556 188854 -1936 188938
rect -2556 188618 -2524 188854
rect -2288 188618 -2204 188854
rect -1968 188618 -1936 188854
rect -2556 171174 -1936 188618
rect -2556 170938 -2524 171174
rect -2288 170938 -2204 171174
rect -1968 170938 -1936 171174
rect -2556 170854 -1936 170938
rect -2556 170618 -2524 170854
rect -2288 170618 -2204 170854
rect -1968 170618 -1936 170854
rect -2556 153174 -1936 170618
rect -2556 152938 -2524 153174
rect -2288 152938 -2204 153174
rect -1968 152938 -1936 153174
rect -2556 152854 -1936 152938
rect -2556 152618 -2524 152854
rect -2288 152618 -2204 152854
rect -1968 152618 -1936 152854
rect -2556 135174 -1936 152618
rect -2556 134938 -2524 135174
rect -2288 134938 -2204 135174
rect -1968 134938 -1936 135174
rect -2556 134854 -1936 134938
rect -2556 134618 -2524 134854
rect -2288 134618 -2204 134854
rect -1968 134618 -1936 134854
rect -2556 117174 -1936 134618
rect -2556 116938 -2524 117174
rect -2288 116938 -2204 117174
rect -1968 116938 -1936 117174
rect -2556 116854 -1936 116938
rect -2556 116618 -2524 116854
rect -2288 116618 -2204 116854
rect -1968 116618 -1936 116854
rect -2556 99174 -1936 116618
rect -2556 98938 -2524 99174
rect -2288 98938 -2204 99174
rect -1968 98938 -1936 99174
rect -2556 98854 -1936 98938
rect -2556 98618 -2524 98854
rect -2288 98618 -2204 98854
rect -1968 98618 -1936 98854
rect -2556 81174 -1936 98618
rect -2556 80938 -2524 81174
rect -2288 80938 -2204 81174
rect -1968 80938 -1936 81174
rect -2556 80854 -1936 80938
rect -2556 80618 -2524 80854
rect -2288 80618 -2204 80854
rect -1968 80618 -1936 80854
rect -2556 63174 -1936 80618
rect -2556 62938 -2524 63174
rect -2288 62938 -2204 63174
rect -1968 62938 -1936 63174
rect -2556 62854 -1936 62938
rect -2556 62618 -2524 62854
rect -2288 62618 -2204 62854
rect -1968 62618 -1936 62854
rect -2556 45174 -1936 62618
rect -2556 44938 -2524 45174
rect -2288 44938 -2204 45174
rect -1968 44938 -1936 45174
rect -2556 44854 -1936 44938
rect -2556 44618 -2524 44854
rect -2288 44618 -2204 44854
rect -1968 44618 -1936 44854
rect -2556 27174 -1936 44618
rect -2556 26938 -2524 27174
rect -2288 26938 -2204 27174
rect -1968 26938 -1936 27174
rect -2556 26854 -1936 26938
rect -2556 26618 -2524 26854
rect -2288 26618 -2204 26854
rect -1968 26618 -1936 26854
rect -2556 9174 -1936 26618
rect -2556 8938 -2524 9174
rect -2288 8938 -2204 9174
rect -1968 8938 -1936 9174
rect -2556 8854 -1936 8938
rect -2556 8618 -2524 8854
rect -2288 8618 -2204 8854
rect -1968 8618 -1936 8854
rect -2556 -1816 -1936 8618
rect -1596 461092 -976 461124
rect -1596 460856 -1564 461092
rect -1328 460856 -1244 461092
rect -1008 460856 -976 461092
rect -1596 460772 -976 460856
rect -1596 460536 -1564 460772
rect -1328 460536 -1244 460772
rect -1008 460536 -976 460772
rect -1596 455454 -976 460536
rect -1596 455218 -1564 455454
rect -1328 455218 -1244 455454
rect -1008 455218 -976 455454
rect -1596 455134 -976 455218
rect -1596 454898 -1564 455134
rect -1328 454898 -1244 455134
rect -1008 454898 -976 455134
rect -1596 437454 -976 454898
rect -1596 437218 -1564 437454
rect -1328 437218 -1244 437454
rect -1008 437218 -976 437454
rect -1596 437134 -976 437218
rect -1596 436898 -1564 437134
rect -1328 436898 -1244 437134
rect -1008 436898 -976 437134
rect -1596 419454 -976 436898
rect -1596 419218 -1564 419454
rect -1328 419218 -1244 419454
rect -1008 419218 -976 419454
rect -1596 419134 -976 419218
rect -1596 418898 -1564 419134
rect -1328 418898 -1244 419134
rect -1008 418898 -976 419134
rect -1596 401454 -976 418898
rect -1596 401218 -1564 401454
rect -1328 401218 -1244 401454
rect -1008 401218 -976 401454
rect -1596 401134 -976 401218
rect -1596 400898 -1564 401134
rect -1328 400898 -1244 401134
rect -1008 400898 -976 401134
rect -1596 383454 -976 400898
rect -1596 383218 -1564 383454
rect -1328 383218 -1244 383454
rect -1008 383218 -976 383454
rect -1596 383134 -976 383218
rect -1596 382898 -1564 383134
rect -1328 382898 -1244 383134
rect -1008 382898 -976 383134
rect -1596 365454 -976 382898
rect -1596 365218 -1564 365454
rect -1328 365218 -1244 365454
rect -1008 365218 -976 365454
rect -1596 365134 -976 365218
rect -1596 364898 -1564 365134
rect -1328 364898 -1244 365134
rect -1008 364898 -976 365134
rect -1596 347454 -976 364898
rect -1596 347218 -1564 347454
rect -1328 347218 -1244 347454
rect -1008 347218 -976 347454
rect -1596 347134 -976 347218
rect -1596 346898 -1564 347134
rect -1328 346898 -1244 347134
rect -1008 346898 -976 347134
rect -1596 329454 -976 346898
rect -1596 329218 -1564 329454
rect -1328 329218 -1244 329454
rect -1008 329218 -976 329454
rect -1596 329134 -976 329218
rect -1596 328898 -1564 329134
rect -1328 328898 -1244 329134
rect -1008 328898 -976 329134
rect -1596 311454 -976 328898
rect -1596 311218 -1564 311454
rect -1328 311218 -1244 311454
rect -1008 311218 -976 311454
rect -1596 311134 -976 311218
rect -1596 310898 -1564 311134
rect -1328 310898 -1244 311134
rect -1008 310898 -976 311134
rect -1596 293454 -976 310898
rect -1596 293218 -1564 293454
rect -1328 293218 -1244 293454
rect -1008 293218 -976 293454
rect -1596 293134 -976 293218
rect -1596 292898 -1564 293134
rect -1328 292898 -1244 293134
rect -1008 292898 -976 293134
rect -1596 275454 -976 292898
rect 4714 461092 5334 464004
rect 4714 460856 4746 461092
rect 4982 460856 5066 461092
rect 5302 460856 5334 461092
rect 4714 460772 5334 460856
rect 4714 460536 4746 460772
rect 4982 460536 5066 460772
rect 5302 460536 5334 460772
rect 4714 455454 5334 460536
rect 4714 455218 4746 455454
rect 4982 455218 5066 455454
rect 5302 455218 5334 455454
rect 4714 455134 5334 455218
rect 4714 454898 4746 455134
rect 4982 454898 5066 455134
rect 5302 454898 5334 455134
rect 4714 437454 5334 454898
rect 4714 437218 4746 437454
rect 4982 437218 5066 437454
rect 5302 437218 5334 437454
rect 4714 437134 5334 437218
rect 4714 436898 4746 437134
rect 4982 436898 5066 437134
rect 5302 436898 5334 437134
rect 4714 419454 5334 436898
rect 4714 419218 4746 419454
rect 4982 419218 5066 419454
rect 5302 419218 5334 419454
rect 4714 419134 5334 419218
rect 4714 418898 4746 419134
rect 4982 418898 5066 419134
rect 5302 418898 5334 419134
rect 4714 401454 5334 418898
rect 4714 401218 4746 401454
rect 4982 401218 5066 401454
rect 5302 401218 5334 401454
rect 4714 401134 5334 401218
rect 4714 400898 4746 401134
rect 4982 400898 5066 401134
rect 5302 400898 5334 401134
rect 4714 383454 5334 400898
rect 4714 383218 4746 383454
rect 4982 383218 5066 383454
rect 5302 383218 5334 383454
rect 4714 383134 5334 383218
rect 4714 382898 4746 383134
rect 4982 382898 5066 383134
rect 5302 382898 5334 383134
rect 4714 365454 5334 382898
rect 4714 365218 4746 365454
rect 4982 365218 5066 365454
rect 5302 365218 5334 365454
rect 4714 365134 5334 365218
rect 4714 364898 4746 365134
rect 4982 364898 5066 365134
rect 5302 364898 5334 365134
rect 4714 347454 5334 364898
rect 4714 347218 4746 347454
rect 4982 347218 5066 347454
rect 5302 347218 5334 347454
rect 4714 347134 5334 347218
rect 4714 346898 4746 347134
rect 4982 346898 5066 347134
rect 5302 346898 5334 347134
rect 4714 329454 5334 346898
rect 4714 329218 4746 329454
rect 4982 329218 5066 329454
rect 5302 329218 5334 329454
rect 4714 329134 5334 329218
rect 4714 328898 4746 329134
rect 4982 328898 5066 329134
rect 5302 328898 5334 329134
rect 4714 311454 5334 328898
rect 4714 311218 4746 311454
rect 4982 311218 5066 311454
rect 5302 311218 5334 311454
rect 4714 311134 5334 311218
rect 4714 310898 4746 311134
rect 4982 310898 5066 311134
rect 5302 310898 5334 311134
rect 4714 293454 5334 310898
rect 4714 293218 4746 293454
rect 4982 293218 5066 293454
rect 5302 293218 5334 293454
rect 4714 293134 5334 293218
rect 4714 292898 4746 293134
rect 4982 292898 5066 293134
rect 5302 292898 5334 293134
rect 59 280532 125 280533
rect 59 280468 60 280532
rect 124 280468 125 280532
rect 59 280467 125 280468
rect -1596 275218 -1564 275454
rect -1328 275218 -1244 275454
rect -1008 275218 -976 275454
rect -1596 275134 -976 275218
rect -1596 274898 -1564 275134
rect -1328 274898 -1244 275134
rect -1008 274898 -976 275134
rect -1596 257454 -976 274898
rect -1596 257218 -1564 257454
rect -1328 257218 -1244 257454
rect -1008 257218 -976 257454
rect -1596 257134 -976 257218
rect -1596 256898 -1564 257134
rect -1328 256898 -1244 257134
rect -1008 256898 -976 257134
rect -1596 239454 -976 256898
rect -1596 239218 -1564 239454
rect -1328 239218 -1244 239454
rect -1008 239218 -976 239454
rect -1596 239134 -976 239218
rect -1596 238898 -1564 239134
rect -1328 238898 -1244 239134
rect -1008 238898 -976 239134
rect -1596 221454 -976 238898
rect -1596 221218 -1564 221454
rect -1328 221218 -1244 221454
rect -1008 221218 -976 221454
rect -1596 221134 -976 221218
rect -1596 220898 -1564 221134
rect -1328 220898 -1244 221134
rect -1008 220898 -976 221134
rect -1596 203454 -976 220898
rect -1596 203218 -1564 203454
rect -1328 203218 -1244 203454
rect -1008 203218 -976 203454
rect -1596 203134 -976 203218
rect -1596 202898 -1564 203134
rect -1328 202898 -1244 203134
rect -1008 202898 -976 203134
rect -1596 185454 -976 202898
rect -1596 185218 -1564 185454
rect -1328 185218 -1244 185454
rect -1008 185218 -976 185454
rect -1596 185134 -976 185218
rect -1596 184898 -1564 185134
rect -1328 184898 -1244 185134
rect -1008 184898 -976 185134
rect -1596 167454 -976 184898
rect -1596 167218 -1564 167454
rect -1328 167218 -1244 167454
rect -1008 167218 -976 167454
rect -1596 167134 -976 167218
rect -1596 166898 -1564 167134
rect -1328 166898 -1244 167134
rect -1008 166898 -976 167134
rect -1596 149454 -976 166898
rect -1596 149218 -1564 149454
rect -1328 149218 -1244 149454
rect -1008 149218 -976 149454
rect -1596 149134 -976 149218
rect -1596 148898 -1564 149134
rect -1328 148898 -1244 149134
rect -1008 148898 -976 149134
rect -1596 131454 -976 148898
rect -1596 131218 -1564 131454
rect -1328 131218 -1244 131454
rect -1008 131218 -976 131454
rect -1596 131134 -976 131218
rect -1596 130898 -1564 131134
rect -1328 130898 -1244 131134
rect -1008 130898 -976 131134
rect -1596 113454 -976 130898
rect -1596 113218 -1564 113454
rect -1328 113218 -1244 113454
rect -1008 113218 -976 113454
rect -1596 113134 -976 113218
rect -1596 112898 -1564 113134
rect -1328 112898 -1244 113134
rect -1008 112898 -976 113134
rect -1596 95454 -976 112898
rect -1596 95218 -1564 95454
rect -1328 95218 -1244 95454
rect -1008 95218 -976 95454
rect -1596 95134 -976 95218
rect -1596 94898 -1564 95134
rect -1328 94898 -1244 95134
rect -1008 94898 -976 95134
rect -1596 77454 -976 94898
rect -1596 77218 -1564 77454
rect -1328 77218 -1244 77454
rect -1008 77218 -976 77454
rect -1596 77134 -976 77218
rect -1596 76898 -1564 77134
rect -1328 76898 -1244 77134
rect -1008 76898 -976 77134
rect -1596 59454 -976 76898
rect 62 74550 122 280467
rect 4714 275454 5334 292898
rect 4714 275218 4746 275454
rect 4982 275218 5066 275454
rect 5302 275218 5334 275454
rect 4714 275134 5334 275218
rect 4714 274898 4746 275134
rect 4982 274898 5066 275134
rect 5302 274898 5334 275134
rect 4714 257454 5334 274898
rect 4714 257218 4746 257454
rect 4982 257218 5066 257454
rect 5302 257218 5334 257454
rect 4714 257134 5334 257218
rect 4714 256898 4746 257134
rect 4982 256898 5066 257134
rect 5302 256898 5334 257134
rect 4714 239454 5334 256898
rect 4714 239218 4746 239454
rect 4982 239218 5066 239454
rect 5302 239218 5334 239454
rect 795 239188 861 239189
rect 795 239124 796 239188
rect 860 239124 861 239188
rect 795 239123 861 239124
rect 4714 239134 5334 239218
rect 798 235517 858 239123
rect 4714 238898 4746 239134
rect 4982 238898 5066 239134
rect 5302 238898 5334 239134
rect 795 235516 861 235517
rect 795 235452 796 235516
rect 860 235452 861 235516
rect 795 235451 861 235452
rect 4714 221454 5334 238898
rect 4714 221218 4746 221454
rect 4982 221218 5066 221454
rect 5302 221218 5334 221454
rect 4714 221134 5334 221218
rect 4714 220898 4746 221134
rect 4982 220898 5066 221134
rect 5302 220898 5334 221134
rect 4714 203454 5334 220898
rect 4714 203218 4746 203454
rect 4982 203218 5066 203454
rect 5302 203218 5334 203454
rect 4714 203134 5334 203218
rect 4714 202898 4746 203134
rect 4982 202898 5066 203134
rect 5302 202898 5334 203134
rect 4714 185454 5334 202898
rect 4714 185218 4746 185454
rect 4982 185218 5066 185454
rect 5302 185218 5334 185454
rect 4714 185134 5334 185218
rect 4714 184898 4746 185134
rect 4982 184898 5066 185134
rect 5302 184898 5334 185134
rect 4714 167454 5334 184898
rect 4714 167218 4746 167454
rect 4982 167218 5066 167454
rect 5302 167218 5334 167454
rect 4714 167134 5334 167218
rect 4714 166898 4746 167134
rect 4982 166898 5066 167134
rect 5302 166898 5334 167134
rect 4714 149454 5334 166898
rect 4714 149218 4746 149454
rect 4982 149218 5066 149454
rect 5302 149218 5334 149454
rect 4714 149134 5334 149218
rect 4714 148898 4746 149134
rect 4982 148898 5066 149134
rect 5302 148898 5334 149134
rect 4714 131454 5334 148898
rect 4714 131218 4746 131454
rect 4982 131218 5066 131454
rect 5302 131218 5334 131454
rect 4714 131134 5334 131218
rect 4714 130898 4746 131134
rect 4982 130898 5066 131134
rect 5302 130898 5334 131134
rect 4714 113454 5334 130898
rect 4714 113218 4746 113454
rect 4982 113218 5066 113454
rect 5302 113218 5334 113454
rect 4714 113134 5334 113218
rect 4714 112898 4746 113134
rect 4982 112898 5066 113134
rect 5302 112898 5334 113134
rect 4714 95454 5334 112898
rect 4714 95218 4746 95454
rect 4982 95218 5066 95454
rect 5302 95218 5334 95454
rect 4714 95134 5334 95218
rect 4714 94898 4746 95134
rect 4982 94898 5066 95134
rect 5302 94898 5334 95134
rect 4714 77454 5334 94898
rect 4714 77218 4746 77454
rect 4982 77218 5066 77454
rect 5302 77218 5334 77454
rect 4714 77134 5334 77218
rect 4714 76898 4746 77134
rect 4982 76898 5066 77134
rect 5302 76898 5334 77134
rect 62 74490 306 74550
rect 246 60298 306 74490
rect -1596 59218 -1564 59454
rect -1328 59218 -1244 59454
rect -1008 59218 -976 59454
rect -1596 59134 -976 59218
rect -1596 58898 -1564 59134
rect -1328 58898 -1244 59134
rect -1008 58898 -976 59134
rect -1596 41454 -976 58898
rect -1596 41218 -1564 41454
rect -1328 41218 -1244 41454
rect -1008 41218 -976 41454
rect -1596 41134 -976 41218
rect -1596 40898 -1564 41134
rect -1328 40898 -1244 41134
rect -1008 40898 -976 41134
rect -1596 23454 -976 40898
rect -1596 23218 -1564 23454
rect -1328 23218 -1244 23454
rect -1008 23218 -976 23454
rect -1596 23134 -976 23218
rect -1596 22898 -1564 23134
rect -1328 22898 -1244 23134
rect -1008 22898 -976 23134
rect -1596 5454 -976 22898
rect -1596 5218 -1564 5454
rect -1328 5218 -1244 5454
rect -1008 5218 -976 5454
rect -1596 5134 -976 5218
rect -1596 4898 -1564 5134
rect -1328 4898 -1244 5134
rect -1008 4898 -976 5134
rect -1596 -856 -976 4898
rect 4714 59454 5334 76898
rect 4714 59218 4746 59454
rect 4982 59218 5066 59454
rect 5302 59218 5334 59454
rect 4714 59134 5334 59218
rect 4714 58898 4746 59134
rect 4982 58898 5066 59134
rect 5302 58898 5334 59134
rect 4714 41454 5334 58898
rect 4714 41218 4746 41454
rect 4982 41218 5066 41454
rect 5302 41218 5334 41454
rect 4714 41134 5334 41218
rect 4714 40898 4746 41134
rect 4982 40898 5066 41134
rect 5302 40898 5334 41134
rect 4714 23454 5334 40898
rect 4714 23218 4746 23454
rect 4982 23218 5066 23454
rect 5302 23218 5334 23454
rect 4714 23134 5334 23218
rect 4714 22898 4746 23134
rect 4982 22898 5066 23134
rect 5302 22898 5334 23134
rect 4714 5454 5334 22898
rect 4714 5218 4746 5454
rect 4982 5218 5066 5454
rect 5302 5218 5334 5454
rect 4714 5134 5334 5218
rect 4714 4898 4746 5134
rect 4982 4898 5066 5134
rect 5302 4898 5334 5134
rect 4714 880 5334 4898
rect 8434 462052 9054 464004
rect 8434 461816 8466 462052
rect 8702 461816 8786 462052
rect 9022 461816 9054 462052
rect 8434 461732 9054 461816
rect 8434 461496 8466 461732
rect 8702 461496 8786 461732
rect 9022 461496 9054 461732
rect 8434 441174 9054 461496
rect 8434 440938 8466 441174
rect 8702 440938 8786 441174
rect 9022 440938 9054 441174
rect 8434 440854 9054 440938
rect 8434 440618 8466 440854
rect 8702 440618 8786 440854
rect 9022 440618 9054 440854
rect 8434 423174 9054 440618
rect 8434 422938 8466 423174
rect 8702 422938 8786 423174
rect 9022 422938 9054 423174
rect 8434 422854 9054 422938
rect 8434 422618 8466 422854
rect 8702 422618 8786 422854
rect 9022 422618 9054 422854
rect 8434 405174 9054 422618
rect 8434 404938 8466 405174
rect 8702 404938 8786 405174
rect 9022 404938 9054 405174
rect 8434 404854 9054 404938
rect 8434 404618 8466 404854
rect 8702 404618 8786 404854
rect 9022 404618 9054 404854
rect 8434 387174 9054 404618
rect 8434 386938 8466 387174
rect 8702 386938 8786 387174
rect 9022 386938 9054 387174
rect 8434 386854 9054 386938
rect 8434 386618 8466 386854
rect 8702 386618 8786 386854
rect 9022 386618 9054 386854
rect 8434 369174 9054 386618
rect 8434 368938 8466 369174
rect 8702 368938 8786 369174
rect 9022 368938 9054 369174
rect 8434 368854 9054 368938
rect 8434 368618 8466 368854
rect 8702 368618 8786 368854
rect 9022 368618 9054 368854
rect 8434 351174 9054 368618
rect 8434 350938 8466 351174
rect 8702 350938 8786 351174
rect 9022 350938 9054 351174
rect 8434 350854 9054 350938
rect 8434 350618 8466 350854
rect 8702 350618 8786 350854
rect 9022 350618 9054 350854
rect 8434 333174 9054 350618
rect 8434 332938 8466 333174
rect 8702 332938 8786 333174
rect 9022 332938 9054 333174
rect 8434 332854 9054 332938
rect 8434 332618 8466 332854
rect 8702 332618 8786 332854
rect 9022 332618 9054 332854
rect 8434 315174 9054 332618
rect 8434 314938 8466 315174
rect 8702 314938 8786 315174
rect 9022 314938 9054 315174
rect 8434 314854 9054 314938
rect 8434 314618 8466 314854
rect 8702 314618 8786 314854
rect 9022 314618 9054 314854
rect 8434 297174 9054 314618
rect 8434 296938 8466 297174
rect 8702 296938 8786 297174
rect 9022 296938 9054 297174
rect 8434 296854 9054 296938
rect 8434 296618 8466 296854
rect 8702 296618 8786 296854
rect 9022 296618 9054 296854
rect 8434 279174 9054 296618
rect 8434 278938 8466 279174
rect 8702 278938 8786 279174
rect 9022 278938 9054 279174
rect 8434 278854 9054 278938
rect 8434 278618 8466 278854
rect 8702 278618 8786 278854
rect 9022 278618 9054 278854
rect 8434 261174 9054 278618
rect 8434 260938 8466 261174
rect 8702 260938 8786 261174
rect 9022 260938 9054 261174
rect 8434 260854 9054 260938
rect 8434 260618 8466 260854
rect 8702 260618 8786 260854
rect 9022 260618 9054 260854
rect 8434 243174 9054 260618
rect 8434 242938 8466 243174
rect 8702 242938 8786 243174
rect 9022 242938 9054 243174
rect 8434 242854 9054 242938
rect 8434 242618 8466 242854
rect 8702 242618 8786 242854
rect 9022 242618 9054 242854
rect 8434 225174 9054 242618
rect 8434 224938 8466 225174
rect 8702 224938 8786 225174
rect 9022 224938 9054 225174
rect 8434 224854 9054 224938
rect 8434 224618 8466 224854
rect 8702 224618 8786 224854
rect 9022 224618 9054 224854
rect 8434 207174 9054 224618
rect 8434 206938 8466 207174
rect 8702 206938 8786 207174
rect 9022 206938 9054 207174
rect 8434 206854 9054 206938
rect 8434 206618 8466 206854
rect 8702 206618 8786 206854
rect 9022 206618 9054 206854
rect 8434 189174 9054 206618
rect 8434 188938 8466 189174
rect 8702 188938 8786 189174
rect 9022 188938 9054 189174
rect 8434 188854 9054 188938
rect 8434 188618 8466 188854
rect 8702 188618 8786 188854
rect 9022 188618 9054 188854
rect 8434 171174 9054 188618
rect 8434 170938 8466 171174
rect 8702 170938 8786 171174
rect 9022 170938 9054 171174
rect 8434 170854 9054 170938
rect 8434 170618 8466 170854
rect 8702 170618 8786 170854
rect 9022 170618 9054 170854
rect 8434 153174 9054 170618
rect 8434 152938 8466 153174
rect 8702 152938 8786 153174
rect 9022 152938 9054 153174
rect 8434 152854 9054 152938
rect 8434 152618 8466 152854
rect 8702 152618 8786 152854
rect 9022 152618 9054 152854
rect 8434 135174 9054 152618
rect 8434 134938 8466 135174
rect 8702 134938 8786 135174
rect 9022 134938 9054 135174
rect 8434 134854 9054 134938
rect 8434 134618 8466 134854
rect 8702 134618 8786 134854
rect 9022 134618 9054 134854
rect 8434 117174 9054 134618
rect 8434 116938 8466 117174
rect 8702 116938 8786 117174
rect 9022 116938 9054 117174
rect 8434 116854 9054 116938
rect 8434 116618 8466 116854
rect 8702 116618 8786 116854
rect 9022 116618 9054 116854
rect 8434 99174 9054 116618
rect 8434 98938 8466 99174
rect 8702 98938 8786 99174
rect 9022 98938 9054 99174
rect 8434 98854 9054 98938
rect 8434 98618 8466 98854
rect 8702 98618 8786 98854
rect 9022 98618 9054 98854
rect 8434 81174 9054 98618
rect 8434 80938 8466 81174
rect 8702 80938 8786 81174
rect 9022 80938 9054 81174
rect 8434 80854 9054 80938
rect 8434 80618 8466 80854
rect 8702 80618 8786 80854
rect 9022 80618 9054 80854
rect 8434 63174 9054 80618
rect 8434 62938 8466 63174
rect 8702 62938 8786 63174
rect 9022 62938 9054 63174
rect 8434 62854 9054 62938
rect 8434 62618 8466 62854
rect 8702 62618 8786 62854
rect 9022 62618 9054 62854
rect 8434 45174 9054 62618
rect 8434 44938 8466 45174
rect 8702 44938 8786 45174
rect 9022 44938 9054 45174
rect 8434 44854 9054 44938
rect 8434 44618 8466 44854
rect 8702 44618 8786 44854
rect 9022 44618 9054 44854
rect 8434 27174 9054 44618
rect 8434 26938 8466 27174
rect 8702 26938 8786 27174
rect 9022 26938 9054 27174
rect 8434 26854 9054 26938
rect 8434 26618 8466 26854
rect 8702 26618 8786 26854
rect 9022 26618 9054 26854
rect 8434 9174 9054 26618
rect 8434 8938 8466 9174
rect 8702 8938 8786 9174
rect 9022 8938 9054 9174
rect 8434 8854 9054 8938
rect 8434 8618 8466 8854
rect 8702 8618 8786 8854
rect 9022 8618 9054 8854
rect 8434 880 9054 8618
rect 12154 463012 12774 464004
rect 12154 462776 12186 463012
rect 12422 462776 12506 463012
rect 12742 462776 12774 463012
rect 12154 462692 12774 462776
rect 12154 462456 12186 462692
rect 12422 462456 12506 462692
rect 12742 462456 12774 462692
rect 12154 444894 12774 462456
rect 12154 444658 12186 444894
rect 12422 444658 12506 444894
rect 12742 444658 12774 444894
rect 12154 444574 12774 444658
rect 12154 444338 12186 444574
rect 12422 444338 12506 444574
rect 12742 444338 12774 444574
rect 12154 426894 12774 444338
rect 12154 426658 12186 426894
rect 12422 426658 12506 426894
rect 12742 426658 12774 426894
rect 12154 426574 12774 426658
rect 12154 426338 12186 426574
rect 12422 426338 12506 426574
rect 12742 426338 12774 426574
rect 12154 408894 12774 426338
rect 12154 408658 12186 408894
rect 12422 408658 12506 408894
rect 12742 408658 12774 408894
rect 12154 408574 12774 408658
rect 12154 408338 12186 408574
rect 12422 408338 12506 408574
rect 12742 408338 12774 408574
rect 12154 390894 12774 408338
rect 12154 390658 12186 390894
rect 12422 390658 12506 390894
rect 12742 390658 12774 390894
rect 12154 390574 12774 390658
rect 12154 390338 12186 390574
rect 12422 390338 12506 390574
rect 12742 390338 12774 390574
rect 12154 372894 12774 390338
rect 12154 372658 12186 372894
rect 12422 372658 12506 372894
rect 12742 372658 12774 372894
rect 12154 372574 12774 372658
rect 12154 372338 12186 372574
rect 12422 372338 12506 372574
rect 12742 372338 12774 372574
rect 12154 354894 12774 372338
rect 12154 354658 12186 354894
rect 12422 354658 12506 354894
rect 12742 354658 12774 354894
rect 12154 354574 12774 354658
rect 12154 354338 12186 354574
rect 12422 354338 12506 354574
rect 12742 354338 12774 354574
rect 12154 336894 12774 354338
rect 12154 336658 12186 336894
rect 12422 336658 12506 336894
rect 12742 336658 12774 336894
rect 12154 336574 12774 336658
rect 12154 336338 12186 336574
rect 12422 336338 12506 336574
rect 12742 336338 12774 336574
rect 12154 318894 12774 336338
rect 12154 318658 12186 318894
rect 12422 318658 12506 318894
rect 12742 318658 12774 318894
rect 12154 318574 12774 318658
rect 12154 318338 12186 318574
rect 12422 318338 12506 318574
rect 12742 318338 12774 318574
rect 12154 300894 12774 318338
rect 12154 300658 12186 300894
rect 12422 300658 12506 300894
rect 12742 300658 12774 300894
rect 12154 300574 12774 300658
rect 12154 300338 12186 300574
rect 12422 300338 12506 300574
rect 12742 300338 12774 300574
rect 12154 282894 12774 300338
rect 12154 282658 12186 282894
rect 12422 282658 12506 282894
rect 12742 282658 12774 282894
rect 12154 282574 12774 282658
rect 12154 282338 12186 282574
rect 12422 282338 12506 282574
rect 12742 282338 12774 282574
rect 12154 264894 12774 282338
rect 12154 264658 12186 264894
rect 12422 264658 12506 264894
rect 12742 264658 12774 264894
rect 12154 264574 12774 264658
rect 12154 264338 12186 264574
rect 12422 264338 12506 264574
rect 12742 264338 12774 264574
rect 12154 246894 12774 264338
rect 12154 246658 12186 246894
rect 12422 246658 12506 246894
rect 12742 246658 12774 246894
rect 12154 246574 12774 246658
rect 12154 246338 12186 246574
rect 12422 246338 12506 246574
rect 12742 246338 12774 246574
rect 12154 228894 12774 246338
rect 12154 228658 12186 228894
rect 12422 228658 12506 228894
rect 12742 228658 12774 228894
rect 12154 228574 12774 228658
rect 12154 228338 12186 228574
rect 12422 228338 12506 228574
rect 12742 228338 12774 228574
rect 12154 210894 12774 228338
rect 12154 210658 12186 210894
rect 12422 210658 12506 210894
rect 12742 210658 12774 210894
rect 12154 210574 12774 210658
rect 12154 210338 12186 210574
rect 12422 210338 12506 210574
rect 12742 210338 12774 210574
rect 12154 192894 12774 210338
rect 12154 192658 12186 192894
rect 12422 192658 12506 192894
rect 12742 192658 12774 192894
rect 12154 192574 12774 192658
rect 12154 192338 12186 192574
rect 12422 192338 12506 192574
rect 12742 192338 12774 192574
rect 12154 174894 12774 192338
rect 12154 174658 12186 174894
rect 12422 174658 12506 174894
rect 12742 174658 12774 174894
rect 12154 174574 12774 174658
rect 12154 174338 12186 174574
rect 12422 174338 12506 174574
rect 12742 174338 12774 174574
rect 12154 156894 12774 174338
rect 12154 156658 12186 156894
rect 12422 156658 12506 156894
rect 12742 156658 12774 156894
rect 12154 156574 12774 156658
rect 12154 156338 12186 156574
rect 12422 156338 12506 156574
rect 12742 156338 12774 156574
rect 12154 138894 12774 156338
rect 12154 138658 12186 138894
rect 12422 138658 12506 138894
rect 12742 138658 12774 138894
rect 12154 138574 12774 138658
rect 12154 138338 12186 138574
rect 12422 138338 12506 138574
rect 12742 138338 12774 138574
rect 12154 120894 12774 138338
rect 12154 120658 12186 120894
rect 12422 120658 12506 120894
rect 12742 120658 12774 120894
rect 12154 120574 12774 120658
rect 12154 120338 12186 120574
rect 12422 120338 12506 120574
rect 12742 120338 12774 120574
rect 12154 102894 12774 120338
rect 12154 102658 12186 102894
rect 12422 102658 12506 102894
rect 12742 102658 12774 102894
rect 12154 102574 12774 102658
rect 12154 102338 12186 102574
rect 12422 102338 12506 102574
rect 12742 102338 12774 102574
rect 12154 84894 12774 102338
rect 12154 84658 12186 84894
rect 12422 84658 12506 84894
rect 12742 84658 12774 84894
rect 12154 84574 12774 84658
rect 12154 84338 12186 84574
rect 12422 84338 12506 84574
rect 12742 84338 12774 84574
rect 12154 66894 12774 84338
rect 12154 66658 12186 66894
rect 12422 66658 12506 66894
rect 12742 66658 12774 66894
rect 12154 66574 12774 66658
rect 12154 66338 12186 66574
rect 12422 66338 12506 66574
rect 12742 66338 12774 66574
rect 12154 48894 12774 66338
rect 12154 48658 12186 48894
rect 12422 48658 12506 48894
rect 12742 48658 12774 48894
rect 12154 48574 12774 48658
rect 12154 48338 12186 48574
rect 12422 48338 12506 48574
rect 12742 48338 12774 48574
rect 12154 30894 12774 48338
rect 12154 30658 12186 30894
rect 12422 30658 12506 30894
rect 12742 30658 12774 30894
rect 12154 30574 12774 30658
rect 12154 30338 12186 30574
rect 12422 30338 12506 30574
rect 12742 30338 12774 30574
rect 12154 12894 12774 30338
rect 12154 12658 12186 12894
rect 12422 12658 12506 12894
rect 12742 12658 12774 12894
rect 12154 12574 12774 12658
rect 12154 12338 12186 12574
rect 12422 12338 12506 12574
rect 12742 12338 12774 12574
rect 12154 880 12774 12338
rect 15874 463972 16494 464004
rect 15874 463736 15906 463972
rect 16142 463736 16226 463972
rect 16462 463736 16494 463972
rect 15874 463652 16494 463736
rect 15874 463416 15906 463652
rect 16142 463416 16226 463652
rect 16462 463416 16494 463652
rect 15874 448614 16494 463416
rect 15874 448378 15906 448614
rect 16142 448378 16226 448614
rect 16462 448378 16494 448614
rect 15874 448294 16494 448378
rect 15874 448058 15906 448294
rect 16142 448058 16226 448294
rect 16462 448058 16494 448294
rect 15874 430614 16494 448058
rect 15874 430378 15906 430614
rect 16142 430378 16226 430614
rect 16462 430378 16494 430614
rect 15874 430294 16494 430378
rect 15874 430058 15906 430294
rect 16142 430058 16226 430294
rect 16462 430058 16494 430294
rect 15874 412614 16494 430058
rect 15874 412378 15906 412614
rect 16142 412378 16226 412614
rect 16462 412378 16494 412614
rect 15874 412294 16494 412378
rect 15874 412058 15906 412294
rect 16142 412058 16226 412294
rect 16462 412058 16494 412294
rect 15874 394614 16494 412058
rect 15874 394378 15906 394614
rect 16142 394378 16226 394614
rect 16462 394378 16494 394614
rect 15874 394294 16494 394378
rect 15874 394058 15906 394294
rect 16142 394058 16226 394294
rect 16462 394058 16494 394294
rect 15874 376614 16494 394058
rect 15874 376378 15906 376614
rect 16142 376378 16226 376614
rect 16462 376378 16494 376614
rect 15874 376294 16494 376378
rect 15874 376058 15906 376294
rect 16142 376058 16226 376294
rect 16462 376058 16494 376294
rect 15874 358614 16494 376058
rect 15874 358378 15906 358614
rect 16142 358378 16226 358614
rect 16462 358378 16494 358614
rect 15874 358294 16494 358378
rect 15874 358058 15906 358294
rect 16142 358058 16226 358294
rect 16462 358058 16494 358294
rect 15874 340614 16494 358058
rect 15874 340378 15906 340614
rect 16142 340378 16226 340614
rect 16462 340378 16494 340614
rect 15874 340294 16494 340378
rect 15874 340058 15906 340294
rect 16142 340058 16226 340294
rect 16462 340058 16494 340294
rect 15874 322614 16494 340058
rect 15874 322378 15906 322614
rect 16142 322378 16226 322614
rect 16462 322378 16494 322614
rect 15874 322294 16494 322378
rect 15874 322058 15906 322294
rect 16142 322058 16226 322294
rect 16462 322058 16494 322294
rect 15874 304614 16494 322058
rect 15874 304378 15906 304614
rect 16142 304378 16226 304614
rect 16462 304378 16494 304614
rect 15874 304294 16494 304378
rect 15874 304058 15906 304294
rect 16142 304058 16226 304294
rect 16462 304058 16494 304294
rect 15874 286614 16494 304058
rect 15874 286378 15906 286614
rect 16142 286378 16226 286614
rect 16462 286378 16494 286614
rect 15874 286294 16494 286378
rect 15874 286058 15906 286294
rect 16142 286058 16226 286294
rect 16462 286058 16494 286294
rect 15874 268614 16494 286058
rect 15874 268378 15906 268614
rect 16142 268378 16226 268614
rect 16462 268378 16494 268614
rect 15874 268294 16494 268378
rect 15874 268058 15906 268294
rect 16142 268058 16226 268294
rect 16462 268058 16494 268294
rect 15874 250614 16494 268058
rect 15874 250378 15906 250614
rect 16142 250378 16226 250614
rect 16462 250378 16494 250614
rect 15874 250294 16494 250378
rect 15874 250058 15906 250294
rect 16142 250058 16226 250294
rect 16462 250058 16494 250294
rect 15874 232614 16494 250058
rect 15874 232378 15906 232614
rect 16142 232378 16226 232614
rect 16462 232378 16494 232614
rect 15874 232294 16494 232378
rect 15874 232058 15906 232294
rect 16142 232058 16226 232294
rect 16462 232058 16494 232294
rect 15874 214614 16494 232058
rect 15874 214378 15906 214614
rect 16142 214378 16226 214614
rect 16462 214378 16494 214614
rect 15874 214294 16494 214378
rect 15874 214058 15906 214294
rect 16142 214058 16226 214294
rect 16462 214058 16494 214294
rect 15874 196614 16494 214058
rect 15874 196378 15906 196614
rect 16142 196378 16226 196614
rect 16462 196378 16494 196614
rect 15874 196294 16494 196378
rect 15874 196058 15906 196294
rect 16142 196058 16226 196294
rect 16462 196058 16494 196294
rect 15874 178614 16494 196058
rect 15874 178378 15906 178614
rect 16142 178378 16226 178614
rect 16462 178378 16494 178614
rect 15874 178294 16494 178378
rect 15874 178058 15906 178294
rect 16142 178058 16226 178294
rect 16462 178058 16494 178294
rect 15874 160614 16494 178058
rect 15874 160378 15906 160614
rect 16142 160378 16226 160614
rect 16462 160378 16494 160614
rect 15874 160294 16494 160378
rect 15874 160058 15906 160294
rect 16142 160058 16226 160294
rect 16462 160058 16494 160294
rect 15874 142614 16494 160058
rect 15874 142378 15906 142614
rect 16142 142378 16226 142614
rect 16462 142378 16494 142614
rect 15874 142294 16494 142378
rect 15874 142058 15906 142294
rect 16142 142058 16226 142294
rect 16462 142058 16494 142294
rect 15874 124614 16494 142058
rect 15874 124378 15906 124614
rect 16142 124378 16226 124614
rect 16462 124378 16494 124614
rect 15874 124294 16494 124378
rect 15874 124058 15906 124294
rect 16142 124058 16226 124294
rect 16462 124058 16494 124294
rect 15874 106614 16494 124058
rect 15874 106378 15906 106614
rect 16142 106378 16226 106614
rect 16462 106378 16494 106614
rect 15874 106294 16494 106378
rect 15874 106058 15906 106294
rect 16142 106058 16226 106294
rect 16462 106058 16494 106294
rect 15874 88614 16494 106058
rect 15874 88378 15906 88614
rect 16142 88378 16226 88614
rect 16462 88378 16494 88614
rect 15874 88294 16494 88378
rect 15874 88058 15906 88294
rect 16142 88058 16226 88294
rect 16462 88058 16494 88294
rect 15874 70614 16494 88058
rect 15874 70378 15906 70614
rect 16142 70378 16226 70614
rect 16462 70378 16494 70614
rect 15874 70294 16494 70378
rect 15874 70058 15906 70294
rect 16142 70058 16226 70294
rect 16462 70058 16494 70294
rect 15874 52614 16494 70058
rect 15874 52378 15906 52614
rect 16142 52378 16226 52614
rect 16462 52378 16494 52614
rect 15874 52294 16494 52378
rect 15874 52058 15906 52294
rect 16142 52058 16226 52294
rect 16462 52058 16494 52294
rect 15874 34614 16494 52058
rect 15874 34378 15906 34614
rect 16142 34378 16226 34614
rect 16462 34378 16494 34614
rect 15874 34294 16494 34378
rect 15874 34058 15906 34294
rect 16142 34058 16226 34294
rect 16462 34058 16494 34294
rect 15874 16614 16494 34058
rect 15874 16378 15906 16614
rect 16142 16378 16226 16614
rect 16462 16378 16494 16614
rect 15874 16294 16494 16378
rect 15874 16058 15906 16294
rect 16142 16058 16226 16294
rect 16462 16058 16494 16294
rect 15874 880 16494 16058
rect 22714 461092 23334 464004
rect 22714 460856 22746 461092
rect 22982 460856 23066 461092
rect 23302 460856 23334 461092
rect 22714 460772 23334 460856
rect 22714 460536 22746 460772
rect 22982 460536 23066 460772
rect 23302 460536 23334 460772
rect 22714 455454 23334 460536
rect 22714 455218 22746 455454
rect 22982 455218 23066 455454
rect 23302 455218 23334 455454
rect 22714 455134 23334 455218
rect 22714 454898 22746 455134
rect 22982 454898 23066 455134
rect 23302 454898 23334 455134
rect 22714 437454 23334 454898
rect 22714 437218 22746 437454
rect 22982 437218 23066 437454
rect 23302 437218 23334 437454
rect 22714 437134 23334 437218
rect 22714 436898 22746 437134
rect 22982 436898 23066 437134
rect 23302 436898 23334 437134
rect 22714 419454 23334 436898
rect 22714 419218 22746 419454
rect 22982 419218 23066 419454
rect 23302 419218 23334 419454
rect 22714 419134 23334 419218
rect 22714 418898 22746 419134
rect 22982 418898 23066 419134
rect 23302 418898 23334 419134
rect 22714 401454 23334 418898
rect 22714 401218 22746 401454
rect 22982 401218 23066 401454
rect 23302 401218 23334 401454
rect 22714 401134 23334 401218
rect 22714 400898 22746 401134
rect 22982 400898 23066 401134
rect 23302 400898 23334 401134
rect 22714 383454 23334 400898
rect 22714 383218 22746 383454
rect 22982 383218 23066 383454
rect 23302 383218 23334 383454
rect 22714 383134 23334 383218
rect 22714 382898 22746 383134
rect 22982 382898 23066 383134
rect 23302 382898 23334 383134
rect 22714 365454 23334 382898
rect 22714 365218 22746 365454
rect 22982 365218 23066 365454
rect 23302 365218 23334 365454
rect 22714 365134 23334 365218
rect 22714 364898 22746 365134
rect 22982 364898 23066 365134
rect 23302 364898 23334 365134
rect 22714 347454 23334 364898
rect 22714 347218 22746 347454
rect 22982 347218 23066 347454
rect 23302 347218 23334 347454
rect 22714 347134 23334 347218
rect 22714 346898 22746 347134
rect 22982 346898 23066 347134
rect 23302 346898 23334 347134
rect 22714 329454 23334 346898
rect 22714 329218 22746 329454
rect 22982 329218 23066 329454
rect 23302 329218 23334 329454
rect 22714 329134 23334 329218
rect 22714 328898 22746 329134
rect 22982 328898 23066 329134
rect 23302 328898 23334 329134
rect 22714 311454 23334 328898
rect 22714 311218 22746 311454
rect 22982 311218 23066 311454
rect 23302 311218 23334 311454
rect 22714 311134 23334 311218
rect 22714 310898 22746 311134
rect 22982 310898 23066 311134
rect 23302 310898 23334 311134
rect 22714 293454 23334 310898
rect 22714 293218 22746 293454
rect 22982 293218 23066 293454
rect 23302 293218 23334 293454
rect 22714 293134 23334 293218
rect 22714 292898 22746 293134
rect 22982 292898 23066 293134
rect 23302 292898 23334 293134
rect 22714 275454 23334 292898
rect 22714 275218 22746 275454
rect 22982 275218 23066 275454
rect 23302 275218 23334 275454
rect 22714 275134 23334 275218
rect 22714 274898 22746 275134
rect 22982 274898 23066 275134
rect 23302 274898 23334 275134
rect 22714 257454 23334 274898
rect 22714 257218 22746 257454
rect 22982 257218 23066 257454
rect 23302 257218 23334 257454
rect 22714 257134 23334 257218
rect 22714 256898 22746 257134
rect 22982 256898 23066 257134
rect 23302 256898 23334 257134
rect 22714 239454 23334 256898
rect 22714 239218 22746 239454
rect 22982 239218 23066 239454
rect 23302 239218 23334 239454
rect 22714 239134 23334 239218
rect 22714 238898 22746 239134
rect 22982 238898 23066 239134
rect 23302 238898 23334 239134
rect 22714 221454 23334 238898
rect 22714 221218 22746 221454
rect 22982 221218 23066 221454
rect 23302 221218 23334 221454
rect 22714 221134 23334 221218
rect 22714 220898 22746 221134
rect 22982 220898 23066 221134
rect 23302 220898 23334 221134
rect 22714 203454 23334 220898
rect 22714 203218 22746 203454
rect 22982 203218 23066 203454
rect 23302 203218 23334 203454
rect 22714 203134 23334 203218
rect 22714 202898 22746 203134
rect 22982 202898 23066 203134
rect 23302 202898 23334 203134
rect 22714 185454 23334 202898
rect 22714 185218 22746 185454
rect 22982 185218 23066 185454
rect 23302 185218 23334 185454
rect 22714 185134 23334 185218
rect 22714 184898 22746 185134
rect 22982 184898 23066 185134
rect 23302 184898 23334 185134
rect 22714 167454 23334 184898
rect 22714 167218 22746 167454
rect 22982 167218 23066 167454
rect 23302 167218 23334 167454
rect 22714 167134 23334 167218
rect 22714 166898 22746 167134
rect 22982 166898 23066 167134
rect 23302 166898 23334 167134
rect 22714 149454 23334 166898
rect 22714 149218 22746 149454
rect 22982 149218 23066 149454
rect 23302 149218 23334 149454
rect 22714 149134 23334 149218
rect 22714 148898 22746 149134
rect 22982 148898 23066 149134
rect 23302 148898 23334 149134
rect 22714 131454 23334 148898
rect 22714 131218 22746 131454
rect 22982 131218 23066 131454
rect 23302 131218 23334 131454
rect 22714 131134 23334 131218
rect 22714 130898 22746 131134
rect 22982 130898 23066 131134
rect 23302 130898 23334 131134
rect 22714 113454 23334 130898
rect 22714 113218 22746 113454
rect 22982 113218 23066 113454
rect 23302 113218 23334 113454
rect 22714 113134 23334 113218
rect 22714 112898 22746 113134
rect 22982 112898 23066 113134
rect 23302 112898 23334 113134
rect 22714 95454 23334 112898
rect 22714 95218 22746 95454
rect 22982 95218 23066 95454
rect 23302 95218 23334 95454
rect 22714 95134 23334 95218
rect 22714 94898 22746 95134
rect 22982 94898 23066 95134
rect 23302 94898 23334 95134
rect 22714 77454 23334 94898
rect 22714 77218 22746 77454
rect 22982 77218 23066 77454
rect 23302 77218 23334 77454
rect 22714 77134 23334 77218
rect 22714 76898 22746 77134
rect 22982 76898 23066 77134
rect 23302 76898 23334 77134
rect 22714 59454 23334 76898
rect 22714 59218 22746 59454
rect 22982 59218 23066 59454
rect 23302 59218 23334 59454
rect 22714 59134 23334 59218
rect 22714 58898 22746 59134
rect 22982 58898 23066 59134
rect 23302 58898 23334 59134
rect 22714 41454 23334 58898
rect 22714 41218 22746 41454
rect 22982 41218 23066 41454
rect 23302 41218 23334 41454
rect 22714 41134 23334 41218
rect 22714 40898 22746 41134
rect 22982 40898 23066 41134
rect 23302 40898 23334 41134
rect 22714 23454 23334 40898
rect 22714 23218 22746 23454
rect 22982 23218 23066 23454
rect 23302 23218 23334 23454
rect 22714 23134 23334 23218
rect 22714 22898 22746 23134
rect 22982 22898 23066 23134
rect 23302 22898 23334 23134
rect 22714 5454 23334 22898
rect 22714 5218 22746 5454
rect 22982 5218 23066 5454
rect 23302 5218 23334 5454
rect 22714 5134 23334 5218
rect 22714 4898 22746 5134
rect 22982 4898 23066 5134
rect 23302 4898 23334 5134
rect 22714 880 23334 4898
rect 26434 462052 27054 464004
rect 26434 461816 26466 462052
rect 26702 461816 26786 462052
rect 27022 461816 27054 462052
rect 26434 461732 27054 461816
rect 26434 461496 26466 461732
rect 26702 461496 26786 461732
rect 27022 461496 27054 461732
rect 26434 441174 27054 461496
rect 26434 440938 26466 441174
rect 26702 440938 26786 441174
rect 27022 440938 27054 441174
rect 26434 440854 27054 440938
rect 26434 440618 26466 440854
rect 26702 440618 26786 440854
rect 27022 440618 27054 440854
rect 26434 423174 27054 440618
rect 26434 422938 26466 423174
rect 26702 422938 26786 423174
rect 27022 422938 27054 423174
rect 26434 422854 27054 422938
rect 26434 422618 26466 422854
rect 26702 422618 26786 422854
rect 27022 422618 27054 422854
rect 26434 405174 27054 422618
rect 26434 404938 26466 405174
rect 26702 404938 26786 405174
rect 27022 404938 27054 405174
rect 26434 404854 27054 404938
rect 26434 404618 26466 404854
rect 26702 404618 26786 404854
rect 27022 404618 27054 404854
rect 26434 387174 27054 404618
rect 26434 386938 26466 387174
rect 26702 386938 26786 387174
rect 27022 386938 27054 387174
rect 26434 386854 27054 386938
rect 26434 386618 26466 386854
rect 26702 386618 26786 386854
rect 27022 386618 27054 386854
rect 26434 369174 27054 386618
rect 26434 368938 26466 369174
rect 26702 368938 26786 369174
rect 27022 368938 27054 369174
rect 26434 368854 27054 368938
rect 26434 368618 26466 368854
rect 26702 368618 26786 368854
rect 27022 368618 27054 368854
rect 26434 351174 27054 368618
rect 26434 350938 26466 351174
rect 26702 350938 26786 351174
rect 27022 350938 27054 351174
rect 26434 350854 27054 350938
rect 26434 350618 26466 350854
rect 26702 350618 26786 350854
rect 27022 350618 27054 350854
rect 26434 333174 27054 350618
rect 26434 332938 26466 333174
rect 26702 332938 26786 333174
rect 27022 332938 27054 333174
rect 26434 332854 27054 332938
rect 26434 332618 26466 332854
rect 26702 332618 26786 332854
rect 27022 332618 27054 332854
rect 26434 315174 27054 332618
rect 26434 314938 26466 315174
rect 26702 314938 26786 315174
rect 27022 314938 27054 315174
rect 26434 314854 27054 314938
rect 26434 314618 26466 314854
rect 26702 314618 26786 314854
rect 27022 314618 27054 314854
rect 26434 297174 27054 314618
rect 26434 296938 26466 297174
rect 26702 296938 26786 297174
rect 27022 296938 27054 297174
rect 26434 296854 27054 296938
rect 26434 296618 26466 296854
rect 26702 296618 26786 296854
rect 27022 296618 27054 296854
rect 26434 279174 27054 296618
rect 26434 278938 26466 279174
rect 26702 278938 26786 279174
rect 27022 278938 27054 279174
rect 26434 278854 27054 278938
rect 26434 278618 26466 278854
rect 26702 278618 26786 278854
rect 27022 278618 27054 278854
rect 26434 261174 27054 278618
rect 26434 260938 26466 261174
rect 26702 260938 26786 261174
rect 27022 260938 27054 261174
rect 26434 260854 27054 260938
rect 26434 260618 26466 260854
rect 26702 260618 26786 260854
rect 27022 260618 27054 260854
rect 26434 243174 27054 260618
rect 26434 242938 26466 243174
rect 26702 242938 26786 243174
rect 27022 242938 27054 243174
rect 26434 242854 27054 242938
rect 26434 242618 26466 242854
rect 26702 242618 26786 242854
rect 27022 242618 27054 242854
rect 26434 225174 27054 242618
rect 26434 224938 26466 225174
rect 26702 224938 26786 225174
rect 27022 224938 27054 225174
rect 26434 224854 27054 224938
rect 26434 224618 26466 224854
rect 26702 224618 26786 224854
rect 27022 224618 27054 224854
rect 26434 207174 27054 224618
rect 26434 206938 26466 207174
rect 26702 206938 26786 207174
rect 27022 206938 27054 207174
rect 26434 206854 27054 206938
rect 26434 206618 26466 206854
rect 26702 206618 26786 206854
rect 27022 206618 27054 206854
rect 26434 189174 27054 206618
rect 26434 188938 26466 189174
rect 26702 188938 26786 189174
rect 27022 188938 27054 189174
rect 26434 188854 27054 188938
rect 26434 188618 26466 188854
rect 26702 188618 26786 188854
rect 27022 188618 27054 188854
rect 26434 171174 27054 188618
rect 26434 170938 26466 171174
rect 26702 170938 26786 171174
rect 27022 170938 27054 171174
rect 26434 170854 27054 170938
rect 26434 170618 26466 170854
rect 26702 170618 26786 170854
rect 27022 170618 27054 170854
rect 26434 153174 27054 170618
rect 26434 152938 26466 153174
rect 26702 152938 26786 153174
rect 27022 152938 27054 153174
rect 26434 152854 27054 152938
rect 26434 152618 26466 152854
rect 26702 152618 26786 152854
rect 27022 152618 27054 152854
rect 26434 135174 27054 152618
rect 26434 134938 26466 135174
rect 26702 134938 26786 135174
rect 27022 134938 27054 135174
rect 26434 134854 27054 134938
rect 26434 134618 26466 134854
rect 26702 134618 26786 134854
rect 27022 134618 27054 134854
rect 26434 117174 27054 134618
rect 26434 116938 26466 117174
rect 26702 116938 26786 117174
rect 27022 116938 27054 117174
rect 26434 116854 27054 116938
rect 26434 116618 26466 116854
rect 26702 116618 26786 116854
rect 27022 116618 27054 116854
rect 26434 99174 27054 116618
rect 26434 98938 26466 99174
rect 26702 98938 26786 99174
rect 27022 98938 27054 99174
rect 26434 98854 27054 98938
rect 26434 98618 26466 98854
rect 26702 98618 26786 98854
rect 27022 98618 27054 98854
rect 26434 81174 27054 98618
rect 26434 80938 26466 81174
rect 26702 80938 26786 81174
rect 27022 80938 27054 81174
rect 26434 80854 27054 80938
rect 26434 80618 26466 80854
rect 26702 80618 26786 80854
rect 27022 80618 27054 80854
rect 26434 63174 27054 80618
rect 26434 62938 26466 63174
rect 26702 62938 26786 63174
rect 27022 62938 27054 63174
rect 26434 62854 27054 62938
rect 26434 62618 26466 62854
rect 26702 62618 26786 62854
rect 27022 62618 27054 62854
rect 26434 45174 27054 62618
rect 26434 44938 26466 45174
rect 26702 44938 26786 45174
rect 27022 44938 27054 45174
rect 26434 44854 27054 44938
rect 26434 44618 26466 44854
rect 26702 44618 26786 44854
rect 27022 44618 27054 44854
rect 26434 27174 27054 44618
rect 26434 26938 26466 27174
rect 26702 26938 26786 27174
rect 27022 26938 27054 27174
rect 26434 26854 27054 26938
rect 26434 26618 26466 26854
rect 26702 26618 26786 26854
rect 27022 26618 27054 26854
rect 26434 9174 27054 26618
rect 26434 8938 26466 9174
rect 26702 8938 26786 9174
rect 27022 8938 27054 9174
rect 26434 8854 27054 8938
rect 26434 8618 26466 8854
rect 26702 8618 26786 8854
rect 27022 8618 27054 8854
rect 26434 880 27054 8618
rect 30154 463012 30774 464004
rect 30154 462776 30186 463012
rect 30422 462776 30506 463012
rect 30742 462776 30774 463012
rect 30154 462692 30774 462776
rect 30154 462456 30186 462692
rect 30422 462456 30506 462692
rect 30742 462456 30774 462692
rect 30154 444894 30774 462456
rect 30154 444658 30186 444894
rect 30422 444658 30506 444894
rect 30742 444658 30774 444894
rect 30154 444574 30774 444658
rect 30154 444338 30186 444574
rect 30422 444338 30506 444574
rect 30742 444338 30774 444574
rect 30154 426894 30774 444338
rect 30154 426658 30186 426894
rect 30422 426658 30506 426894
rect 30742 426658 30774 426894
rect 30154 426574 30774 426658
rect 30154 426338 30186 426574
rect 30422 426338 30506 426574
rect 30742 426338 30774 426574
rect 30154 408894 30774 426338
rect 30154 408658 30186 408894
rect 30422 408658 30506 408894
rect 30742 408658 30774 408894
rect 30154 408574 30774 408658
rect 30154 408338 30186 408574
rect 30422 408338 30506 408574
rect 30742 408338 30774 408574
rect 30154 390894 30774 408338
rect 30154 390658 30186 390894
rect 30422 390658 30506 390894
rect 30742 390658 30774 390894
rect 30154 390574 30774 390658
rect 30154 390338 30186 390574
rect 30422 390338 30506 390574
rect 30742 390338 30774 390574
rect 30154 372894 30774 390338
rect 30154 372658 30186 372894
rect 30422 372658 30506 372894
rect 30742 372658 30774 372894
rect 30154 372574 30774 372658
rect 30154 372338 30186 372574
rect 30422 372338 30506 372574
rect 30742 372338 30774 372574
rect 30154 354894 30774 372338
rect 30154 354658 30186 354894
rect 30422 354658 30506 354894
rect 30742 354658 30774 354894
rect 30154 354574 30774 354658
rect 30154 354338 30186 354574
rect 30422 354338 30506 354574
rect 30742 354338 30774 354574
rect 30154 336894 30774 354338
rect 30154 336658 30186 336894
rect 30422 336658 30506 336894
rect 30742 336658 30774 336894
rect 30154 336574 30774 336658
rect 30154 336338 30186 336574
rect 30422 336338 30506 336574
rect 30742 336338 30774 336574
rect 30154 318894 30774 336338
rect 30154 318658 30186 318894
rect 30422 318658 30506 318894
rect 30742 318658 30774 318894
rect 30154 318574 30774 318658
rect 30154 318338 30186 318574
rect 30422 318338 30506 318574
rect 30742 318338 30774 318574
rect 30154 300894 30774 318338
rect 30154 300658 30186 300894
rect 30422 300658 30506 300894
rect 30742 300658 30774 300894
rect 30154 300574 30774 300658
rect 30154 300338 30186 300574
rect 30422 300338 30506 300574
rect 30742 300338 30774 300574
rect 30154 282894 30774 300338
rect 30154 282658 30186 282894
rect 30422 282658 30506 282894
rect 30742 282658 30774 282894
rect 30154 282574 30774 282658
rect 30154 282338 30186 282574
rect 30422 282338 30506 282574
rect 30742 282338 30774 282574
rect 30154 264894 30774 282338
rect 30154 264658 30186 264894
rect 30422 264658 30506 264894
rect 30742 264658 30774 264894
rect 30154 264574 30774 264658
rect 30154 264338 30186 264574
rect 30422 264338 30506 264574
rect 30742 264338 30774 264574
rect 30154 246894 30774 264338
rect 30154 246658 30186 246894
rect 30422 246658 30506 246894
rect 30742 246658 30774 246894
rect 30154 246574 30774 246658
rect 30154 246338 30186 246574
rect 30422 246338 30506 246574
rect 30742 246338 30774 246574
rect 30154 228894 30774 246338
rect 30154 228658 30186 228894
rect 30422 228658 30506 228894
rect 30742 228658 30774 228894
rect 30154 228574 30774 228658
rect 30154 228338 30186 228574
rect 30422 228338 30506 228574
rect 30742 228338 30774 228574
rect 30154 210894 30774 228338
rect 30154 210658 30186 210894
rect 30422 210658 30506 210894
rect 30742 210658 30774 210894
rect 30154 210574 30774 210658
rect 30154 210338 30186 210574
rect 30422 210338 30506 210574
rect 30742 210338 30774 210574
rect 30154 192894 30774 210338
rect 30154 192658 30186 192894
rect 30422 192658 30506 192894
rect 30742 192658 30774 192894
rect 30154 192574 30774 192658
rect 30154 192338 30186 192574
rect 30422 192338 30506 192574
rect 30742 192338 30774 192574
rect 30154 174894 30774 192338
rect 30154 174658 30186 174894
rect 30422 174658 30506 174894
rect 30742 174658 30774 174894
rect 30154 174574 30774 174658
rect 30154 174338 30186 174574
rect 30422 174338 30506 174574
rect 30742 174338 30774 174574
rect 30154 156894 30774 174338
rect 30154 156658 30186 156894
rect 30422 156658 30506 156894
rect 30742 156658 30774 156894
rect 30154 156574 30774 156658
rect 30154 156338 30186 156574
rect 30422 156338 30506 156574
rect 30742 156338 30774 156574
rect 30154 138894 30774 156338
rect 30154 138658 30186 138894
rect 30422 138658 30506 138894
rect 30742 138658 30774 138894
rect 30154 138574 30774 138658
rect 30154 138338 30186 138574
rect 30422 138338 30506 138574
rect 30742 138338 30774 138574
rect 30154 120894 30774 138338
rect 30154 120658 30186 120894
rect 30422 120658 30506 120894
rect 30742 120658 30774 120894
rect 30154 120574 30774 120658
rect 30154 120338 30186 120574
rect 30422 120338 30506 120574
rect 30742 120338 30774 120574
rect 30154 102894 30774 120338
rect 30154 102658 30186 102894
rect 30422 102658 30506 102894
rect 30742 102658 30774 102894
rect 30154 102574 30774 102658
rect 30154 102338 30186 102574
rect 30422 102338 30506 102574
rect 30742 102338 30774 102574
rect 30154 84894 30774 102338
rect 30154 84658 30186 84894
rect 30422 84658 30506 84894
rect 30742 84658 30774 84894
rect 30154 84574 30774 84658
rect 30154 84338 30186 84574
rect 30422 84338 30506 84574
rect 30742 84338 30774 84574
rect 30154 66894 30774 84338
rect 30154 66658 30186 66894
rect 30422 66658 30506 66894
rect 30742 66658 30774 66894
rect 30154 66574 30774 66658
rect 30154 66338 30186 66574
rect 30422 66338 30506 66574
rect 30742 66338 30774 66574
rect 30154 48894 30774 66338
rect 30154 48658 30186 48894
rect 30422 48658 30506 48894
rect 30742 48658 30774 48894
rect 30154 48574 30774 48658
rect 30154 48338 30186 48574
rect 30422 48338 30506 48574
rect 30742 48338 30774 48574
rect 30154 30894 30774 48338
rect 30154 30658 30186 30894
rect 30422 30658 30506 30894
rect 30742 30658 30774 30894
rect 30154 30574 30774 30658
rect 30154 30338 30186 30574
rect 30422 30338 30506 30574
rect 30742 30338 30774 30574
rect 30154 12894 30774 30338
rect 30154 12658 30186 12894
rect 30422 12658 30506 12894
rect 30742 12658 30774 12894
rect 30154 12574 30774 12658
rect 30154 12338 30186 12574
rect 30422 12338 30506 12574
rect 30742 12338 30774 12574
rect 30154 880 30774 12338
rect 33874 463972 34494 464004
rect 33874 463736 33906 463972
rect 34142 463736 34226 463972
rect 34462 463736 34494 463972
rect 33874 463652 34494 463736
rect 33874 463416 33906 463652
rect 34142 463416 34226 463652
rect 34462 463416 34494 463652
rect 33874 448614 34494 463416
rect 33874 448378 33906 448614
rect 34142 448378 34226 448614
rect 34462 448378 34494 448614
rect 33874 448294 34494 448378
rect 33874 448058 33906 448294
rect 34142 448058 34226 448294
rect 34462 448058 34494 448294
rect 33874 430614 34494 448058
rect 33874 430378 33906 430614
rect 34142 430378 34226 430614
rect 34462 430378 34494 430614
rect 33874 430294 34494 430378
rect 33874 430058 33906 430294
rect 34142 430058 34226 430294
rect 34462 430058 34494 430294
rect 33874 412614 34494 430058
rect 33874 412378 33906 412614
rect 34142 412378 34226 412614
rect 34462 412378 34494 412614
rect 33874 412294 34494 412378
rect 33874 412058 33906 412294
rect 34142 412058 34226 412294
rect 34462 412058 34494 412294
rect 33874 394614 34494 412058
rect 33874 394378 33906 394614
rect 34142 394378 34226 394614
rect 34462 394378 34494 394614
rect 33874 394294 34494 394378
rect 33874 394058 33906 394294
rect 34142 394058 34226 394294
rect 34462 394058 34494 394294
rect 33874 376614 34494 394058
rect 33874 376378 33906 376614
rect 34142 376378 34226 376614
rect 34462 376378 34494 376614
rect 33874 376294 34494 376378
rect 33874 376058 33906 376294
rect 34142 376058 34226 376294
rect 34462 376058 34494 376294
rect 33874 358614 34494 376058
rect 33874 358378 33906 358614
rect 34142 358378 34226 358614
rect 34462 358378 34494 358614
rect 33874 358294 34494 358378
rect 33874 358058 33906 358294
rect 34142 358058 34226 358294
rect 34462 358058 34494 358294
rect 33874 340614 34494 358058
rect 33874 340378 33906 340614
rect 34142 340378 34226 340614
rect 34462 340378 34494 340614
rect 33874 340294 34494 340378
rect 33874 340058 33906 340294
rect 34142 340058 34226 340294
rect 34462 340058 34494 340294
rect 33874 322614 34494 340058
rect 33874 322378 33906 322614
rect 34142 322378 34226 322614
rect 34462 322378 34494 322614
rect 33874 322294 34494 322378
rect 33874 322058 33906 322294
rect 34142 322058 34226 322294
rect 34462 322058 34494 322294
rect 33874 304614 34494 322058
rect 33874 304378 33906 304614
rect 34142 304378 34226 304614
rect 34462 304378 34494 304614
rect 33874 304294 34494 304378
rect 33874 304058 33906 304294
rect 34142 304058 34226 304294
rect 34462 304058 34494 304294
rect 33874 286614 34494 304058
rect 33874 286378 33906 286614
rect 34142 286378 34226 286614
rect 34462 286378 34494 286614
rect 33874 286294 34494 286378
rect 33874 286058 33906 286294
rect 34142 286058 34226 286294
rect 34462 286058 34494 286294
rect 33874 268614 34494 286058
rect 33874 268378 33906 268614
rect 34142 268378 34226 268614
rect 34462 268378 34494 268614
rect 33874 268294 34494 268378
rect 33874 268058 33906 268294
rect 34142 268058 34226 268294
rect 34462 268058 34494 268294
rect 33874 250614 34494 268058
rect 33874 250378 33906 250614
rect 34142 250378 34226 250614
rect 34462 250378 34494 250614
rect 33874 250294 34494 250378
rect 33874 250058 33906 250294
rect 34142 250058 34226 250294
rect 34462 250058 34494 250294
rect 33874 232614 34494 250058
rect 33874 232378 33906 232614
rect 34142 232378 34226 232614
rect 34462 232378 34494 232614
rect 33874 232294 34494 232378
rect 33874 232058 33906 232294
rect 34142 232058 34226 232294
rect 34462 232058 34494 232294
rect 33874 214614 34494 232058
rect 33874 214378 33906 214614
rect 34142 214378 34226 214614
rect 34462 214378 34494 214614
rect 33874 214294 34494 214378
rect 33874 214058 33906 214294
rect 34142 214058 34226 214294
rect 34462 214058 34494 214294
rect 33874 196614 34494 214058
rect 33874 196378 33906 196614
rect 34142 196378 34226 196614
rect 34462 196378 34494 196614
rect 33874 196294 34494 196378
rect 33874 196058 33906 196294
rect 34142 196058 34226 196294
rect 34462 196058 34494 196294
rect 33874 178614 34494 196058
rect 33874 178378 33906 178614
rect 34142 178378 34226 178614
rect 34462 178378 34494 178614
rect 33874 178294 34494 178378
rect 33874 178058 33906 178294
rect 34142 178058 34226 178294
rect 34462 178058 34494 178294
rect 33874 160614 34494 178058
rect 33874 160378 33906 160614
rect 34142 160378 34226 160614
rect 34462 160378 34494 160614
rect 33874 160294 34494 160378
rect 33874 160058 33906 160294
rect 34142 160058 34226 160294
rect 34462 160058 34494 160294
rect 33874 142614 34494 160058
rect 33874 142378 33906 142614
rect 34142 142378 34226 142614
rect 34462 142378 34494 142614
rect 33874 142294 34494 142378
rect 33874 142058 33906 142294
rect 34142 142058 34226 142294
rect 34462 142058 34494 142294
rect 33874 124614 34494 142058
rect 33874 124378 33906 124614
rect 34142 124378 34226 124614
rect 34462 124378 34494 124614
rect 33874 124294 34494 124378
rect 33874 124058 33906 124294
rect 34142 124058 34226 124294
rect 34462 124058 34494 124294
rect 33874 106614 34494 124058
rect 33874 106378 33906 106614
rect 34142 106378 34226 106614
rect 34462 106378 34494 106614
rect 33874 106294 34494 106378
rect 33874 106058 33906 106294
rect 34142 106058 34226 106294
rect 34462 106058 34494 106294
rect 33874 88614 34494 106058
rect 33874 88378 33906 88614
rect 34142 88378 34226 88614
rect 34462 88378 34494 88614
rect 33874 88294 34494 88378
rect 33874 88058 33906 88294
rect 34142 88058 34226 88294
rect 34462 88058 34494 88294
rect 33874 70614 34494 88058
rect 33874 70378 33906 70614
rect 34142 70378 34226 70614
rect 34462 70378 34494 70614
rect 33874 70294 34494 70378
rect 33874 70058 33906 70294
rect 34142 70058 34226 70294
rect 34462 70058 34494 70294
rect 33874 52614 34494 70058
rect 33874 52378 33906 52614
rect 34142 52378 34226 52614
rect 34462 52378 34494 52614
rect 33874 52294 34494 52378
rect 33874 52058 33906 52294
rect 34142 52058 34226 52294
rect 34462 52058 34494 52294
rect 33874 34614 34494 52058
rect 33874 34378 33906 34614
rect 34142 34378 34226 34614
rect 34462 34378 34494 34614
rect 33874 34294 34494 34378
rect 33874 34058 33906 34294
rect 34142 34058 34226 34294
rect 34462 34058 34494 34294
rect 33874 16614 34494 34058
rect 33874 16378 33906 16614
rect 34142 16378 34226 16614
rect 34462 16378 34494 16614
rect 33874 16294 34494 16378
rect 33874 16058 33906 16294
rect 34142 16058 34226 16294
rect 34462 16058 34494 16294
rect 33874 880 34494 16058
rect 40714 461092 41334 464004
rect 40714 460856 40746 461092
rect 40982 460856 41066 461092
rect 41302 460856 41334 461092
rect 40714 460772 41334 460856
rect 40714 460536 40746 460772
rect 40982 460536 41066 460772
rect 41302 460536 41334 460772
rect 40714 455454 41334 460536
rect 40714 455218 40746 455454
rect 40982 455218 41066 455454
rect 41302 455218 41334 455454
rect 40714 455134 41334 455218
rect 40714 454898 40746 455134
rect 40982 454898 41066 455134
rect 41302 454898 41334 455134
rect 40714 437454 41334 454898
rect 40714 437218 40746 437454
rect 40982 437218 41066 437454
rect 41302 437218 41334 437454
rect 40714 437134 41334 437218
rect 40714 436898 40746 437134
rect 40982 436898 41066 437134
rect 41302 436898 41334 437134
rect 40714 419454 41334 436898
rect 40714 419218 40746 419454
rect 40982 419218 41066 419454
rect 41302 419218 41334 419454
rect 40714 419134 41334 419218
rect 40714 418898 40746 419134
rect 40982 418898 41066 419134
rect 41302 418898 41334 419134
rect 40714 401454 41334 418898
rect 40714 401218 40746 401454
rect 40982 401218 41066 401454
rect 41302 401218 41334 401454
rect 40714 401134 41334 401218
rect 40714 400898 40746 401134
rect 40982 400898 41066 401134
rect 41302 400898 41334 401134
rect 40714 383454 41334 400898
rect 40714 383218 40746 383454
rect 40982 383218 41066 383454
rect 41302 383218 41334 383454
rect 40714 383134 41334 383218
rect 40714 382898 40746 383134
rect 40982 382898 41066 383134
rect 41302 382898 41334 383134
rect 40714 365454 41334 382898
rect 40714 365218 40746 365454
rect 40982 365218 41066 365454
rect 41302 365218 41334 365454
rect 40714 365134 41334 365218
rect 40714 364898 40746 365134
rect 40982 364898 41066 365134
rect 41302 364898 41334 365134
rect 40714 347454 41334 364898
rect 40714 347218 40746 347454
rect 40982 347218 41066 347454
rect 41302 347218 41334 347454
rect 40714 347134 41334 347218
rect 40714 346898 40746 347134
rect 40982 346898 41066 347134
rect 41302 346898 41334 347134
rect 40714 329454 41334 346898
rect 40714 329218 40746 329454
rect 40982 329218 41066 329454
rect 41302 329218 41334 329454
rect 40714 329134 41334 329218
rect 40714 328898 40746 329134
rect 40982 328898 41066 329134
rect 41302 328898 41334 329134
rect 40714 311454 41334 328898
rect 40714 311218 40746 311454
rect 40982 311218 41066 311454
rect 41302 311218 41334 311454
rect 40714 311134 41334 311218
rect 40714 310898 40746 311134
rect 40982 310898 41066 311134
rect 41302 310898 41334 311134
rect 40714 293454 41334 310898
rect 40714 293218 40746 293454
rect 40982 293218 41066 293454
rect 41302 293218 41334 293454
rect 40714 293134 41334 293218
rect 40714 292898 40746 293134
rect 40982 292898 41066 293134
rect 41302 292898 41334 293134
rect 40714 275454 41334 292898
rect 40714 275218 40746 275454
rect 40982 275218 41066 275454
rect 41302 275218 41334 275454
rect 40714 275134 41334 275218
rect 40714 274898 40746 275134
rect 40982 274898 41066 275134
rect 41302 274898 41334 275134
rect 40714 257454 41334 274898
rect 40714 257218 40746 257454
rect 40982 257218 41066 257454
rect 41302 257218 41334 257454
rect 40714 257134 41334 257218
rect 40714 256898 40746 257134
rect 40982 256898 41066 257134
rect 41302 256898 41334 257134
rect 40714 239454 41334 256898
rect 40714 239218 40746 239454
rect 40982 239218 41066 239454
rect 41302 239218 41334 239454
rect 40714 239134 41334 239218
rect 40714 238898 40746 239134
rect 40982 238898 41066 239134
rect 41302 238898 41334 239134
rect 40714 221454 41334 238898
rect 40714 221218 40746 221454
rect 40982 221218 41066 221454
rect 41302 221218 41334 221454
rect 40714 221134 41334 221218
rect 40714 220898 40746 221134
rect 40982 220898 41066 221134
rect 41302 220898 41334 221134
rect 40714 203454 41334 220898
rect 40714 203218 40746 203454
rect 40982 203218 41066 203454
rect 41302 203218 41334 203454
rect 40714 203134 41334 203218
rect 40714 202898 40746 203134
rect 40982 202898 41066 203134
rect 41302 202898 41334 203134
rect 40714 185454 41334 202898
rect 40714 185218 40746 185454
rect 40982 185218 41066 185454
rect 41302 185218 41334 185454
rect 40714 185134 41334 185218
rect 40714 184898 40746 185134
rect 40982 184898 41066 185134
rect 41302 184898 41334 185134
rect 40714 167454 41334 184898
rect 40714 167218 40746 167454
rect 40982 167218 41066 167454
rect 41302 167218 41334 167454
rect 40714 167134 41334 167218
rect 40714 166898 40746 167134
rect 40982 166898 41066 167134
rect 41302 166898 41334 167134
rect 40714 149454 41334 166898
rect 40714 149218 40746 149454
rect 40982 149218 41066 149454
rect 41302 149218 41334 149454
rect 40714 149134 41334 149218
rect 40714 148898 40746 149134
rect 40982 148898 41066 149134
rect 41302 148898 41334 149134
rect 40714 131454 41334 148898
rect 40714 131218 40746 131454
rect 40982 131218 41066 131454
rect 41302 131218 41334 131454
rect 40714 131134 41334 131218
rect 40714 130898 40746 131134
rect 40982 130898 41066 131134
rect 41302 130898 41334 131134
rect 40714 113454 41334 130898
rect 40714 113218 40746 113454
rect 40982 113218 41066 113454
rect 41302 113218 41334 113454
rect 40714 113134 41334 113218
rect 40714 112898 40746 113134
rect 40982 112898 41066 113134
rect 41302 112898 41334 113134
rect 40714 95454 41334 112898
rect 40714 95218 40746 95454
rect 40982 95218 41066 95454
rect 41302 95218 41334 95454
rect 40714 95134 41334 95218
rect 40714 94898 40746 95134
rect 40982 94898 41066 95134
rect 41302 94898 41334 95134
rect 40714 77454 41334 94898
rect 40714 77218 40746 77454
rect 40982 77218 41066 77454
rect 41302 77218 41334 77454
rect 40714 77134 41334 77218
rect 40714 76898 40746 77134
rect 40982 76898 41066 77134
rect 41302 76898 41334 77134
rect 40714 59454 41334 76898
rect 40714 59218 40746 59454
rect 40982 59218 41066 59454
rect 41302 59218 41334 59454
rect 40714 59134 41334 59218
rect 40714 58898 40746 59134
rect 40982 58898 41066 59134
rect 41302 58898 41334 59134
rect 40714 41454 41334 58898
rect 40714 41218 40746 41454
rect 40982 41218 41066 41454
rect 41302 41218 41334 41454
rect 40714 41134 41334 41218
rect 40714 40898 40746 41134
rect 40982 40898 41066 41134
rect 41302 40898 41334 41134
rect 40714 23454 41334 40898
rect 40714 23218 40746 23454
rect 40982 23218 41066 23454
rect 41302 23218 41334 23454
rect 40714 23134 41334 23218
rect 40714 22898 40746 23134
rect 40982 22898 41066 23134
rect 41302 22898 41334 23134
rect 40714 5454 41334 22898
rect 40714 5218 40746 5454
rect 40982 5218 41066 5454
rect 41302 5218 41334 5454
rect 40714 5134 41334 5218
rect 40714 4898 40746 5134
rect 40982 4898 41066 5134
rect 41302 4898 41334 5134
rect 40714 880 41334 4898
rect 44434 462052 45054 464004
rect 44434 461816 44466 462052
rect 44702 461816 44786 462052
rect 45022 461816 45054 462052
rect 44434 461732 45054 461816
rect 44434 461496 44466 461732
rect 44702 461496 44786 461732
rect 45022 461496 45054 461732
rect 44434 441174 45054 461496
rect 44434 440938 44466 441174
rect 44702 440938 44786 441174
rect 45022 440938 45054 441174
rect 44434 440854 45054 440938
rect 44434 440618 44466 440854
rect 44702 440618 44786 440854
rect 45022 440618 45054 440854
rect 44434 423174 45054 440618
rect 44434 422938 44466 423174
rect 44702 422938 44786 423174
rect 45022 422938 45054 423174
rect 44434 422854 45054 422938
rect 44434 422618 44466 422854
rect 44702 422618 44786 422854
rect 45022 422618 45054 422854
rect 44434 405174 45054 422618
rect 44434 404938 44466 405174
rect 44702 404938 44786 405174
rect 45022 404938 45054 405174
rect 44434 404854 45054 404938
rect 44434 404618 44466 404854
rect 44702 404618 44786 404854
rect 45022 404618 45054 404854
rect 44434 387174 45054 404618
rect 44434 386938 44466 387174
rect 44702 386938 44786 387174
rect 45022 386938 45054 387174
rect 44434 386854 45054 386938
rect 44434 386618 44466 386854
rect 44702 386618 44786 386854
rect 45022 386618 45054 386854
rect 44434 369174 45054 386618
rect 44434 368938 44466 369174
rect 44702 368938 44786 369174
rect 45022 368938 45054 369174
rect 44434 368854 45054 368938
rect 44434 368618 44466 368854
rect 44702 368618 44786 368854
rect 45022 368618 45054 368854
rect 44434 351174 45054 368618
rect 44434 350938 44466 351174
rect 44702 350938 44786 351174
rect 45022 350938 45054 351174
rect 44434 350854 45054 350938
rect 44434 350618 44466 350854
rect 44702 350618 44786 350854
rect 45022 350618 45054 350854
rect 44434 333174 45054 350618
rect 44434 332938 44466 333174
rect 44702 332938 44786 333174
rect 45022 332938 45054 333174
rect 44434 332854 45054 332938
rect 44434 332618 44466 332854
rect 44702 332618 44786 332854
rect 45022 332618 45054 332854
rect 44434 315174 45054 332618
rect 44434 314938 44466 315174
rect 44702 314938 44786 315174
rect 45022 314938 45054 315174
rect 44434 314854 45054 314938
rect 44434 314618 44466 314854
rect 44702 314618 44786 314854
rect 45022 314618 45054 314854
rect 44434 297174 45054 314618
rect 44434 296938 44466 297174
rect 44702 296938 44786 297174
rect 45022 296938 45054 297174
rect 44434 296854 45054 296938
rect 44434 296618 44466 296854
rect 44702 296618 44786 296854
rect 45022 296618 45054 296854
rect 44434 279174 45054 296618
rect 44434 278938 44466 279174
rect 44702 278938 44786 279174
rect 45022 278938 45054 279174
rect 44434 278854 45054 278938
rect 44434 278618 44466 278854
rect 44702 278618 44786 278854
rect 45022 278618 45054 278854
rect 44434 261174 45054 278618
rect 44434 260938 44466 261174
rect 44702 260938 44786 261174
rect 45022 260938 45054 261174
rect 44434 260854 45054 260938
rect 44434 260618 44466 260854
rect 44702 260618 44786 260854
rect 45022 260618 45054 260854
rect 44434 243174 45054 260618
rect 44434 242938 44466 243174
rect 44702 242938 44786 243174
rect 45022 242938 45054 243174
rect 44434 242854 45054 242938
rect 44434 242618 44466 242854
rect 44702 242618 44786 242854
rect 45022 242618 45054 242854
rect 44434 225174 45054 242618
rect 44434 224938 44466 225174
rect 44702 224938 44786 225174
rect 45022 224938 45054 225174
rect 44434 224854 45054 224938
rect 44434 224618 44466 224854
rect 44702 224618 44786 224854
rect 45022 224618 45054 224854
rect 44434 207174 45054 224618
rect 44434 206938 44466 207174
rect 44702 206938 44786 207174
rect 45022 206938 45054 207174
rect 44434 206854 45054 206938
rect 44434 206618 44466 206854
rect 44702 206618 44786 206854
rect 45022 206618 45054 206854
rect 44434 189174 45054 206618
rect 44434 188938 44466 189174
rect 44702 188938 44786 189174
rect 45022 188938 45054 189174
rect 44434 188854 45054 188938
rect 44434 188618 44466 188854
rect 44702 188618 44786 188854
rect 45022 188618 45054 188854
rect 44434 171174 45054 188618
rect 44434 170938 44466 171174
rect 44702 170938 44786 171174
rect 45022 170938 45054 171174
rect 44434 170854 45054 170938
rect 44434 170618 44466 170854
rect 44702 170618 44786 170854
rect 45022 170618 45054 170854
rect 44434 153174 45054 170618
rect 44434 152938 44466 153174
rect 44702 152938 44786 153174
rect 45022 152938 45054 153174
rect 44434 152854 45054 152938
rect 44434 152618 44466 152854
rect 44702 152618 44786 152854
rect 45022 152618 45054 152854
rect 44434 135174 45054 152618
rect 44434 134938 44466 135174
rect 44702 134938 44786 135174
rect 45022 134938 45054 135174
rect 44434 134854 45054 134938
rect 44434 134618 44466 134854
rect 44702 134618 44786 134854
rect 45022 134618 45054 134854
rect 44434 117174 45054 134618
rect 44434 116938 44466 117174
rect 44702 116938 44786 117174
rect 45022 116938 45054 117174
rect 44434 116854 45054 116938
rect 44434 116618 44466 116854
rect 44702 116618 44786 116854
rect 45022 116618 45054 116854
rect 44434 99174 45054 116618
rect 44434 98938 44466 99174
rect 44702 98938 44786 99174
rect 45022 98938 45054 99174
rect 44434 98854 45054 98938
rect 44434 98618 44466 98854
rect 44702 98618 44786 98854
rect 45022 98618 45054 98854
rect 44434 81174 45054 98618
rect 44434 80938 44466 81174
rect 44702 80938 44786 81174
rect 45022 80938 45054 81174
rect 44434 80854 45054 80938
rect 44434 80618 44466 80854
rect 44702 80618 44786 80854
rect 45022 80618 45054 80854
rect 44434 63174 45054 80618
rect 44434 62938 44466 63174
rect 44702 62938 44786 63174
rect 45022 62938 45054 63174
rect 44434 62854 45054 62938
rect 44434 62618 44466 62854
rect 44702 62618 44786 62854
rect 45022 62618 45054 62854
rect 44434 45174 45054 62618
rect 44434 44938 44466 45174
rect 44702 44938 44786 45174
rect 45022 44938 45054 45174
rect 44434 44854 45054 44938
rect 44434 44618 44466 44854
rect 44702 44618 44786 44854
rect 45022 44618 45054 44854
rect 44434 27174 45054 44618
rect 44434 26938 44466 27174
rect 44702 26938 44786 27174
rect 45022 26938 45054 27174
rect 44434 26854 45054 26938
rect 44434 26618 44466 26854
rect 44702 26618 44786 26854
rect 45022 26618 45054 26854
rect 44434 9174 45054 26618
rect 44434 8938 44466 9174
rect 44702 8938 44786 9174
rect 45022 8938 45054 9174
rect 44434 8854 45054 8938
rect 44434 8618 44466 8854
rect 44702 8618 44786 8854
rect 45022 8618 45054 8854
rect 44434 880 45054 8618
rect 48154 463012 48774 464004
rect 48154 462776 48186 463012
rect 48422 462776 48506 463012
rect 48742 462776 48774 463012
rect 48154 462692 48774 462776
rect 48154 462456 48186 462692
rect 48422 462456 48506 462692
rect 48742 462456 48774 462692
rect 48154 444894 48774 462456
rect 48154 444658 48186 444894
rect 48422 444658 48506 444894
rect 48742 444658 48774 444894
rect 48154 444574 48774 444658
rect 48154 444338 48186 444574
rect 48422 444338 48506 444574
rect 48742 444338 48774 444574
rect 48154 426894 48774 444338
rect 48154 426658 48186 426894
rect 48422 426658 48506 426894
rect 48742 426658 48774 426894
rect 48154 426574 48774 426658
rect 48154 426338 48186 426574
rect 48422 426338 48506 426574
rect 48742 426338 48774 426574
rect 48154 408894 48774 426338
rect 48154 408658 48186 408894
rect 48422 408658 48506 408894
rect 48742 408658 48774 408894
rect 48154 408574 48774 408658
rect 48154 408338 48186 408574
rect 48422 408338 48506 408574
rect 48742 408338 48774 408574
rect 48154 390894 48774 408338
rect 48154 390658 48186 390894
rect 48422 390658 48506 390894
rect 48742 390658 48774 390894
rect 48154 390574 48774 390658
rect 48154 390338 48186 390574
rect 48422 390338 48506 390574
rect 48742 390338 48774 390574
rect 48154 372894 48774 390338
rect 48154 372658 48186 372894
rect 48422 372658 48506 372894
rect 48742 372658 48774 372894
rect 48154 372574 48774 372658
rect 48154 372338 48186 372574
rect 48422 372338 48506 372574
rect 48742 372338 48774 372574
rect 48154 354894 48774 372338
rect 48154 354658 48186 354894
rect 48422 354658 48506 354894
rect 48742 354658 48774 354894
rect 48154 354574 48774 354658
rect 48154 354338 48186 354574
rect 48422 354338 48506 354574
rect 48742 354338 48774 354574
rect 48154 336894 48774 354338
rect 48154 336658 48186 336894
rect 48422 336658 48506 336894
rect 48742 336658 48774 336894
rect 48154 336574 48774 336658
rect 48154 336338 48186 336574
rect 48422 336338 48506 336574
rect 48742 336338 48774 336574
rect 48154 318894 48774 336338
rect 48154 318658 48186 318894
rect 48422 318658 48506 318894
rect 48742 318658 48774 318894
rect 48154 318574 48774 318658
rect 48154 318338 48186 318574
rect 48422 318338 48506 318574
rect 48742 318338 48774 318574
rect 48154 300894 48774 318338
rect 48154 300658 48186 300894
rect 48422 300658 48506 300894
rect 48742 300658 48774 300894
rect 48154 300574 48774 300658
rect 48154 300338 48186 300574
rect 48422 300338 48506 300574
rect 48742 300338 48774 300574
rect 48154 282894 48774 300338
rect 48154 282658 48186 282894
rect 48422 282658 48506 282894
rect 48742 282658 48774 282894
rect 48154 282574 48774 282658
rect 48154 282338 48186 282574
rect 48422 282338 48506 282574
rect 48742 282338 48774 282574
rect 48154 264894 48774 282338
rect 48154 264658 48186 264894
rect 48422 264658 48506 264894
rect 48742 264658 48774 264894
rect 48154 264574 48774 264658
rect 48154 264338 48186 264574
rect 48422 264338 48506 264574
rect 48742 264338 48774 264574
rect 48154 246894 48774 264338
rect 48154 246658 48186 246894
rect 48422 246658 48506 246894
rect 48742 246658 48774 246894
rect 48154 246574 48774 246658
rect 48154 246338 48186 246574
rect 48422 246338 48506 246574
rect 48742 246338 48774 246574
rect 48154 228894 48774 246338
rect 48154 228658 48186 228894
rect 48422 228658 48506 228894
rect 48742 228658 48774 228894
rect 48154 228574 48774 228658
rect 48154 228338 48186 228574
rect 48422 228338 48506 228574
rect 48742 228338 48774 228574
rect 48154 210894 48774 228338
rect 48154 210658 48186 210894
rect 48422 210658 48506 210894
rect 48742 210658 48774 210894
rect 48154 210574 48774 210658
rect 48154 210338 48186 210574
rect 48422 210338 48506 210574
rect 48742 210338 48774 210574
rect 48154 192894 48774 210338
rect 48154 192658 48186 192894
rect 48422 192658 48506 192894
rect 48742 192658 48774 192894
rect 48154 192574 48774 192658
rect 48154 192338 48186 192574
rect 48422 192338 48506 192574
rect 48742 192338 48774 192574
rect 48154 174894 48774 192338
rect 48154 174658 48186 174894
rect 48422 174658 48506 174894
rect 48742 174658 48774 174894
rect 48154 174574 48774 174658
rect 48154 174338 48186 174574
rect 48422 174338 48506 174574
rect 48742 174338 48774 174574
rect 48154 156894 48774 174338
rect 48154 156658 48186 156894
rect 48422 156658 48506 156894
rect 48742 156658 48774 156894
rect 48154 156574 48774 156658
rect 48154 156338 48186 156574
rect 48422 156338 48506 156574
rect 48742 156338 48774 156574
rect 48154 138894 48774 156338
rect 48154 138658 48186 138894
rect 48422 138658 48506 138894
rect 48742 138658 48774 138894
rect 48154 138574 48774 138658
rect 48154 138338 48186 138574
rect 48422 138338 48506 138574
rect 48742 138338 48774 138574
rect 48154 120894 48774 138338
rect 48154 120658 48186 120894
rect 48422 120658 48506 120894
rect 48742 120658 48774 120894
rect 48154 120574 48774 120658
rect 48154 120338 48186 120574
rect 48422 120338 48506 120574
rect 48742 120338 48774 120574
rect 48154 102894 48774 120338
rect 48154 102658 48186 102894
rect 48422 102658 48506 102894
rect 48742 102658 48774 102894
rect 48154 102574 48774 102658
rect 48154 102338 48186 102574
rect 48422 102338 48506 102574
rect 48742 102338 48774 102574
rect 48154 84894 48774 102338
rect 48154 84658 48186 84894
rect 48422 84658 48506 84894
rect 48742 84658 48774 84894
rect 48154 84574 48774 84658
rect 48154 84338 48186 84574
rect 48422 84338 48506 84574
rect 48742 84338 48774 84574
rect 48154 66894 48774 84338
rect 48154 66658 48186 66894
rect 48422 66658 48506 66894
rect 48742 66658 48774 66894
rect 48154 66574 48774 66658
rect 48154 66338 48186 66574
rect 48422 66338 48506 66574
rect 48742 66338 48774 66574
rect 48154 48894 48774 66338
rect 48154 48658 48186 48894
rect 48422 48658 48506 48894
rect 48742 48658 48774 48894
rect 48154 48574 48774 48658
rect 48154 48338 48186 48574
rect 48422 48338 48506 48574
rect 48742 48338 48774 48574
rect 48154 30894 48774 48338
rect 48154 30658 48186 30894
rect 48422 30658 48506 30894
rect 48742 30658 48774 30894
rect 48154 30574 48774 30658
rect 48154 30338 48186 30574
rect 48422 30338 48506 30574
rect 48742 30338 48774 30574
rect 48154 12894 48774 30338
rect 48154 12658 48186 12894
rect 48422 12658 48506 12894
rect 48742 12658 48774 12894
rect 48154 12574 48774 12658
rect 48154 12338 48186 12574
rect 48422 12338 48506 12574
rect 48742 12338 48774 12574
rect 4939 0 9719 638
rect 14918 0 19698 638
rect 28939 0 33719 638
rect 38918 0 43698 638
rect -1596 -1092 -1564 -856
rect -1328 -1092 -1244 -856
rect -1008 -1092 -976 -856
rect -1596 -1176 -976 -1092
rect -1596 -1412 -1564 -1176
rect -1328 -1412 -1244 -1176
rect -1008 -1412 -976 -1176
rect -1596 -1444 -976 -1412
rect -2556 -2052 -2524 -1816
rect -2288 -2052 -2204 -1816
rect -1968 -2052 -1936 -1816
rect -2556 -2136 -1936 -2052
rect -2556 -2372 -2524 -2136
rect -2288 -2372 -2204 -2136
rect -1968 -2372 -1936 -2136
rect -2556 -2404 -1936 -2372
rect -3516 -3012 -3484 -2776
rect -3248 -3012 -3164 -2776
rect -2928 -3012 -2896 -2776
rect -3516 -3096 -2896 -3012
rect -3516 -3332 -3484 -3096
rect -3248 -3332 -3164 -3096
rect -2928 -3332 -2896 -3096
rect -3516 -3364 -2896 -3332
rect 48154 -2776 48774 12338
rect 48154 -3012 48186 -2776
rect 48422 -3012 48506 -2776
rect 48742 -3012 48774 -2776
rect 48154 -3096 48774 -3012
rect 48154 -3332 48186 -3096
rect 48422 -3332 48506 -3096
rect 48742 -3332 48774 -3096
rect -4476 -3972 -4444 -3736
rect -4208 -3972 -4124 -3736
rect -3888 -3972 -3856 -3736
rect -4476 -4056 -3856 -3972
rect -4476 -4292 -4444 -4056
rect -4208 -4292 -4124 -4056
rect -3888 -4292 -3856 -4056
rect -4476 -4324 -3856 -4292
rect 48154 -4324 48774 -3332
rect 51874 463972 52494 464004
rect 51874 463736 51906 463972
rect 52142 463736 52226 463972
rect 52462 463736 52494 463972
rect 51874 463652 52494 463736
rect 51874 463416 51906 463652
rect 52142 463416 52226 463652
rect 52462 463416 52494 463652
rect 51874 448614 52494 463416
rect 51874 448378 51906 448614
rect 52142 448378 52226 448614
rect 52462 448378 52494 448614
rect 51874 448294 52494 448378
rect 51874 448058 51906 448294
rect 52142 448058 52226 448294
rect 52462 448058 52494 448294
rect 51874 430614 52494 448058
rect 51874 430378 51906 430614
rect 52142 430378 52226 430614
rect 52462 430378 52494 430614
rect 51874 430294 52494 430378
rect 51874 430058 51906 430294
rect 52142 430058 52226 430294
rect 52462 430058 52494 430294
rect 51874 412614 52494 430058
rect 51874 412378 51906 412614
rect 52142 412378 52226 412614
rect 52462 412378 52494 412614
rect 51874 412294 52494 412378
rect 51874 412058 51906 412294
rect 52142 412058 52226 412294
rect 52462 412058 52494 412294
rect 51874 394614 52494 412058
rect 51874 394378 51906 394614
rect 52142 394378 52226 394614
rect 52462 394378 52494 394614
rect 51874 394294 52494 394378
rect 51874 394058 51906 394294
rect 52142 394058 52226 394294
rect 52462 394058 52494 394294
rect 51874 376614 52494 394058
rect 51874 376378 51906 376614
rect 52142 376378 52226 376614
rect 52462 376378 52494 376614
rect 51874 376294 52494 376378
rect 51874 376058 51906 376294
rect 52142 376058 52226 376294
rect 52462 376058 52494 376294
rect 51874 358614 52494 376058
rect 51874 358378 51906 358614
rect 52142 358378 52226 358614
rect 52462 358378 52494 358614
rect 51874 358294 52494 358378
rect 51874 358058 51906 358294
rect 52142 358058 52226 358294
rect 52462 358058 52494 358294
rect 51874 340614 52494 358058
rect 51874 340378 51906 340614
rect 52142 340378 52226 340614
rect 52462 340378 52494 340614
rect 51874 340294 52494 340378
rect 51874 340058 51906 340294
rect 52142 340058 52226 340294
rect 52462 340058 52494 340294
rect 51874 322614 52494 340058
rect 51874 322378 51906 322614
rect 52142 322378 52226 322614
rect 52462 322378 52494 322614
rect 51874 322294 52494 322378
rect 51874 322058 51906 322294
rect 52142 322058 52226 322294
rect 52462 322058 52494 322294
rect 51874 304614 52494 322058
rect 51874 304378 51906 304614
rect 52142 304378 52226 304614
rect 52462 304378 52494 304614
rect 51874 304294 52494 304378
rect 51874 304058 51906 304294
rect 52142 304058 52226 304294
rect 52462 304058 52494 304294
rect 51874 286614 52494 304058
rect 51874 286378 51906 286614
rect 52142 286378 52226 286614
rect 52462 286378 52494 286614
rect 51874 286294 52494 286378
rect 51874 286058 51906 286294
rect 52142 286058 52226 286294
rect 52462 286058 52494 286294
rect 51874 268614 52494 286058
rect 51874 268378 51906 268614
rect 52142 268378 52226 268614
rect 52462 268378 52494 268614
rect 51874 268294 52494 268378
rect 51874 268058 51906 268294
rect 52142 268058 52226 268294
rect 52462 268058 52494 268294
rect 51874 250614 52494 268058
rect 51874 250378 51906 250614
rect 52142 250378 52226 250614
rect 52462 250378 52494 250614
rect 51874 250294 52494 250378
rect 51874 250058 51906 250294
rect 52142 250058 52226 250294
rect 52462 250058 52494 250294
rect 51874 232614 52494 250058
rect 51874 232378 51906 232614
rect 52142 232378 52226 232614
rect 52462 232378 52494 232614
rect 51874 232294 52494 232378
rect 51874 232058 51906 232294
rect 52142 232058 52226 232294
rect 52462 232058 52494 232294
rect 51874 214614 52494 232058
rect 51874 214378 51906 214614
rect 52142 214378 52226 214614
rect 52462 214378 52494 214614
rect 51874 214294 52494 214378
rect 51874 214058 51906 214294
rect 52142 214058 52226 214294
rect 52462 214058 52494 214294
rect 51874 196614 52494 214058
rect 51874 196378 51906 196614
rect 52142 196378 52226 196614
rect 52462 196378 52494 196614
rect 51874 196294 52494 196378
rect 51874 196058 51906 196294
rect 52142 196058 52226 196294
rect 52462 196058 52494 196294
rect 51874 178614 52494 196058
rect 51874 178378 51906 178614
rect 52142 178378 52226 178614
rect 52462 178378 52494 178614
rect 51874 178294 52494 178378
rect 51874 178058 51906 178294
rect 52142 178058 52226 178294
rect 52462 178058 52494 178294
rect 51874 160614 52494 178058
rect 51874 160378 51906 160614
rect 52142 160378 52226 160614
rect 52462 160378 52494 160614
rect 51874 160294 52494 160378
rect 51874 160058 51906 160294
rect 52142 160058 52226 160294
rect 52462 160058 52494 160294
rect 51874 142614 52494 160058
rect 51874 142378 51906 142614
rect 52142 142378 52226 142614
rect 52462 142378 52494 142614
rect 51874 142294 52494 142378
rect 51874 142058 51906 142294
rect 52142 142058 52226 142294
rect 52462 142058 52494 142294
rect 51874 124614 52494 142058
rect 51874 124378 51906 124614
rect 52142 124378 52226 124614
rect 52462 124378 52494 124614
rect 51874 124294 52494 124378
rect 51874 124058 51906 124294
rect 52142 124058 52226 124294
rect 52462 124058 52494 124294
rect 51874 106614 52494 124058
rect 51874 106378 51906 106614
rect 52142 106378 52226 106614
rect 52462 106378 52494 106614
rect 51874 106294 52494 106378
rect 51874 106058 51906 106294
rect 52142 106058 52226 106294
rect 52462 106058 52494 106294
rect 51874 88614 52494 106058
rect 51874 88378 51906 88614
rect 52142 88378 52226 88614
rect 52462 88378 52494 88614
rect 51874 88294 52494 88378
rect 51874 88058 51906 88294
rect 52142 88058 52226 88294
rect 52462 88058 52494 88294
rect 51874 70614 52494 88058
rect 51874 70378 51906 70614
rect 52142 70378 52226 70614
rect 52462 70378 52494 70614
rect 51874 70294 52494 70378
rect 51874 70058 51906 70294
rect 52142 70058 52226 70294
rect 52462 70058 52494 70294
rect 51874 52614 52494 70058
rect 51874 52378 51906 52614
rect 52142 52378 52226 52614
rect 52462 52378 52494 52614
rect 51874 52294 52494 52378
rect 51874 52058 51906 52294
rect 52142 52058 52226 52294
rect 52462 52058 52494 52294
rect 51874 34614 52494 52058
rect 51874 34378 51906 34614
rect 52142 34378 52226 34614
rect 52462 34378 52494 34614
rect 51874 34294 52494 34378
rect 51874 34058 51906 34294
rect 52142 34058 52226 34294
rect 52462 34058 52494 34294
rect 51874 16614 52494 34058
rect 51874 16378 51906 16614
rect 52142 16378 52226 16614
rect 52462 16378 52494 16614
rect 51874 16294 52494 16378
rect 51874 16058 51906 16294
rect 52142 16058 52226 16294
rect 52462 16058 52494 16294
rect 51874 -3736 52494 16058
rect 51874 -3972 51906 -3736
rect 52142 -3972 52226 -3736
rect 52462 -3972 52494 -3736
rect 51874 -4056 52494 -3972
rect 51874 -4292 51906 -4056
rect 52142 -4292 52226 -4056
rect 52462 -4292 52494 -4056
rect 51874 -4324 52494 -4292
rect 58714 461092 59334 464004
rect 58714 460856 58746 461092
rect 58982 460856 59066 461092
rect 59302 460856 59334 461092
rect 58714 460772 59334 460856
rect 58714 460536 58746 460772
rect 58982 460536 59066 460772
rect 59302 460536 59334 460772
rect 58714 455454 59334 460536
rect 58714 455218 58746 455454
rect 58982 455218 59066 455454
rect 59302 455218 59334 455454
rect 58714 455134 59334 455218
rect 58714 454898 58746 455134
rect 58982 454898 59066 455134
rect 59302 454898 59334 455134
rect 58714 437454 59334 454898
rect 58714 437218 58746 437454
rect 58982 437218 59066 437454
rect 59302 437218 59334 437454
rect 58714 437134 59334 437218
rect 58714 436898 58746 437134
rect 58982 436898 59066 437134
rect 59302 436898 59334 437134
rect 58714 419454 59334 436898
rect 58714 419218 58746 419454
rect 58982 419218 59066 419454
rect 59302 419218 59334 419454
rect 58714 419134 59334 419218
rect 58714 418898 58746 419134
rect 58982 418898 59066 419134
rect 59302 418898 59334 419134
rect 58714 401454 59334 418898
rect 58714 401218 58746 401454
rect 58982 401218 59066 401454
rect 59302 401218 59334 401454
rect 58714 401134 59334 401218
rect 58714 400898 58746 401134
rect 58982 400898 59066 401134
rect 59302 400898 59334 401134
rect 58714 383454 59334 400898
rect 58714 383218 58746 383454
rect 58982 383218 59066 383454
rect 59302 383218 59334 383454
rect 58714 383134 59334 383218
rect 58714 382898 58746 383134
rect 58982 382898 59066 383134
rect 59302 382898 59334 383134
rect 58714 365454 59334 382898
rect 58714 365218 58746 365454
rect 58982 365218 59066 365454
rect 59302 365218 59334 365454
rect 58714 365134 59334 365218
rect 58714 364898 58746 365134
rect 58982 364898 59066 365134
rect 59302 364898 59334 365134
rect 58714 347454 59334 364898
rect 58714 347218 58746 347454
rect 58982 347218 59066 347454
rect 59302 347218 59334 347454
rect 58714 347134 59334 347218
rect 58714 346898 58746 347134
rect 58982 346898 59066 347134
rect 59302 346898 59334 347134
rect 58714 329454 59334 346898
rect 58714 329218 58746 329454
rect 58982 329218 59066 329454
rect 59302 329218 59334 329454
rect 58714 329134 59334 329218
rect 58714 328898 58746 329134
rect 58982 328898 59066 329134
rect 59302 328898 59334 329134
rect 58714 311454 59334 328898
rect 58714 311218 58746 311454
rect 58982 311218 59066 311454
rect 59302 311218 59334 311454
rect 58714 311134 59334 311218
rect 58714 310898 58746 311134
rect 58982 310898 59066 311134
rect 59302 310898 59334 311134
rect 58714 293454 59334 310898
rect 58714 293218 58746 293454
rect 58982 293218 59066 293454
rect 59302 293218 59334 293454
rect 58714 293134 59334 293218
rect 58714 292898 58746 293134
rect 58982 292898 59066 293134
rect 59302 292898 59334 293134
rect 58714 275454 59334 292898
rect 58714 275218 58746 275454
rect 58982 275218 59066 275454
rect 59302 275218 59334 275454
rect 58714 275134 59334 275218
rect 58714 274898 58746 275134
rect 58982 274898 59066 275134
rect 59302 274898 59334 275134
rect 58714 257454 59334 274898
rect 58714 257218 58746 257454
rect 58982 257218 59066 257454
rect 59302 257218 59334 257454
rect 58714 257134 59334 257218
rect 58714 256898 58746 257134
rect 58982 256898 59066 257134
rect 59302 256898 59334 257134
rect 58714 239454 59334 256898
rect 58714 239218 58746 239454
rect 58982 239218 59066 239454
rect 59302 239218 59334 239454
rect 58714 239134 59334 239218
rect 58714 238898 58746 239134
rect 58982 238898 59066 239134
rect 59302 238898 59334 239134
rect 58714 221454 59334 238898
rect 58714 221218 58746 221454
rect 58982 221218 59066 221454
rect 59302 221218 59334 221454
rect 58714 221134 59334 221218
rect 58714 220898 58746 221134
rect 58982 220898 59066 221134
rect 59302 220898 59334 221134
rect 58714 203454 59334 220898
rect 58714 203218 58746 203454
rect 58982 203218 59066 203454
rect 59302 203218 59334 203454
rect 58714 203134 59334 203218
rect 58714 202898 58746 203134
rect 58982 202898 59066 203134
rect 59302 202898 59334 203134
rect 58714 185454 59334 202898
rect 58714 185218 58746 185454
rect 58982 185218 59066 185454
rect 59302 185218 59334 185454
rect 58714 185134 59334 185218
rect 58714 184898 58746 185134
rect 58982 184898 59066 185134
rect 59302 184898 59334 185134
rect 58714 167454 59334 184898
rect 58714 167218 58746 167454
rect 58982 167218 59066 167454
rect 59302 167218 59334 167454
rect 58714 167134 59334 167218
rect 58714 166898 58746 167134
rect 58982 166898 59066 167134
rect 59302 166898 59334 167134
rect 58714 149454 59334 166898
rect 58714 149218 58746 149454
rect 58982 149218 59066 149454
rect 59302 149218 59334 149454
rect 58714 149134 59334 149218
rect 58714 148898 58746 149134
rect 58982 148898 59066 149134
rect 59302 148898 59334 149134
rect 58714 131454 59334 148898
rect 58714 131218 58746 131454
rect 58982 131218 59066 131454
rect 59302 131218 59334 131454
rect 58714 131134 59334 131218
rect 58714 130898 58746 131134
rect 58982 130898 59066 131134
rect 59302 130898 59334 131134
rect 58714 113454 59334 130898
rect 58714 113218 58746 113454
rect 58982 113218 59066 113454
rect 59302 113218 59334 113454
rect 58714 113134 59334 113218
rect 58714 112898 58746 113134
rect 58982 112898 59066 113134
rect 59302 112898 59334 113134
rect 58714 95454 59334 112898
rect 58714 95218 58746 95454
rect 58982 95218 59066 95454
rect 59302 95218 59334 95454
rect 58714 95134 59334 95218
rect 58714 94898 58746 95134
rect 58982 94898 59066 95134
rect 59302 94898 59334 95134
rect 58714 77454 59334 94898
rect 58714 77218 58746 77454
rect 58982 77218 59066 77454
rect 59302 77218 59334 77454
rect 58714 77134 59334 77218
rect 58714 76898 58746 77134
rect 58982 76898 59066 77134
rect 59302 76898 59334 77134
rect 58714 59454 59334 76898
rect 58714 59218 58746 59454
rect 58982 59218 59066 59454
rect 59302 59218 59334 59454
rect 58714 59134 59334 59218
rect 58714 58898 58746 59134
rect 58982 58898 59066 59134
rect 59302 58898 59334 59134
rect 58714 41454 59334 58898
rect 58714 41218 58746 41454
rect 58982 41218 59066 41454
rect 59302 41218 59334 41454
rect 58714 41134 59334 41218
rect 58714 40898 58746 41134
rect 58982 40898 59066 41134
rect 59302 40898 59334 41134
rect 58714 23454 59334 40898
rect 58714 23218 58746 23454
rect 58982 23218 59066 23454
rect 59302 23218 59334 23454
rect 58714 23134 59334 23218
rect 58714 22898 58746 23134
rect 58982 22898 59066 23134
rect 59302 22898 59334 23134
rect 58714 5454 59334 22898
rect 58714 5218 58746 5454
rect 58982 5218 59066 5454
rect 59302 5218 59334 5454
rect 58714 5134 59334 5218
rect 58714 4898 58746 5134
rect 58982 4898 59066 5134
rect 59302 4898 59334 5134
rect 58714 -856 59334 4898
rect 58714 -1092 58746 -856
rect 58982 -1092 59066 -856
rect 59302 -1092 59334 -856
rect 58714 -1176 59334 -1092
rect 58714 -1412 58746 -1176
rect 58982 -1412 59066 -1176
rect 59302 -1412 59334 -1176
rect 58714 -4324 59334 -1412
rect 62434 462052 63054 464004
rect 62434 461816 62466 462052
rect 62702 461816 62786 462052
rect 63022 461816 63054 462052
rect 62434 461732 63054 461816
rect 62434 461496 62466 461732
rect 62702 461496 62786 461732
rect 63022 461496 63054 461732
rect 62434 441174 63054 461496
rect 62434 440938 62466 441174
rect 62702 440938 62786 441174
rect 63022 440938 63054 441174
rect 62434 440854 63054 440938
rect 62434 440618 62466 440854
rect 62702 440618 62786 440854
rect 63022 440618 63054 440854
rect 62434 423174 63054 440618
rect 62434 422938 62466 423174
rect 62702 422938 62786 423174
rect 63022 422938 63054 423174
rect 62434 422854 63054 422938
rect 62434 422618 62466 422854
rect 62702 422618 62786 422854
rect 63022 422618 63054 422854
rect 62434 405174 63054 422618
rect 62434 404938 62466 405174
rect 62702 404938 62786 405174
rect 63022 404938 63054 405174
rect 62434 404854 63054 404938
rect 62434 404618 62466 404854
rect 62702 404618 62786 404854
rect 63022 404618 63054 404854
rect 62434 387174 63054 404618
rect 62434 386938 62466 387174
rect 62702 386938 62786 387174
rect 63022 386938 63054 387174
rect 62434 386854 63054 386938
rect 62434 386618 62466 386854
rect 62702 386618 62786 386854
rect 63022 386618 63054 386854
rect 62434 369174 63054 386618
rect 62434 368938 62466 369174
rect 62702 368938 62786 369174
rect 63022 368938 63054 369174
rect 62434 368854 63054 368938
rect 62434 368618 62466 368854
rect 62702 368618 62786 368854
rect 63022 368618 63054 368854
rect 62434 351174 63054 368618
rect 62434 350938 62466 351174
rect 62702 350938 62786 351174
rect 63022 350938 63054 351174
rect 62434 350854 63054 350938
rect 62434 350618 62466 350854
rect 62702 350618 62786 350854
rect 63022 350618 63054 350854
rect 62434 333174 63054 350618
rect 62434 332938 62466 333174
rect 62702 332938 62786 333174
rect 63022 332938 63054 333174
rect 62434 332854 63054 332938
rect 62434 332618 62466 332854
rect 62702 332618 62786 332854
rect 63022 332618 63054 332854
rect 62434 315174 63054 332618
rect 62434 314938 62466 315174
rect 62702 314938 62786 315174
rect 63022 314938 63054 315174
rect 62434 314854 63054 314938
rect 62434 314618 62466 314854
rect 62702 314618 62786 314854
rect 63022 314618 63054 314854
rect 62434 297174 63054 314618
rect 62434 296938 62466 297174
rect 62702 296938 62786 297174
rect 63022 296938 63054 297174
rect 62434 296854 63054 296938
rect 62434 296618 62466 296854
rect 62702 296618 62786 296854
rect 63022 296618 63054 296854
rect 62434 279174 63054 296618
rect 62434 278938 62466 279174
rect 62702 278938 62786 279174
rect 63022 278938 63054 279174
rect 62434 278854 63054 278938
rect 62434 278618 62466 278854
rect 62702 278618 62786 278854
rect 63022 278618 63054 278854
rect 62434 261174 63054 278618
rect 62434 260938 62466 261174
rect 62702 260938 62786 261174
rect 63022 260938 63054 261174
rect 62434 260854 63054 260938
rect 62434 260618 62466 260854
rect 62702 260618 62786 260854
rect 63022 260618 63054 260854
rect 62434 243174 63054 260618
rect 62434 242938 62466 243174
rect 62702 242938 62786 243174
rect 63022 242938 63054 243174
rect 62434 242854 63054 242938
rect 62434 242618 62466 242854
rect 62702 242618 62786 242854
rect 63022 242618 63054 242854
rect 62434 225174 63054 242618
rect 62434 224938 62466 225174
rect 62702 224938 62786 225174
rect 63022 224938 63054 225174
rect 62434 224854 63054 224938
rect 62434 224618 62466 224854
rect 62702 224618 62786 224854
rect 63022 224618 63054 224854
rect 62434 207174 63054 224618
rect 62434 206938 62466 207174
rect 62702 206938 62786 207174
rect 63022 206938 63054 207174
rect 62434 206854 63054 206938
rect 62434 206618 62466 206854
rect 62702 206618 62786 206854
rect 63022 206618 63054 206854
rect 62434 189174 63054 206618
rect 62434 188938 62466 189174
rect 62702 188938 62786 189174
rect 63022 188938 63054 189174
rect 62434 188854 63054 188938
rect 62434 188618 62466 188854
rect 62702 188618 62786 188854
rect 63022 188618 63054 188854
rect 62434 171174 63054 188618
rect 62434 170938 62466 171174
rect 62702 170938 62786 171174
rect 63022 170938 63054 171174
rect 62434 170854 63054 170938
rect 62434 170618 62466 170854
rect 62702 170618 62786 170854
rect 63022 170618 63054 170854
rect 62434 153174 63054 170618
rect 62434 152938 62466 153174
rect 62702 152938 62786 153174
rect 63022 152938 63054 153174
rect 62434 152854 63054 152938
rect 62434 152618 62466 152854
rect 62702 152618 62786 152854
rect 63022 152618 63054 152854
rect 62434 135174 63054 152618
rect 62434 134938 62466 135174
rect 62702 134938 62786 135174
rect 63022 134938 63054 135174
rect 62434 134854 63054 134938
rect 62434 134618 62466 134854
rect 62702 134618 62786 134854
rect 63022 134618 63054 134854
rect 62434 117174 63054 134618
rect 62434 116938 62466 117174
rect 62702 116938 62786 117174
rect 63022 116938 63054 117174
rect 62434 116854 63054 116938
rect 62434 116618 62466 116854
rect 62702 116618 62786 116854
rect 63022 116618 63054 116854
rect 62434 99174 63054 116618
rect 62434 98938 62466 99174
rect 62702 98938 62786 99174
rect 63022 98938 63054 99174
rect 62434 98854 63054 98938
rect 62434 98618 62466 98854
rect 62702 98618 62786 98854
rect 63022 98618 63054 98854
rect 62434 81174 63054 98618
rect 62434 80938 62466 81174
rect 62702 80938 62786 81174
rect 63022 80938 63054 81174
rect 62434 80854 63054 80938
rect 62434 80618 62466 80854
rect 62702 80618 62786 80854
rect 63022 80618 63054 80854
rect 62434 63174 63054 80618
rect 62434 62938 62466 63174
rect 62702 62938 62786 63174
rect 63022 62938 63054 63174
rect 62434 62854 63054 62938
rect 62434 62618 62466 62854
rect 62702 62618 62786 62854
rect 63022 62618 63054 62854
rect 62434 45174 63054 62618
rect 62434 44938 62466 45174
rect 62702 44938 62786 45174
rect 63022 44938 63054 45174
rect 62434 44854 63054 44938
rect 62434 44618 62466 44854
rect 62702 44618 62786 44854
rect 63022 44618 63054 44854
rect 62434 27174 63054 44618
rect 62434 26938 62466 27174
rect 62702 26938 62786 27174
rect 63022 26938 63054 27174
rect 62434 26854 63054 26938
rect 62434 26618 62466 26854
rect 62702 26618 62786 26854
rect 63022 26618 63054 26854
rect 62434 9174 63054 26618
rect 62434 8938 62466 9174
rect 62702 8938 62786 9174
rect 63022 8938 63054 9174
rect 62434 8854 63054 8938
rect 62434 8618 62466 8854
rect 62702 8618 62786 8854
rect 63022 8618 63054 8854
rect 62434 -1816 63054 8618
rect 62434 -2052 62466 -1816
rect 62702 -2052 62786 -1816
rect 63022 -2052 63054 -1816
rect 62434 -2136 63054 -2052
rect 62434 -2372 62466 -2136
rect 62702 -2372 62786 -2136
rect 63022 -2372 63054 -2136
rect 62434 -4324 63054 -2372
rect 66154 463012 66774 464004
rect 66154 462776 66186 463012
rect 66422 462776 66506 463012
rect 66742 462776 66774 463012
rect 66154 462692 66774 462776
rect 66154 462456 66186 462692
rect 66422 462456 66506 462692
rect 66742 462456 66774 462692
rect 66154 444894 66774 462456
rect 66154 444658 66186 444894
rect 66422 444658 66506 444894
rect 66742 444658 66774 444894
rect 66154 444574 66774 444658
rect 66154 444338 66186 444574
rect 66422 444338 66506 444574
rect 66742 444338 66774 444574
rect 66154 426894 66774 444338
rect 66154 426658 66186 426894
rect 66422 426658 66506 426894
rect 66742 426658 66774 426894
rect 66154 426574 66774 426658
rect 66154 426338 66186 426574
rect 66422 426338 66506 426574
rect 66742 426338 66774 426574
rect 66154 408894 66774 426338
rect 66154 408658 66186 408894
rect 66422 408658 66506 408894
rect 66742 408658 66774 408894
rect 66154 408574 66774 408658
rect 66154 408338 66186 408574
rect 66422 408338 66506 408574
rect 66742 408338 66774 408574
rect 66154 390894 66774 408338
rect 66154 390658 66186 390894
rect 66422 390658 66506 390894
rect 66742 390658 66774 390894
rect 66154 390574 66774 390658
rect 66154 390338 66186 390574
rect 66422 390338 66506 390574
rect 66742 390338 66774 390574
rect 66154 372894 66774 390338
rect 66154 372658 66186 372894
rect 66422 372658 66506 372894
rect 66742 372658 66774 372894
rect 66154 372574 66774 372658
rect 66154 372338 66186 372574
rect 66422 372338 66506 372574
rect 66742 372338 66774 372574
rect 66154 354894 66774 372338
rect 66154 354658 66186 354894
rect 66422 354658 66506 354894
rect 66742 354658 66774 354894
rect 66154 354574 66774 354658
rect 66154 354338 66186 354574
rect 66422 354338 66506 354574
rect 66742 354338 66774 354574
rect 66154 336894 66774 354338
rect 66154 336658 66186 336894
rect 66422 336658 66506 336894
rect 66742 336658 66774 336894
rect 66154 336574 66774 336658
rect 66154 336338 66186 336574
rect 66422 336338 66506 336574
rect 66742 336338 66774 336574
rect 66154 318894 66774 336338
rect 66154 318658 66186 318894
rect 66422 318658 66506 318894
rect 66742 318658 66774 318894
rect 66154 318574 66774 318658
rect 66154 318338 66186 318574
rect 66422 318338 66506 318574
rect 66742 318338 66774 318574
rect 66154 300894 66774 318338
rect 66154 300658 66186 300894
rect 66422 300658 66506 300894
rect 66742 300658 66774 300894
rect 66154 300574 66774 300658
rect 66154 300338 66186 300574
rect 66422 300338 66506 300574
rect 66742 300338 66774 300574
rect 66154 282894 66774 300338
rect 66154 282658 66186 282894
rect 66422 282658 66506 282894
rect 66742 282658 66774 282894
rect 66154 282574 66774 282658
rect 66154 282338 66186 282574
rect 66422 282338 66506 282574
rect 66742 282338 66774 282574
rect 66154 264894 66774 282338
rect 66154 264658 66186 264894
rect 66422 264658 66506 264894
rect 66742 264658 66774 264894
rect 66154 264574 66774 264658
rect 66154 264338 66186 264574
rect 66422 264338 66506 264574
rect 66742 264338 66774 264574
rect 66154 246894 66774 264338
rect 66154 246658 66186 246894
rect 66422 246658 66506 246894
rect 66742 246658 66774 246894
rect 66154 246574 66774 246658
rect 66154 246338 66186 246574
rect 66422 246338 66506 246574
rect 66742 246338 66774 246574
rect 66154 228894 66774 246338
rect 66154 228658 66186 228894
rect 66422 228658 66506 228894
rect 66742 228658 66774 228894
rect 66154 228574 66774 228658
rect 66154 228338 66186 228574
rect 66422 228338 66506 228574
rect 66742 228338 66774 228574
rect 66154 210894 66774 228338
rect 66154 210658 66186 210894
rect 66422 210658 66506 210894
rect 66742 210658 66774 210894
rect 66154 210574 66774 210658
rect 66154 210338 66186 210574
rect 66422 210338 66506 210574
rect 66742 210338 66774 210574
rect 66154 192894 66774 210338
rect 66154 192658 66186 192894
rect 66422 192658 66506 192894
rect 66742 192658 66774 192894
rect 66154 192574 66774 192658
rect 66154 192338 66186 192574
rect 66422 192338 66506 192574
rect 66742 192338 66774 192574
rect 66154 174894 66774 192338
rect 66154 174658 66186 174894
rect 66422 174658 66506 174894
rect 66742 174658 66774 174894
rect 66154 174574 66774 174658
rect 66154 174338 66186 174574
rect 66422 174338 66506 174574
rect 66742 174338 66774 174574
rect 66154 156894 66774 174338
rect 66154 156658 66186 156894
rect 66422 156658 66506 156894
rect 66742 156658 66774 156894
rect 66154 156574 66774 156658
rect 66154 156338 66186 156574
rect 66422 156338 66506 156574
rect 66742 156338 66774 156574
rect 66154 138894 66774 156338
rect 66154 138658 66186 138894
rect 66422 138658 66506 138894
rect 66742 138658 66774 138894
rect 66154 138574 66774 138658
rect 66154 138338 66186 138574
rect 66422 138338 66506 138574
rect 66742 138338 66774 138574
rect 66154 120894 66774 138338
rect 66154 120658 66186 120894
rect 66422 120658 66506 120894
rect 66742 120658 66774 120894
rect 66154 120574 66774 120658
rect 66154 120338 66186 120574
rect 66422 120338 66506 120574
rect 66742 120338 66774 120574
rect 66154 102894 66774 120338
rect 66154 102658 66186 102894
rect 66422 102658 66506 102894
rect 66742 102658 66774 102894
rect 66154 102574 66774 102658
rect 66154 102338 66186 102574
rect 66422 102338 66506 102574
rect 66742 102338 66774 102574
rect 66154 84894 66774 102338
rect 66154 84658 66186 84894
rect 66422 84658 66506 84894
rect 66742 84658 66774 84894
rect 66154 84574 66774 84658
rect 66154 84338 66186 84574
rect 66422 84338 66506 84574
rect 66742 84338 66774 84574
rect 66154 66894 66774 84338
rect 66154 66658 66186 66894
rect 66422 66658 66506 66894
rect 66742 66658 66774 66894
rect 66154 66574 66774 66658
rect 66154 66338 66186 66574
rect 66422 66338 66506 66574
rect 66742 66338 66774 66574
rect 66154 48894 66774 66338
rect 66154 48658 66186 48894
rect 66422 48658 66506 48894
rect 66742 48658 66774 48894
rect 66154 48574 66774 48658
rect 66154 48338 66186 48574
rect 66422 48338 66506 48574
rect 66742 48338 66774 48574
rect 66154 30894 66774 48338
rect 66154 30658 66186 30894
rect 66422 30658 66506 30894
rect 66742 30658 66774 30894
rect 66154 30574 66774 30658
rect 66154 30338 66186 30574
rect 66422 30338 66506 30574
rect 66742 30338 66774 30574
rect 66154 12894 66774 30338
rect 66154 12658 66186 12894
rect 66422 12658 66506 12894
rect 66742 12658 66774 12894
rect 66154 12574 66774 12658
rect 66154 12338 66186 12574
rect 66422 12338 66506 12574
rect 66742 12338 66774 12574
rect 66154 -2776 66774 12338
rect 66154 -3012 66186 -2776
rect 66422 -3012 66506 -2776
rect 66742 -3012 66774 -2776
rect 66154 -3096 66774 -3012
rect 66154 -3332 66186 -3096
rect 66422 -3332 66506 -3096
rect 66742 -3332 66774 -3096
rect 66154 -4324 66774 -3332
rect 69874 463972 70494 464004
rect 69874 463736 69906 463972
rect 70142 463736 70226 463972
rect 70462 463736 70494 463972
rect 69874 463652 70494 463736
rect 69874 463416 69906 463652
rect 70142 463416 70226 463652
rect 70462 463416 70494 463652
rect 69874 448614 70494 463416
rect 69874 448378 69906 448614
rect 70142 448378 70226 448614
rect 70462 448378 70494 448614
rect 69874 448294 70494 448378
rect 69874 448058 69906 448294
rect 70142 448058 70226 448294
rect 70462 448058 70494 448294
rect 69874 430614 70494 448058
rect 69874 430378 69906 430614
rect 70142 430378 70226 430614
rect 70462 430378 70494 430614
rect 69874 430294 70494 430378
rect 69874 430058 69906 430294
rect 70142 430058 70226 430294
rect 70462 430058 70494 430294
rect 69874 412614 70494 430058
rect 69874 412378 69906 412614
rect 70142 412378 70226 412614
rect 70462 412378 70494 412614
rect 69874 412294 70494 412378
rect 69874 412058 69906 412294
rect 70142 412058 70226 412294
rect 70462 412058 70494 412294
rect 69874 394614 70494 412058
rect 69874 394378 69906 394614
rect 70142 394378 70226 394614
rect 70462 394378 70494 394614
rect 69874 394294 70494 394378
rect 69874 394058 69906 394294
rect 70142 394058 70226 394294
rect 70462 394058 70494 394294
rect 69874 376614 70494 394058
rect 69874 376378 69906 376614
rect 70142 376378 70226 376614
rect 70462 376378 70494 376614
rect 69874 376294 70494 376378
rect 69874 376058 69906 376294
rect 70142 376058 70226 376294
rect 70462 376058 70494 376294
rect 69874 358614 70494 376058
rect 69874 358378 69906 358614
rect 70142 358378 70226 358614
rect 70462 358378 70494 358614
rect 69874 358294 70494 358378
rect 69874 358058 69906 358294
rect 70142 358058 70226 358294
rect 70462 358058 70494 358294
rect 69874 340614 70494 358058
rect 69874 340378 69906 340614
rect 70142 340378 70226 340614
rect 70462 340378 70494 340614
rect 69874 340294 70494 340378
rect 69874 340058 69906 340294
rect 70142 340058 70226 340294
rect 70462 340058 70494 340294
rect 69874 322614 70494 340058
rect 69874 322378 69906 322614
rect 70142 322378 70226 322614
rect 70462 322378 70494 322614
rect 69874 322294 70494 322378
rect 69874 322058 69906 322294
rect 70142 322058 70226 322294
rect 70462 322058 70494 322294
rect 69874 304614 70494 322058
rect 69874 304378 69906 304614
rect 70142 304378 70226 304614
rect 70462 304378 70494 304614
rect 69874 304294 70494 304378
rect 69874 304058 69906 304294
rect 70142 304058 70226 304294
rect 70462 304058 70494 304294
rect 69874 286614 70494 304058
rect 69874 286378 69906 286614
rect 70142 286378 70226 286614
rect 70462 286378 70494 286614
rect 69874 286294 70494 286378
rect 69874 286058 69906 286294
rect 70142 286058 70226 286294
rect 70462 286058 70494 286294
rect 69874 268614 70494 286058
rect 69874 268378 69906 268614
rect 70142 268378 70226 268614
rect 70462 268378 70494 268614
rect 69874 268294 70494 268378
rect 69874 268058 69906 268294
rect 70142 268058 70226 268294
rect 70462 268058 70494 268294
rect 69874 250614 70494 268058
rect 69874 250378 69906 250614
rect 70142 250378 70226 250614
rect 70462 250378 70494 250614
rect 69874 250294 70494 250378
rect 69874 250058 69906 250294
rect 70142 250058 70226 250294
rect 70462 250058 70494 250294
rect 69874 232614 70494 250058
rect 69874 232378 69906 232614
rect 70142 232378 70226 232614
rect 70462 232378 70494 232614
rect 69874 232294 70494 232378
rect 69874 232058 69906 232294
rect 70142 232058 70226 232294
rect 70462 232058 70494 232294
rect 69874 214614 70494 232058
rect 69874 214378 69906 214614
rect 70142 214378 70226 214614
rect 70462 214378 70494 214614
rect 69874 214294 70494 214378
rect 69874 214058 69906 214294
rect 70142 214058 70226 214294
rect 70462 214058 70494 214294
rect 69874 196614 70494 214058
rect 69874 196378 69906 196614
rect 70142 196378 70226 196614
rect 70462 196378 70494 196614
rect 69874 196294 70494 196378
rect 69874 196058 69906 196294
rect 70142 196058 70226 196294
rect 70462 196058 70494 196294
rect 69874 178614 70494 196058
rect 69874 178378 69906 178614
rect 70142 178378 70226 178614
rect 70462 178378 70494 178614
rect 69874 178294 70494 178378
rect 69874 178058 69906 178294
rect 70142 178058 70226 178294
rect 70462 178058 70494 178294
rect 69874 160614 70494 178058
rect 69874 160378 69906 160614
rect 70142 160378 70226 160614
rect 70462 160378 70494 160614
rect 69874 160294 70494 160378
rect 69874 160058 69906 160294
rect 70142 160058 70226 160294
rect 70462 160058 70494 160294
rect 69874 142614 70494 160058
rect 69874 142378 69906 142614
rect 70142 142378 70226 142614
rect 70462 142378 70494 142614
rect 69874 142294 70494 142378
rect 69874 142058 69906 142294
rect 70142 142058 70226 142294
rect 70462 142058 70494 142294
rect 69874 124614 70494 142058
rect 69874 124378 69906 124614
rect 70142 124378 70226 124614
rect 70462 124378 70494 124614
rect 69874 124294 70494 124378
rect 69874 124058 69906 124294
rect 70142 124058 70226 124294
rect 70462 124058 70494 124294
rect 69874 106614 70494 124058
rect 69874 106378 69906 106614
rect 70142 106378 70226 106614
rect 70462 106378 70494 106614
rect 69874 106294 70494 106378
rect 69874 106058 69906 106294
rect 70142 106058 70226 106294
rect 70462 106058 70494 106294
rect 69874 88614 70494 106058
rect 69874 88378 69906 88614
rect 70142 88378 70226 88614
rect 70462 88378 70494 88614
rect 69874 88294 70494 88378
rect 69874 88058 69906 88294
rect 70142 88058 70226 88294
rect 70462 88058 70494 88294
rect 69874 70614 70494 88058
rect 69874 70378 69906 70614
rect 70142 70378 70226 70614
rect 70462 70378 70494 70614
rect 69874 70294 70494 70378
rect 69874 70058 69906 70294
rect 70142 70058 70226 70294
rect 70462 70058 70494 70294
rect 69874 52614 70494 70058
rect 69874 52378 69906 52614
rect 70142 52378 70226 52614
rect 70462 52378 70494 52614
rect 69874 52294 70494 52378
rect 69874 52058 69906 52294
rect 70142 52058 70226 52294
rect 70462 52058 70494 52294
rect 69874 34614 70494 52058
rect 69874 34378 69906 34614
rect 70142 34378 70226 34614
rect 70462 34378 70494 34614
rect 69874 34294 70494 34378
rect 69874 34058 69906 34294
rect 70142 34058 70226 34294
rect 70462 34058 70494 34294
rect 69874 16614 70494 34058
rect 69874 16378 69906 16614
rect 70142 16378 70226 16614
rect 70462 16378 70494 16614
rect 69874 16294 70494 16378
rect 69874 16058 69906 16294
rect 70142 16058 70226 16294
rect 70462 16058 70494 16294
rect 69874 -3736 70494 16058
rect 69874 -3972 69906 -3736
rect 70142 -3972 70226 -3736
rect 70462 -3972 70494 -3736
rect 69874 -4056 70494 -3972
rect 69874 -4292 69906 -4056
rect 70142 -4292 70226 -4056
rect 70462 -4292 70494 -4056
rect 69874 -4324 70494 -4292
rect 76714 461092 77334 464004
rect 76714 460856 76746 461092
rect 76982 460856 77066 461092
rect 77302 460856 77334 461092
rect 76714 460772 77334 460856
rect 76714 460536 76746 460772
rect 76982 460536 77066 460772
rect 77302 460536 77334 460772
rect 76714 455454 77334 460536
rect 76714 455218 76746 455454
rect 76982 455218 77066 455454
rect 77302 455218 77334 455454
rect 76714 455134 77334 455218
rect 76714 454898 76746 455134
rect 76982 454898 77066 455134
rect 77302 454898 77334 455134
rect 76714 437454 77334 454898
rect 76714 437218 76746 437454
rect 76982 437218 77066 437454
rect 77302 437218 77334 437454
rect 76714 437134 77334 437218
rect 76714 436898 76746 437134
rect 76982 436898 77066 437134
rect 77302 436898 77334 437134
rect 76714 419454 77334 436898
rect 76714 419218 76746 419454
rect 76982 419218 77066 419454
rect 77302 419218 77334 419454
rect 76714 419134 77334 419218
rect 76714 418898 76746 419134
rect 76982 418898 77066 419134
rect 77302 418898 77334 419134
rect 76714 401454 77334 418898
rect 76714 401218 76746 401454
rect 76982 401218 77066 401454
rect 77302 401218 77334 401454
rect 76714 401134 77334 401218
rect 76714 400898 76746 401134
rect 76982 400898 77066 401134
rect 77302 400898 77334 401134
rect 76714 383454 77334 400898
rect 76714 383218 76746 383454
rect 76982 383218 77066 383454
rect 77302 383218 77334 383454
rect 76714 383134 77334 383218
rect 76714 382898 76746 383134
rect 76982 382898 77066 383134
rect 77302 382898 77334 383134
rect 76714 365454 77334 382898
rect 76714 365218 76746 365454
rect 76982 365218 77066 365454
rect 77302 365218 77334 365454
rect 76714 365134 77334 365218
rect 76714 364898 76746 365134
rect 76982 364898 77066 365134
rect 77302 364898 77334 365134
rect 76714 347454 77334 364898
rect 76714 347218 76746 347454
rect 76982 347218 77066 347454
rect 77302 347218 77334 347454
rect 76714 347134 77334 347218
rect 76714 346898 76746 347134
rect 76982 346898 77066 347134
rect 77302 346898 77334 347134
rect 76714 329454 77334 346898
rect 76714 329218 76746 329454
rect 76982 329218 77066 329454
rect 77302 329218 77334 329454
rect 76714 329134 77334 329218
rect 76714 328898 76746 329134
rect 76982 328898 77066 329134
rect 77302 328898 77334 329134
rect 76714 311454 77334 328898
rect 76714 311218 76746 311454
rect 76982 311218 77066 311454
rect 77302 311218 77334 311454
rect 76714 311134 77334 311218
rect 76714 310898 76746 311134
rect 76982 310898 77066 311134
rect 77302 310898 77334 311134
rect 76714 293454 77334 310898
rect 76714 293218 76746 293454
rect 76982 293218 77066 293454
rect 77302 293218 77334 293454
rect 76714 293134 77334 293218
rect 76714 292898 76746 293134
rect 76982 292898 77066 293134
rect 77302 292898 77334 293134
rect 76714 275454 77334 292898
rect 76714 275218 76746 275454
rect 76982 275218 77066 275454
rect 77302 275218 77334 275454
rect 76714 275134 77334 275218
rect 76714 274898 76746 275134
rect 76982 274898 77066 275134
rect 77302 274898 77334 275134
rect 76714 257454 77334 274898
rect 76714 257218 76746 257454
rect 76982 257218 77066 257454
rect 77302 257218 77334 257454
rect 76714 257134 77334 257218
rect 76714 256898 76746 257134
rect 76982 256898 77066 257134
rect 77302 256898 77334 257134
rect 76714 239454 77334 256898
rect 76714 239218 76746 239454
rect 76982 239218 77066 239454
rect 77302 239218 77334 239454
rect 76714 239134 77334 239218
rect 76714 238898 76746 239134
rect 76982 238898 77066 239134
rect 77302 238898 77334 239134
rect 76714 221454 77334 238898
rect 76714 221218 76746 221454
rect 76982 221218 77066 221454
rect 77302 221218 77334 221454
rect 76714 221134 77334 221218
rect 76714 220898 76746 221134
rect 76982 220898 77066 221134
rect 77302 220898 77334 221134
rect 76714 203454 77334 220898
rect 76714 203218 76746 203454
rect 76982 203218 77066 203454
rect 77302 203218 77334 203454
rect 76714 203134 77334 203218
rect 76714 202898 76746 203134
rect 76982 202898 77066 203134
rect 77302 202898 77334 203134
rect 76714 185454 77334 202898
rect 76714 185218 76746 185454
rect 76982 185218 77066 185454
rect 77302 185218 77334 185454
rect 76714 185134 77334 185218
rect 76714 184898 76746 185134
rect 76982 184898 77066 185134
rect 77302 184898 77334 185134
rect 76714 167454 77334 184898
rect 76714 167218 76746 167454
rect 76982 167218 77066 167454
rect 77302 167218 77334 167454
rect 76714 167134 77334 167218
rect 76714 166898 76746 167134
rect 76982 166898 77066 167134
rect 77302 166898 77334 167134
rect 76714 149454 77334 166898
rect 76714 149218 76746 149454
rect 76982 149218 77066 149454
rect 77302 149218 77334 149454
rect 76714 149134 77334 149218
rect 76714 148898 76746 149134
rect 76982 148898 77066 149134
rect 77302 148898 77334 149134
rect 76714 131454 77334 148898
rect 76714 131218 76746 131454
rect 76982 131218 77066 131454
rect 77302 131218 77334 131454
rect 76714 131134 77334 131218
rect 76714 130898 76746 131134
rect 76982 130898 77066 131134
rect 77302 130898 77334 131134
rect 76714 113454 77334 130898
rect 76714 113218 76746 113454
rect 76982 113218 77066 113454
rect 77302 113218 77334 113454
rect 76714 113134 77334 113218
rect 76714 112898 76746 113134
rect 76982 112898 77066 113134
rect 77302 112898 77334 113134
rect 76714 95454 77334 112898
rect 76714 95218 76746 95454
rect 76982 95218 77066 95454
rect 77302 95218 77334 95454
rect 76714 95134 77334 95218
rect 76714 94898 76746 95134
rect 76982 94898 77066 95134
rect 77302 94898 77334 95134
rect 76714 77454 77334 94898
rect 76714 77218 76746 77454
rect 76982 77218 77066 77454
rect 77302 77218 77334 77454
rect 76714 77134 77334 77218
rect 76714 76898 76746 77134
rect 76982 76898 77066 77134
rect 77302 76898 77334 77134
rect 76714 59454 77334 76898
rect 76714 59218 76746 59454
rect 76982 59218 77066 59454
rect 77302 59218 77334 59454
rect 76714 59134 77334 59218
rect 76714 58898 76746 59134
rect 76982 58898 77066 59134
rect 77302 58898 77334 59134
rect 76714 41454 77334 58898
rect 76714 41218 76746 41454
rect 76982 41218 77066 41454
rect 77302 41218 77334 41454
rect 76714 41134 77334 41218
rect 76714 40898 76746 41134
rect 76982 40898 77066 41134
rect 77302 40898 77334 41134
rect 76714 23454 77334 40898
rect 76714 23218 76746 23454
rect 76982 23218 77066 23454
rect 77302 23218 77334 23454
rect 76714 23134 77334 23218
rect 76714 22898 76746 23134
rect 76982 22898 77066 23134
rect 77302 22898 77334 23134
rect 76714 5454 77334 22898
rect 76714 5218 76746 5454
rect 76982 5218 77066 5454
rect 77302 5218 77334 5454
rect 76714 5134 77334 5218
rect 76714 4898 76746 5134
rect 76982 4898 77066 5134
rect 77302 4898 77334 5134
rect 76714 -856 77334 4898
rect 76714 -1092 76746 -856
rect 76982 -1092 77066 -856
rect 77302 -1092 77334 -856
rect 76714 -1176 77334 -1092
rect 76714 -1412 76746 -1176
rect 76982 -1412 77066 -1176
rect 77302 -1412 77334 -1176
rect 76714 -4324 77334 -1412
rect 80434 462052 81054 464004
rect 80434 461816 80466 462052
rect 80702 461816 80786 462052
rect 81022 461816 81054 462052
rect 80434 461732 81054 461816
rect 80434 461496 80466 461732
rect 80702 461496 80786 461732
rect 81022 461496 81054 461732
rect 80434 441174 81054 461496
rect 80434 440938 80466 441174
rect 80702 440938 80786 441174
rect 81022 440938 81054 441174
rect 80434 440854 81054 440938
rect 80434 440618 80466 440854
rect 80702 440618 80786 440854
rect 81022 440618 81054 440854
rect 80434 423174 81054 440618
rect 80434 422938 80466 423174
rect 80702 422938 80786 423174
rect 81022 422938 81054 423174
rect 80434 422854 81054 422938
rect 80434 422618 80466 422854
rect 80702 422618 80786 422854
rect 81022 422618 81054 422854
rect 80434 405174 81054 422618
rect 80434 404938 80466 405174
rect 80702 404938 80786 405174
rect 81022 404938 81054 405174
rect 80434 404854 81054 404938
rect 80434 404618 80466 404854
rect 80702 404618 80786 404854
rect 81022 404618 81054 404854
rect 80434 387174 81054 404618
rect 80434 386938 80466 387174
rect 80702 386938 80786 387174
rect 81022 386938 81054 387174
rect 80434 386854 81054 386938
rect 80434 386618 80466 386854
rect 80702 386618 80786 386854
rect 81022 386618 81054 386854
rect 80434 369174 81054 386618
rect 80434 368938 80466 369174
rect 80702 368938 80786 369174
rect 81022 368938 81054 369174
rect 80434 368854 81054 368938
rect 80434 368618 80466 368854
rect 80702 368618 80786 368854
rect 81022 368618 81054 368854
rect 80434 351174 81054 368618
rect 80434 350938 80466 351174
rect 80702 350938 80786 351174
rect 81022 350938 81054 351174
rect 80434 350854 81054 350938
rect 80434 350618 80466 350854
rect 80702 350618 80786 350854
rect 81022 350618 81054 350854
rect 80434 333174 81054 350618
rect 80434 332938 80466 333174
rect 80702 332938 80786 333174
rect 81022 332938 81054 333174
rect 80434 332854 81054 332938
rect 80434 332618 80466 332854
rect 80702 332618 80786 332854
rect 81022 332618 81054 332854
rect 80434 315174 81054 332618
rect 80434 314938 80466 315174
rect 80702 314938 80786 315174
rect 81022 314938 81054 315174
rect 80434 314854 81054 314938
rect 80434 314618 80466 314854
rect 80702 314618 80786 314854
rect 81022 314618 81054 314854
rect 80434 297174 81054 314618
rect 80434 296938 80466 297174
rect 80702 296938 80786 297174
rect 81022 296938 81054 297174
rect 80434 296854 81054 296938
rect 80434 296618 80466 296854
rect 80702 296618 80786 296854
rect 81022 296618 81054 296854
rect 80434 279174 81054 296618
rect 80434 278938 80466 279174
rect 80702 278938 80786 279174
rect 81022 278938 81054 279174
rect 80434 278854 81054 278938
rect 80434 278618 80466 278854
rect 80702 278618 80786 278854
rect 81022 278618 81054 278854
rect 80434 261174 81054 278618
rect 80434 260938 80466 261174
rect 80702 260938 80786 261174
rect 81022 260938 81054 261174
rect 80434 260854 81054 260938
rect 80434 260618 80466 260854
rect 80702 260618 80786 260854
rect 81022 260618 81054 260854
rect 80434 243174 81054 260618
rect 80434 242938 80466 243174
rect 80702 242938 80786 243174
rect 81022 242938 81054 243174
rect 80434 242854 81054 242938
rect 80434 242618 80466 242854
rect 80702 242618 80786 242854
rect 81022 242618 81054 242854
rect 80434 225174 81054 242618
rect 80434 224938 80466 225174
rect 80702 224938 80786 225174
rect 81022 224938 81054 225174
rect 80434 224854 81054 224938
rect 80434 224618 80466 224854
rect 80702 224618 80786 224854
rect 81022 224618 81054 224854
rect 80434 207174 81054 224618
rect 80434 206938 80466 207174
rect 80702 206938 80786 207174
rect 81022 206938 81054 207174
rect 80434 206854 81054 206938
rect 80434 206618 80466 206854
rect 80702 206618 80786 206854
rect 81022 206618 81054 206854
rect 80434 189174 81054 206618
rect 80434 188938 80466 189174
rect 80702 188938 80786 189174
rect 81022 188938 81054 189174
rect 80434 188854 81054 188938
rect 80434 188618 80466 188854
rect 80702 188618 80786 188854
rect 81022 188618 81054 188854
rect 80434 171174 81054 188618
rect 80434 170938 80466 171174
rect 80702 170938 80786 171174
rect 81022 170938 81054 171174
rect 80434 170854 81054 170938
rect 80434 170618 80466 170854
rect 80702 170618 80786 170854
rect 81022 170618 81054 170854
rect 80434 153174 81054 170618
rect 80434 152938 80466 153174
rect 80702 152938 80786 153174
rect 81022 152938 81054 153174
rect 80434 152854 81054 152938
rect 80434 152618 80466 152854
rect 80702 152618 80786 152854
rect 81022 152618 81054 152854
rect 80434 135174 81054 152618
rect 80434 134938 80466 135174
rect 80702 134938 80786 135174
rect 81022 134938 81054 135174
rect 80434 134854 81054 134938
rect 80434 134618 80466 134854
rect 80702 134618 80786 134854
rect 81022 134618 81054 134854
rect 80434 117174 81054 134618
rect 80434 116938 80466 117174
rect 80702 116938 80786 117174
rect 81022 116938 81054 117174
rect 80434 116854 81054 116938
rect 80434 116618 80466 116854
rect 80702 116618 80786 116854
rect 81022 116618 81054 116854
rect 80434 99174 81054 116618
rect 80434 98938 80466 99174
rect 80702 98938 80786 99174
rect 81022 98938 81054 99174
rect 80434 98854 81054 98938
rect 80434 98618 80466 98854
rect 80702 98618 80786 98854
rect 81022 98618 81054 98854
rect 80434 81174 81054 98618
rect 80434 80938 80466 81174
rect 80702 80938 80786 81174
rect 81022 80938 81054 81174
rect 80434 80854 81054 80938
rect 80434 80618 80466 80854
rect 80702 80618 80786 80854
rect 81022 80618 81054 80854
rect 80434 63174 81054 80618
rect 80434 62938 80466 63174
rect 80702 62938 80786 63174
rect 81022 62938 81054 63174
rect 80434 62854 81054 62938
rect 80434 62618 80466 62854
rect 80702 62618 80786 62854
rect 81022 62618 81054 62854
rect 80434 45174 81054 62618
rect 80434 44938 80466 45174
rect 80702 44938 80786 45174
rect 81022 44938 81054 45174
rect 80434 44854 81054 44938
rect 80434 44618 80466 44854
rect 80702 44618 80786 44854
rect 81022 44618 81054 44854
rect 80434 27174 81054 44618
rect 80434 26938 80466 27174
rect 80702 26938 80786 27174
rect 81022 26938 81054 27174
rect 80434 26854 81054 26938
rect 80434 26618 80466 26854
rect 80702 26618 80786 26854
rect 81022 26618 81054 26854
rect 80434 9174 81054 26618
rect 80434 8938 80466 9174
rect 80702 8938 80786 9174
rect 81022 8938 81054 9174
rect 80434 8854 81054 8938
rect 80434 8618 80466 8854
rect 80702 8618 80786 8854
rect 81022 8618 81054 8854
rect 80434 -1816 81054 8618
rect 80434 -2052 80466 -1816
rect 80702 -2052 80786 -1816
rect 81022 -2052 81054 -1816
rect 80434 -2136 81054 -2052
rect 80434 -2372 80466 -2136
rect 80702 -2372 80786 -2136
rect 81022 -2372 81054 -2136
rect 80434 -4324 81054 -2372
rect 84154 463012 84774 464004
rect 84154 462776 84186 463012
rect 84422 462776 84506 463012
rect 84742 462776 84774 463012
rect 84154 462692 84774 462776
rect 84154 462456 84186 462692
rect 84422 462456 84506 462692
rect 84742 462456 84774 462692
rect 84154 444894 84774 462456
rect 84154 444658 84186 444894
rect 84422 444658 84506 444894
rect 84742 444658 84774 444894
rect 84154 444574 84774 444658
rect 84154 444338 84186 444574
rect 84422 444338 84506 444574
rect 84742 444338 84774 444574
rect 84154 426894 84774 444338
rect 84154 426658 84186 426894
rect 84422 426658 84506 426894
rect 84742 426658 84774 426894
rect 84154 426574 84774 426658
rect 84154 426338 84186 426574
rect 84422 426338 84506 426574
rect 84742 426338 84774 426574
rect 84154 408894 84774 426338
rect 84154 408658 84186 408894
rect 84422 408658 84506 408894
rect 84742 408658 84774 408894
rect 84154 408574 84774 408658
rect 84154 408338 84186 408574
rect 84422 408338 84506 408574
rect 84742 408338 84774 408574
rect 84154 390894 84774 408338
rect 84154 390658 84186 390894
rect 84422 390658 84506 390894
rect 84742 390658 84774 390894
rect 84154 390574 84774 390658
rect 84154 390338 84186 390574
rect 84422 390338 84506 390574
rect 84742 390338 84774 390574
rect 84154 372894 84774 390338
rect 84154 372658 84186 372894
rect 84422 372658 84506 372894
rect 84742 372658 84774 372894
rect 84154 372574 84774 372658
rect 84154 372338 84186 372574
rect 84422 372338 84506 372574
rect 84742 372338 84774 372574
rect 84154 354894 84774 372338
rect 84154 354658 84186 354894
rect 84422 354658 84506 354894
rect 84742 354658 84774 354894
rect 84154 354574 84774 354658
rect 84154 354338 84186 354574
rect 84422 354338 84506 354574
rect 84742 354338 84774 354574
rect 84154 336894 84774 354338
rect 84154 336658 84186 336894
rect 84422 336658 84506 336894
rect 84742 336658 84774 336894
rect 84154 336574 84774 336658
rect 84154 336338 84186 336574
rect 84422 336338 84506 336574
rect 84742 336338 84774 336574
rect 84154 318894 84774 336338
rect 84154 318658 84186 318894
rect 84422 318658 84506 318894
rect 84742 318658 84774 318894
rect 84154 318574 84774 318658
rect 84154 318338 84186 318574
rect 84422 318338 84506 318574
rect 84742 318338 84774 318574
rect 84154 300894 84774 318338
rect 84154 300658 84186 300894
rect 84422 300658 84506 300894
rect 84742 300658 84774 300894
rect 84154 300574 84774 300658
rect 84154 300338 84186 300574
rect 84422 300338 84506 300574
rect 84742 300338 84774 300574
rect 84154 282894 84774 300338
rect 84154 282658 84186 282894
rect 84422 282658 84506 282894
rect 84742 282658 84774 282894
rect 84154 282574 84774 282658
rect 84154 282338 84186 282574
rect 84422 282338 84506 282574
rect 84742 282338 84774 282574
rect 84154 264894 84774 282338
rect 84154 264658 84186 264894
rect 84422 264658 84506 264894
rect 84742 264658 84774 264894
rect 84154 264574 84774 264658
rect 84154 264338 84186 264574
rect 84422 264338 84506 264574
rect 84742 264338 84774 264574
rect 84154 246894 84774 264338
rect 84154 246658 84186 246894
rect 84422 246658 84506 246894
rect 84742 246658 84774 246894
rect 84154 246574 84774 246658
rect 84154 246338 84186 246574
rect 84422 246338 84506 246574
rect 84742 246338 84774 246574
rect 84154 228894 84774 246338
rect 84154 228658 84186 228894
rect 84422 228658 84506 228894
rect 84742 228658 84774 228894
rect 84154 228574 84774 228658
rect 84154 228338 84186 228574
rect 84422 228338 84506 228574
rect 84742 228338 84774 228574
rect 84154 210894 84774 228338
rect 84154 210658 84186 210894
rect 84422 210658 84506 210894
rect 84742 210658 84774 210894
rect 84154 210574 84774 210658
rect 84154 210338 84186 210574
rect 84422 210338 84506 210574
rect 84742 210338 84774 210574
rect 84154 192894 84774 210338
rect 84154 192658 84186 192894
rect 84422 192658 84506 192894
rect 84742 192658 84774 192894
rect 84154 192574 84774 192658
rect 84154 192338 84186 192574
rect 84422 192338 84506 192574
rect 84742 192338 84774 192574
rect 84154 174894 84774 192338
rect 84154 174658 84186 174894
rect 84422 174658 84506 174894
rect 84742 174658 84774 174894
rect 84154 174574 84774 174658
rect 84154 174338 84186 174574
rect 84422 174338 84506 174574
rect 84742 174338 84774 174574
rect 84154 156894 84774 174338
rect 84154 156658 84186 156894
rect 84422 156658 84506 156894
rect 84742 156658 84774 156894
rect 84154 156574 84774 156658
rect 84154 156338 84186 156574
rect 84422 156338 84506 156574
rect 84742 156338 84774 156574
rect 84154 138894 84774 156338
rect 84154 138658 84186 138894
rect 84422 138658 84506 138894
rect 84742 138658 84774 138894
rect 84154 138574 84774 138658
rect 84154 138338 84186 138574
rect 84422 138338 84506 138574
rect 84742 138338 84774 138574
rect 84154 120894 84774 138338
rect 84154 120658 84186 120894
rect 84422 120658 84506 120894
rect 84742 120658 84774 120894
rect 84154 120574 84774 120658
rect 84154 120338 84186 120574
rect 84422 120338 84506 120574
rect 84742 120338 84774 120574
rect 84154 102894 84774 120338
rect 84154 102658 84186 102894
rect 84422 102658 84506 102894
rect 84742 102658 84774 102894
rect 84154 102574 84774 102658
rect 84154 102338 84186 102574
rect 84422 102338 84506 102574
rect 84742 102338 84774 102574
rect 84154 84894 84774 102338
rect 84154 84658 84186 84894
rect 84422 84658 84506 84894
rect 84742 84658 84774 84894
rect 84154 84574 84774 84658
rect 84154 84338 84186 84574
rect 84422 84338 84506 84574
rect 84742 84338 84774 84574
rect 84154 66894 84774 84338
rect 84154 66658 84186 66894
rect 84422 66658 84506 66894
rect 84742 66658 84774 66894
rect 84154 66574 84774 66658
rect 84154 66338 84186 66574
rect 84422 66338 84506 66574
rect 84742 66338 84774 66574
rect 84154 48894 84774 66338
rect 84154 48658 84186 48894
rect 84422 48658 84506 48894
rect 84742 48658 84774 48894
rect 84154 48574 84774 48658
rect 84154 48338 84186 48574
rect 84422 48338 84506 48574
rect 84742 48338 84774 48574
rect 84154 30894 84774 48338
rect 84154 30658 84186 30894
rect 84422 30658 84506 30894
rect 84742 30658 84774 30894
rect 84154 30574 84774 30658
rect 84154 30338 84186 30574
rect 84422 30338 84506 30574
rect 84742 30338 84774 30574
rect 84154 12894 84774 30338
rect 84154 12658 84186 12894
rect 84422 12658 84506 12894
rect 84742 12658 84774 12894
rect 84154 12574 84774 12658
rect 84154 12338 84186 12574
rect 84422 12338 84506 12574
rect 84742 12338 84774 12574
rect 84154 -2776 84774 12338
rect 84154 -3012 84186 -2776
rect 84422 -3012 84506 -2776
rect 84742 -3012 84774 -2776
rect 84154 -3096 84774 -3012
rect 84154 -3332 84186 -3096
rect 84422 -3332 84506 -3096
rect 84742 -3332 84774 -3096
rect 84154 -4324 84774 -3332
rect 87874 463972 88494 464004
rect 87874 463736 87906 463972
rect 88142 463736 88226 463972
rect 88462 463736 88494 463972
rect 87874 463652 88494 463736
rect 87874 463416 87906 463652
rect 88142 463416 88226 463652
rect 88462 463416 88494 463652
rect 87874 448614 88494 463416
rect 87874 448378 87906 448614
rect 88142 448378 88226 448614
rect 88462 448378 88494 448614
rect 87874 448294 88494 448378
rect 87874 448058 87906 448294
rect 88142 448058 88226 448294
rect 88462 448058 88494 448294
rect 87874 430614 88494 448058
rect 87874 430378 87906 430614
rect 88142 430378 88226 430614
rect 88462 430378 88494 430614
rect 87874 430294 88494 430378
rect 87874 430058 87906 430294
rect 88142 430058 88226 430294
rect 88462 430058 88494 430294
rect 87874 412614 88494 430058
rect 87874 412378 87906 412614
rect 88142 412378 88226 412614
rect 88462 412378 88494 412614
rect 87874 412294 88494 412378
rect 87874 412058 87906 412294
rect 88142 412058 88226 412294
rect 88462 412058 88494 412294
rect 87874 394614 88494 412058
rect 87874 394378 87906 394614
rect 88142 394378 88226 394614
rect 88462 394378 88494 394614
rect 87874 394294 88494 394378
rect 87874 394058 87906 394294
rect 88142 394058 88226 394294
rect 88462 394058 88494 394294
rect 87874 376614 88494 394058
rect 87874 376378 87906 376614
rect 88142 376378 88226 376614
rect 88462 376378 88494 376614
rect 87874 376294 88494 376378
rect 87874 376058 87906 376294
rect 88142 376058 88226 376294
rect 88462 376058 88494 376294
rect 87874 358614 88494 376058
rect 87874 358378 87906 358614
rect 88142 358378 88226 358614
rect 88462 358378 88494 358614
rect 87874 358294 88494 358378
rect 87874 358058 87906 358294
rect 88142 358058 88226 358294
rect 88462 358058 88494 358294
rect 87874 340614 88494 358058
rect 87874 340378 87906 340614
rect 88142 340378 88226 340614
rect 88462 340378 88494 340614
rect 87874 340294 88494 340378
rect 87874 340058 87906 340294
rect 88142 340058 88226 340294
rect 88462 340058 88494 340294
rect 87874 322614 88494 340058
rect 87874 322378 87906 322614
rect 88142 322378 88226 322614
rect 88462 322378 88494 322614
rect 87874 322294 88494 322378
rect 87874 322058 87906 322294
rect 88142 322058 88226 322294
rect 88462 322058 88494 322294
rect 87874 304614 88494 322058
rect 87874 304378 87906 304614
rect 88142 304378 88226 304614
rect 88462 304378 88494 304614
rect 87874 304294 88494 304378
rect 87874 304058 87906 304294
rect 88142 304058 88226 304294
rect 88462 304058 88494 304294
rect 87874 286614 88494 304058
rect 87874 286378 87906 286614
rect 88142 286378 88226 286614
rect 88462 286378 88494 286614
rect 87874 286294 88494 286378
rect 87874 286058 87906 286294
rect 88142 286058 88226 286294
rect 88462 286058 88494 286294
rect 87874 268614 88494 286058
rect 87874 268378 87906 268614
rect 88142 268378 88226 268614
rect 88462 268378 88494 268614
rect 87874 268294 88494 268378
rect 87874 268058 87906 268294
rect 88142 268058 88226 268294
rect 88462 268058 88494 268294
rect 87874 250614 88494 268058
rect 87874 250378 87906 250614
rect 88142 250378 88226 250614
rect 88462 250378 88494 250614
rect 87874 250294 88494 250378
rect 87874 250058 87906 250294
rect 88142 250058 88226 250294
rect 88462 250058 88494 250294
rect 87874 232614 88494 250058
rect 87874 232378 87906 232614
rect 88142 232378 88226 232614
rect 88462 232378 88494 232614
rect 87874 232294 88494 232378
rect 87874 232058 87906 232294
rect 88142 232058 88226 232294
rect 88462 232058 88494 232294
rect 87874 214614 88494 232058
rect 87874 214378 87906 214614
rect 88142 214378 88226 214614
rect 88462 214378 88494 214614
rect 87874 214294 88494 214378
rect 87874 214058 87906 214294
rect 88142 214058 88226 214294
rect 88462 214058 88494 214294
rect 87874 196614 88494 214058
rect 87874 196378 87906 196614
rect 88142 196378 88226 196614
rect 88462 196378 88494 196614
rect 87874 196294 88494 196378
rect 87874 196058 87906 196294
rect 88142 196058 88226 196294
rect 88462 196058 88494 196294
rect 87874 178614 88494 196058
rect 87874 178378 87906 178614
rect 88142 178378 88226 178614
rect 88462 178378 88494 178614
rect 87874 178294 88494 178378
rect 87874 178058 87906 178294
rect 88142 178058 88226 178294
rect 88462 178058 88494 178294
rect 87874 160614 88494 178058
rect 87874 160378 87906 160614
rect 88142 160378 88226 160614
rect 88462 160378 88494 160614
rect 87874 160294 88494 160378
rect 87874 160058 87906 160294
rect 88142 160058 88226 160294
rect 88462 160058 88494 160294
rect 87874 142614 88494 160058
rect 87874 142378 87906 142614
rect 88142 142378 88226 142614
rect 88462 142378 88494 142614
rect 87874 142294 88494 142378
rect 87874 142058 87906 142294
rect 88142 142058 88226 142294
rect 88462 142058 88494 142294
rect 87874 124614 88494 142058
rect 87874 124378 87906 124614
rect 88142 124378 88226 124614
rect 88462 124378 88494 124614
rect 87874 124294 88494 124378
rect 87874 124058 87906 124294
rect 88142 124058 88226 124294
rect 88462 124058 88494 124294
rect 87874 106614 88494 124058
rect 87874 106378 87906 106614
rect 88142 106378 88226 106614
rect 88462 106378 88494 106614
rect 87874 106294 88494 106378
rect 87874 106058 87906 106294
rect 88142 106058 88226 106294
rect 88462 106058 88494 106294
rect 87874 88614 88494 106058
rect 87874 88378 87906 88614
rect 88142 88378 88226 88614
rect 88462 88378 88494 88614
rect 87874 88294 88494 88378
rect 87874 88058 87906 88294
rect 88142 88058 88226 88294
rect 88462 88058 88494 88294
rect 87874 70614 88494 88058
rect 87874 70378 87906 70614
rect 88142 70378 88226 70614
rect 88462 70378 88494 70614
rect 87874 70294 88494 70378
rect 87874 70058 87906 70294
rect 88142 70058 88226 70294
rect 88462 70058 88494 70294
rect 87874 52614 88494 70058
rect 94714 461092 95334 464004
rect 94714 460856 94746 461092
rect 94982 460856 95066 461092
rect 95302 460856 95334 461092
rect 94714 460772 95334 460856
rect 94714 460536 94746 460772
rect 94982 460536 95066 460772
rect 95302 460536 95334 460772
rect 94714 455454 95334 460536
rect 94714 455218 94746 455454
rect 94982 455218 95066 455454
rect 95302 455218 95334 455454
rect 94714 455134 95334 455218
rect 94714 454898 94746 455134
rect 94982 454898 95066 455134
rect 95302 454898 95334 455134
rect 94714 437454 95334 454898
rect 94714 437218 94746 437454
rect 94982 437218 95066 437454
rect 95302 437218 95334 437454
rect 94714 437134 95334 437218
rect 94714 436898 94746 437134
rect 94982 436898 95066 437134
rect 95302 436898 95334 437134
rect 94714 419454 95334 436898
rect 94714 419218 94746 419454
rect 94982 419218 95066 419454
rect 95302 419218 95334 419454
rect 94714 419134 95334 419218
rect 94714 418898 94746 419134
rect 94982 418898 95066 419134
rect 95302 418898 95334 419134
rect 94714 401454 95334 418898
rect 94714 401218 94746 401454
rect 94982 401218 95066 401454
rect 95302 401218 95334 401454
rect 94714 401134 95334 401218
rect 94714 400898 94746 401134
rect 94982 400898 95066 401134
rect 95302 400898 95334 401134
rect 94714 383454 95334 400898
rect 94714 383218 94746 383454
rect 94982 383218 95066 383454
rect 95302 383218 95334 383454
rect 94714 383134 95334 383218
rect 94714 382898 94746 383134
rect 94982 382898 95066 383134
rect 95302 382898 95334 383134
rect 94714 365454 95334 382898
rect 94714 365218 94746 365454
rect 94982 365218 95066 365454
rect 95302 365218 95334 365454
rect 94714 365134 95334 365218
rect 94714 364898 94746 365134
rect 94982 364898 95066 365134
rect 95302 364898 95334 365134
rect 94714 347454 95334 364898
rect 94714 347218 94746 347454
rect 94982 347218 95066 347454
rect 95302 347218 95334 347454
rect 94714 347134 95334 347218
rect 94714 346898 94746 347134
rect 94982 346898 95066 347134
rect 95302 346898 95334 347134
rect 94714 329454 95334 346898
rect 94714 329218 94746 329454
rect 94982 329218 95066 329454
rect 95302 329218 95334 329454
rect 94714 329134 95334 329218
rect 94714 328898 94746 329134
rect 94982 328898 95066 329134
rect 95302 328898 95334 329134
rect 94714 311454 95334 328898
rect 94714 311218 94746 311454
rect 94982 311218 95066 311454
rect 95302 311218 95334 311454
rect 94714 311134 95334 311218
rect 94714 310898 94746 311134
rect 94982 310898 95066 311134
rect 95302 310898 95334 311134
rect 94714 293454 95334 310898
rect 94714 293218 94746 293454
rect 94982 293218 95066 293454
rect 95302 293218 95334 293454
rect 94714 293134 95334 293218
rect 94714 292898 94746 293134
rect 94982 292898 95066 293134
rect 95302 292898 95334 293134
rect 94714 275454 95334 292898
rect 94714 275218 94746 275454
rect 94982 275218 95066 275454
rect 95302 275218 95334 275454
rect 94714 275134 95334 275218
rect 94714 274898 94746 275134
rect 94982 274898 95066 275134
rect 95302 274898 95334 275134
rect 94714 257454 95334 274898
rect 94714 257218 94746 257454
rect 94982 257218 95066 257454
rect 95302 257218 95334 257454
rect 94714 257134 95334 257218
rect 94714 256898 94746 257134
rect 94982 256898 95066 257134
rect 95302 256898 95334 257134
rect 94714 239454 95334 256898
rect 94714 239218 94746 239454
rect 94982 239218 95066 239454
rect 95302 239218 95334 239454
rect 94714 239134 95334 239218
rect 94714 238898 94746 239134
rect 94982 238898 95066 239134
rect 95302 238898 95334 239134
rect 94714 221454 95334 238898
rect 94714 221218 94746 221454
rect 94982 221218 95066 221454
rect 95302 221218 95334 221454
rect 94714 221134 95334 221218
rect 94714 220898 94746 221134
rect 94982 220898 95066 221134
rect 95302 220898 95334 221134
rect 94714 203454 95334 220898
rect 94714 203218 94746 203454
rect 94982 203218 95066 203454
rect 95302 203218 95334 203454
rect 94714 203134 95334 203218
rect 94714 202898 94746 203134
rect 94982 202898 95066 203134
rect 95302 202898 95334 203134
rect 94714 185454 95334 202898
rect 94714 185218 94746 185454
rect 94982 185218 95066 185454
rect 95302 185218 95334 185454
rect 94714 185134 95334 185218
rect 94714 184898 94746 185134
rect 94982 184898 95066 185134
rect 95302 184898 95334 185134
rect 94714 167454 95334 184898
rect 94714 167218 94746 167454
rect 94982 167218 95066 167454
rect 95302 167218 95334 167454
rect 94714 167134 95334 167218
rect 94714 166898 94746 167134
rect 94982 166898 95066 167134
rect 95302 166898 95334 167134
rect 94714 149454 95334 166898
rect 94714 149218 94746 149454
rect 94982 149218 95066 149454
rect 95302 149218 95334 149454
rect 94714 149134 95334 149218
rect 94714 148898 94746 149134
rect 94982 148898 95066 149134
rect 95302 148898 95334 149134
rect 94714 131454 95334 148898
rect 94714 131218 94746 131454
rect 94982 131218 95066 131454
rect 95302 131218 95334 131454
rect 94714 131134 95334 131218
rect 94714 130898 94746 131134
rect 94982 130898 95066 131134
rect 95302 130898 95334 131134
rect 94714 113454 95334 130898
rect 94714 113218 94746 113454
rect 94982 113218 95066 113454
rect 95302 113218 95334 113454
rect 94714 113134 95334 113218
rect 94714 112898 94746 113134
rect 94982 112898 95066 113134
rect 95302 112898 95334 113134
rect 94714 95454 95334 112898
rect 94714 95218 94746 95454
rect 94982 95218 95066 95454
rect 95302 95218 95334 95454
rect 94714 95134 95334 95218
rect 94714 94898 94746 95134
rect 94982 94898 95066 95134
rect 95302 94898 95334 95134
rect 94714 77454 95334 94898
rect 94714 77218 94746 77454
rect 94982 77218 95066 77454
rect 95302 77218 95334 77454
rect 94714 77134 95334 77218
rect 94714 76898 94746 77134
rect 94982 76898 95066 77134
rect 95302 76898 95334 77134
rect 94714 59724 95334 76898
rect 98434 462052 99054 464004
rect 98434 461816 98466 462052
rect 98702 461816 98786 462052
rect 99022 461816 99054 462052
rect 98434 461732 99054 461816
rect 98434 461496 98466 461732
rect 98702 461496 98786 461732
rect 99022 461496 99054 461732
rect 98434 441174 99054 461496
rect 98434 440938 98466 441174
rect 98702 440938 98786 441174
rect 99022 440938 99054 441174
rect 98434 440854 99054 440938
rect 98434 440618 98466 440854
rect 98702 440618 98786 440854
rect 99022 440618 99054 440854
rect 98434 423174 99054 440618
rect 98434 422938 98466 423174
rect 98702 422938 98786 423174
rect 99022 422938 99054 423174
rect 98434 422854 99054 422938
rect 98434 422618 98466 422854
rect 98702 422618 98786 422854
rect 99022 422618 99054 422854
rect 98434 405174 99054 422618
rect 98434 404938 98466 405174
rect 98702 404938 98786 405174
rect 99022 404938 99054 405174
rect 98434 404854 99054 404938
rect 98434 404618 98466 404854
rect 98702 404618 98786 404854
rect 99022 404618 99054 404854
rect 98434 387174 99054 404618
rect 98434 386938 98466 387174
rect 98702 386938 98786 387174
rect 99022 386938 99054 387174
rect 98434 386854 99054 386938
rect 98434 386618 98466 386854
rect 98702 386618 98786 386854
rect 99022 386618 99054 386854
rect 98434 369174 99054 386618
rect 98434 368938 98466 369174
rect 98702 368938 98786 369174
rect 99022 368938 99054 369174
rect 98434 368854 99054 368938
rect 98434 368618 98466 368854
rect 98702 368618 98786 368854
rect 99022 368618 99054 368854
rect 98434 351174 99054 368618
rect 98434 350938 98466 351174
rect 98702 350938 98786 351174
rect 99022 350938 99054 351174
rect 98434 350854 99054 350938
rect 98434 350618 98466 350854
rect 98702 350618 98786 350854
rect 99022 350618 99054 350854
rect 98434 333174 99054 350618
rect 98434 332938 98466 333174
rect 98702 332938 98786 333174
rect 99022 332938 99054 333174
rect 98434 332854 99054 332938
rect 98434 332618 98466 332854
rect 98702 332618 98786 332854
rect 99022 332618 99054 332854
rect 98434 315174 99054 332618
rect 98434 314938 98466 315174
rect 98702 314938 98786 315174
rect 99022 314938 99054 315174
rect 98434 314854 99054 314938
rect 98434 314618 98466 314854
rect 98702 314618 98786 314854
rect 99022 314618 99054 314854
rect 98434 297174 99054 314618
rect 98434 296938 98466 297174
rect 98702 296938 98786 297174
rect 99022 296938 99054 297174
rect 98434 296854 99054 296938
rect 98434 296618 98466 296854
rect 98702 296618 98786 296854
rect 99022 296618 99054 296854
rect 98434 279174 99054 296618
rect 98434 278938 98466 279174
rect 98702 278938 98786 279174
rect 99022 278938 99054 279174
rect 98434 278854 99054 278938
rect 98434 278618 98466 278854
rect 98702 278618 98786 278854
rect 99022 278618 99054 278854
rect 98434 261174 99054 278618
rect 98434 260938 98466 261174
rect 98702 260938 98786 261174
rect 99022 260938 99054 261174
rect 98434 260854 99054 260938
rect 98434 260618 98466 260854
rect 98702 260618 98786 260854
rect 99022 260618 99054 260854
rect 98434 243174 99054 260618
rect 98434 242938 98466 243174
rect 98702 242938 98786 243174
rect 99022 242938 99054 243174
rect 98434 242854 99054 242938
rect 98434 242618 98466 242854
rect 98702 242618 98786 242854
rect 99022 242618 99054 242854
rect 98434 225174 99054 242618
rect 98434 224938 98466 225174
rect 98702 224938 98786 225174
rect 99022 224938 99054 225174
rect 98434 224854 99054 224938
rect 98434 224618 98466 224854
rect 98702 224618 98786 224854
rect 99022 224618 99054 224854
rect 98434 207174 99054 224618
rect 98434 206938 98466 207174
rect 98702 206938 98786 207174
rect 99022 206938 99054 207174
rect 98434 206854 99054 206938
rect 98434 206618 98466 206854
rect 98702 206618 98786 206854
rect 99022 206618 99054 206854
rect 98434 189174 99054 206618
rect 98434 188938 98466 189174
rect 98702 188938 98786 189174
rect 99022 188938 99054 189174
rect 98434 188854 99054 188938
rect 98434 188618 98466 188854
rect 98702 188618 98786 188854
rect 99022 188618 99054 188854
rect 98434 171174 99054 188618
rect 98434 170938 98466 171174
rect 98702 170938 98786 171174
rect 99022 170938 99054 171174
rect 98434 170854 99054 170938
rect 98434 170618 98466 170854
rect 98702 170618 98786 170854
rect 99022 170618 99054 170854
rect 98434 153174 99054 170618
rect 98434 152938 98466 153174
rect 98702 152938 98786 153174
rect 99022 152938 99054 153174
rect 98434 152854 99054 152938
rect 98434 152618 98466 152854
rect 98702 152618 98786 152854
rect 99022 152618 99054 152854
rect 98434 135174 99054 152618
rect 98434 134938 98466 135174
rect 98702 134938 98786 135174
rect 99022 134938 99054 135174
rect 98434 134854 99054 134938
rect 98434 134618 98466 134854
rect 98702 134618 98786 134854
rect 99022 134618 99054 134854
rect 98434 117174 99054 134618
rect 98434 116938 98466 117174
rect 98702 116938 98786 117174
rect 99022 116938 99054 117174
rect 98434 116854 99054 116938
rect 98434 116618 98466 116854
rect 98702 116618 98786 116854
rect 99022 116618 99054 116854
rect 98434 99174 99054 116618
rect 98434 98938 98466 99174
rect 98702 98938 98786 99174
rect 99022 98938 99054 99174
rect 98434 98854 99054 98938
rect 98434 98618 98466 98854
rect 98702 98618 98786 98854
rect 99022 98618 99054 98854
rect 98434 81174 99054 98618
rect 98434 80938 98466 81174
rect 98702 80938 98786 81174
rect 99022 80938 99054 81174
rect 98434 80854 99054 80938
rect 98434 80618 98466 80854
rect 98702 80618 98786 80854
rect 99022 80618 99054 80854
rect 98434 63174 99054 80618
rect 98434 62938 98466 63174
rect 98702 62938 98786 63174
rect 99022 62938 99054 63174
rect 98434 62854 99054 62938
rect 98434 62618 98466 62854
rect 98702 62618 98786 62854
rect 99022 62618 99054 62854
rect 98434 58629 99054 62618
rect 102154 463012 102774 464004
rect 102154 462776 102186 463012
rect 102422 462776 102506 463012
rect 102742 462776 102774 463012
rect 102154 462692 102774 462776
rect 102154 462456 102186 462692
rect 102422 462456 102506 462692
rect 102742 462456 102774 462692
rect 102154 444894 102774 462456
rect 102154 444658 102186 444894
rect 102422 444658 102506 444894
rect 102742 444658 102774 444894
rect 102154 444574 102774 444658
rect 102154 444338 102186 444574
rect 102422 444338 102506 444574
rect 102742 444338 102774 444574
rect 102154 426894 102774 444338
rect 102154 426658 102186 426894
rect 102422 426658 102506 426894
rect 102742 426658 102774 426894
rect 102154 426574 102774 426658
rect 102154 426338 102186 426574
rect 102422 426338 102506 426574
rect 102742 426338 102774 426574
rect 102154 408894 102774 426338
rect 102154 408658 102186 408894
rect 102422 408658 102506 408894
rect 102742 408658 102774 408894
rect 102154 408574 102774 408658
rect 102154 408338 102186 408574
rect 102422 408338 102506 408574
rect 102742 408338 102774 408574
rect 102154 390894 102774 408338
rect 102154 390658 102186 390894
rect 102422 390658 102506 390894
rect 102742 390658 102774 390894
rect 102154 390574 102774 390658
rect 102154 390338 102186 390574
rect 102422 390338 102506 390574
rect 102742 390338 102774 390574
rect 102154 372894 102774 390338
rect 102154 372658 102186 372894
rect 102422 372658 102506 372894
rect 102742 372658 102774 372894
rect 102154 372574 102774 372658
rect 102154 372338 102186 372574
rect 102422 372338 102506 372574
rect 102742 372338 102774 372574
rect 102154 354894 102774 372338
rect 102154 354658 102186 354894
rect 102422 354658 102506 354894
rect 102742 354658 102774 354894
rect 102154 354574 102774 354658
rect 102154 354338 102186 354574
rect 102422 354338 102506 354574
rect 102742 354338 102774 354574
rect 102154 336894 102774 354338
rect 102154 336658 102186 336894
rect 102422 336658 102506 336894
rect 102742 336658 102774 336894
rect 102154 336574 102774 336658
rect 102154 336338 102186 336574
rect 102422 336338 102506 336574
rect 102742 336338 102774 336574
rect 102154 318894 102774 336338
rect 102154 318658 102186 318894
rect 102422 318658 102506 318894
rect 102742 318658 102774 318894
rect 102154 318574 102774 318658
rect 102154 318338 102186 318574
rect 102422 318338 102506 318574
rect 102742 318338 102774 318574
rect 102154 300894 102774 318338
rect 102154 300658 102186 300894
rect 102422 300658 102506 300894
rect 102742 300658 102774 300894
rect 102154 300574 102774 300658
rect 102154 300338 102186 300574
rect 102422 300338 102506 300574
rect 102742 300338 102774 300574
rect 102154 282894 102774 300338
rect 102154 282658 102186 282894
rect 102422 282658 102506 282894
rect 102742 282658 102774 282894
rect 102154 282574 102774 282658
rect 102154 282338 102186 282574
rect 102422 282338 102506 282574
rect 102742 282338 102774 282574
rect 102154 264894 102774 282338
rect 102154 264658 102186 264894
rect 102422 264658 102506 264894
rect 102742 264658 102774 264894
rect 102154 264574 102774 264658
rect 102154 264338 102186 264574
rect 102422 264338 102506 264574
rect 102742 264338 102774 264574
rect 102154 246894 102774 264338
rect 102154 246658 102186 246894
rect 102422 246658 102506 246894
rect 102742 246658 102774 246894
rect 102154 246574 102774 246658
rect 102154 246338 102186 246574
rect 102422 246338 102506 246574
rect 102742 246338 102774 246574
rect 102154 228894 102774 246338
rect 102154 228658 102186 228894
rect 102422 228658 102506 228894
rect 102742 228658 102774 228894
rect 102154 228574 102774 228658
rect 102154 228338 102186 228574
rect 102422 228338 102506 228574
rect 102742 228338 102774 228574
rect 102154 210894 102774 228338
rect 102154 210658 102186 210894
rect 102422 210658 102506 210894
rect 102742 210658 102774 210894
rect 102154 210574 102774 210658
rect 102154 210338 102186 210574
rect 102422 210338 102506 210574
rect 102742 210338 102774 210574
rect 102154 192894 102774 210338
rect 102154 192658 102186 192894
rect 102422 192658 102506 192894
rect 102742 192658 102774 192894
rect 102154 192574 102774 192658
rect 102154 192338 102186 192574
rect 102422 192338 102506 192574
rect 102742 192338 102774 192574
rect 102154 174894 102774 192338
rect 102154 174658 102186 174894
rect 102422 174658 102506 174894
rect 102742 174658 102774 174894
rect 102154 174574 102774 174658
rect 102154 174338 102186 174574
rect 102422 174338 102506 174574
rect 102742 174338 102774 174574
rect 102154 156894 102774 174338
rect 102154 156658 102186 156894
rect 102422 156658 102506 156894
rect 102742 156658 102774 156894
rect 102154 156574 102774 156658
rect 102154 156338 102186 156574
rect 102422 156338 102506 156574
rect 102742 156338 102774 156574
rect 102154 138894 102774 156338
rect 102154 138658 102186 138894
rect 102422 138658 102506 138894
rect 102742 138658 102774 138894
rect 102154 138574 102774 138658
rect 102154 138338 102186 138574
rect 102422 138338 102506 138574
rect 102742 138338 102774 138574
rect 102154 120894 102774 138338
rect 102154 120658 102186 120894
rect 102422 120658 102506 120894
rect 102742 120658 102774 120894
rect 102154 120574 102774 120658
rect 102154 120338 102186 120574
rect 102422 120338 102506 120574
rect 102742 120338 102774 120574
rect 102154 102894 102774 120338
rect 102154 102658 102186 102894
rect 102422 102658 102506 102894
rect 102742 102658 102774 102894
rect 102154 102574 102774 102658
rect 102154 102338 102186 102574
rect 102422 102338 102506 102574
rect 102742 102338 102774 102574
rect 102154 84894 102774 102338
rect 102154 84658 102186 84894
rect 102422 84658 102506 84894
rect 102742 84658 102774 84894
rect 102154 84574 102774 84658
rect 102154 84338 102186 84574
rect 102422 84338 102506 84574
rect 102742 84338 102774 84574
rect 102154 66894 102774 84338
rect 102154 66658 102186 66894
rect 102422 66658 102506 66894
rect 102742 66658 102774 66894
rect 102154 66574 102774 66658
rect 102154 66338 102186 66574
rect 102422 66338 102506 66574
rect 102742 66338 102774 66574
rect 102154 58629 102774 66338
rect 105874 463972 106494 464004
rect 105874 463736 105906 463972
rect 106142 463736 106226 463972
rect 106462 463736 106494 463972
rect 105874 463652 106494 463736
rect 105874 463416 105906 463652
rect 106142 463416 106226 463652
rect 106462 463416 106494 463652
rect 105874 448614 106494 463416
rect 105874 448378 105906 448614
rect 106142 448378 106226 448614
rect 106462 448378 106494 448614
rect 105874 448294 106494 448378
rect 105874 448058 105906 448294
rect 106142 448058 106226 448294
rect 106462 448058 106494 448294
rect 105874 430614 106494 448058
rect 105874 430378 105906 430614
rect 106142 430378 106226 430614
rect 106462 430378 106494 430614
rect 105874 430294 106494 430378
rect 105874 430058 105906 430294
rect 106142 430058 106226 430294
rect 106462 430058 106494 430294
rect 105874 412614 106494 430058
rect 105874 412378 105906 412614
rect 106142 412378 106226 412614
rect 106462 412378 106494 412614
rect 105874 412294 106494 412378
rect 105874 412058 105906 412294
rect 106142 412058 106226 412294
rect 106462 412058 106494 412294
rect 105874 394614 106494 412058
rect 105874 394378 105906 394614
rect 106142 394378 106226 394614
rect 106462 394378 106494 394614
rect 105874 394294 106494 394378
rect 105874 394058 105906 394294
rect 106142 394058 106226 394294
rect 106462 394058 106494 394294
rect 105874 376614 106494 394058
rect 105874 376378 105906 376614
rect 106142 376378 106226 376614
rect 106462 376378 106494 376614
rect 105874 376294 106494 376378
rect 105874 376058 105906 376294
rect 106142 376058 106226 376294
rect 106462 376058 106494 376294
rect 105874 358614 106494 376058
rect 105874 358378 105906 358614
rect 106142 358378 106226 358614
rect 106462 358378 106494 358614
rect 105874 358294 106494 358378
rect 105874 358058 105906 358294
rect 106142 358058 106226 358294
rect 106462 358058 106494 358294
rect 105874 340614 106494 358058
rect 105874 340378 105906 340614
rect 106142 340378 106226 340614
rect 106462 340378 106494 340614
rect 105874 340294 106494 340378
rect 105874 340058 105906 340294
rect 106142 340058 106226 340294
rect 106462 340058 106494 340294
rect 105874 322614 106494 340058
rect 105874 322378 105906 322614
rect 106142 322378 106226 322614
rect 106462 322378 106494 322614
rect 105874 322294 106494 322378
rect 105874 322058 105906 322294
rect 106142 322058 106226 322294
rect 106462 322058 106494 322294
rect 105874 304614 106494 322058
rect 105874 304378 105906 304614
rect 106142 304378 106226 304614
rect 106462 304378 106494 304614
rect 105874 304294 106494 304378
rect 105874 304058 105906 304294
rect 106142 304058 106226 304294
rect 106462 304058 106494 304294
rect 105874 286614 106494 304058
rect 105874 286378 105906 286614
rect 106142 286378 106226 286614
rect 106462 286378 106494 286614
rect 105874 286294 106494 286378
rect 105874 286058 105906 286294
rect 106142 286058 106226 286294
rect 106462 286058 106494 286294
rect 105874 268614 106494 286058
rect 105874 268378 105906 268614
rect 106142 268378 106226 268614
rect 106462 268378 106494 268614
rect 105874 268294 106494 268378
rect 105874 268058 105906 268294
rect 106142 268058 106226 268294
rect 106462 268058 106494 268294
rect 105874 250614 106494 268058
rect 105874 250378 105906 250614
rect 106142 250378 106226 250614
rect 106462 250378 106494 250614
rect 105874 250294 106494 250378
rect 105874 250058 105906 250294
rect 106142 250058 106226 250294
rect 106462 250058 106494 250294
rect 105874 232614 106494 250058
rect 105874 232378 105906 232614
rect 106142 232378 106226 232614
rect 106462 232378 106494 232614
rect 105874 232294 106494 232378
rect 105874 232058 105906 232294
rect 106142 232058 106226 232294
rect 106462 232058 106494 232294
rect 105874 214614 106494 232058
rect 105874 214378 105906 214614
rect 106142 214378 106226 214614
rect 106462 214378 106494 214614
rect 105874 214294 106494 214378
rect 105874 214058 105906 214294
rect 106142 214058 106226 214294
rect 106462 214058 106494 214294
rect 105874 196614 106494 214058
rect 105874 196378 105906 196614
rect 106142 196378 106226 196614
rect 106462 196378 106494 196614
rect 105874 196294 106494 196378
rect 105874 196058 105906 196294
rect 106142 196058 106226 196294
rect 106462 196058 106494 196294
rect 105874 178614 106494 196058
rect 105874 178378 105906 178614
rect 106142 178378 106226 178614
rect 106462 178378 106494 178614
rect 105874 178294 106494 178378
rect 105874 178058 105906 178294
rect 106142 178058 106226 178294
rect 106462 178058 106494 178294
rect 105874 160614 106494 178058
rect 105874 160378 105906 160614
rect 106142 160378 106226 160614
rect 106462 160378 106494 160614
rect 105874 160294 106494 160378
rect 105874 160058 105906 160294
rect 106142 160058 106226 160294
rect 106462 160058 106494 160294
rect 105874 142614 106494 160058
rect 105874 142378 105906 142614
rect 106142 142378 106226 142614
rect 106462 142378 106494 142614
rect 105874 142294 106494 142378
rect 105874 142058 105906 142294
rect 106142 142058 106226 142294
rect 106462 142058 106494 142294
rect 105874 124614 106494 142058
rect 105874 124378 105906 124614
rect 106142 124378 106226 124614
rect 106462 124378 106494 124614
rect 105874 124294 106494 124378
rect 105874 124058 105906 124294
rect 106142 124058 106226 124294
rect 106462 124058 106494 124294
rect 105874 106614 106494 124058
rect 105874 106378 105906 106614
rect 106142 106378 106226 106614
rect 106462 106378 106494 106614
rect 105874 106294 106494 106378
rect 105874 106058 105906 106294
rect 106142 106058 106226 106294
rect 106462 106058 106494 106294
rect 105874 88614 106494 106058
rect 105874 88378 105906 88614
rect 106142 88378 106226 88614
rect 106462 88378 106494 88614
rect 105874 88294 106494 88378
rect 105874 88058 105906 88294
rect 106142 88058 106226 88294
rect 106462 88058 106494 88294
rect 105874 70614 106494 88058
rect 105874 70378 105906 70614
rect 106142 70378 106226 70614
rect 106462 70378 106494 70614
rect 105874 70294 106494 70378
rect 105874 70058 105906 70294
rect 106142 70058 106226 70294
rect 106462 70058 106494 70294
rect 105874 58629 106494 70058
rect 112714 461092 113334 464004
rect 112714 460856 112746 461092
rect 112982 460856 113066 461092
rect 113302 460856 113334 461092
rect 112714 460772 113334 460856
rect 112714 460536 112746 460772
rect 112982 460536 113066 460772
rect 113302 460536 113334 460772
rect 112714 455454 113334 460536
rect 112714 455218 112746 455454
rect 112982 455218 113066 455454
rect 113302 455218 113334 455454
rect 112714 455134 113334 455218
rect 112714 454898 112746 455134
rect 112982 454898 113066 455134
rect 113302 454898 113334 455134
rect 112714 437454 113334 454898
rect 112714 437218 112746 437454
rect 112982 437218 113066 437454
rect 113302 437218 113334 437454
rect 112714 437134 113334 437218
rect 112714 436898 112746 437134
rect 112982 436898 113066 437134
rect 113302 436898 113334 437134
rect 112714 419454 113334 436898
rect 112714 419218 112746 419454
rect 112982 419218 113066 419454
rect 113302 419218 113334 419454
rect 112714 419134 113334 419218
rect 112714 418898 112746 419134
rect 112982 418898 113066 419134
rect 113302 418898 113334 419134
rect 112714 401454 113334 418898
rect 112714 401218 112746 401454
rect 112982 401218 113066 401454
rect 113302 401218 113334 401454
rect 112714 401134 113334 401218
rect 112714 400898 112746 401134
rect 112982 400898 113066 401134
rect 113302 400898 113334 401134
rect 112714 383454 113334 400898
rect 112714 383218 112746 383454
rect 112982 383218 113066 383454
rect 113302 383218 113334 383454
rect 112714 383134 113334 383218
rect 112714 382898 112746 383134
rect 112982 382898 113066 383134
rect 113302 382898 113334 383134
rect 112714 365454 113334 382898
rect 112714 365218 112746 365454
rect 112982 365218 113066 365454
rect 113302 365218 113334 365454
rect 112714 365134 113334 365218
rect 112714 364898 112746 365134
rect 112982 364898 113066 365134
rect 113302 364898 113334 365134
rect 112714 347454 113334 364898
rect 112714 347218 112746 347454
rect 112982 347218 113066 347454
rect 113302 347218 113334 347454
rect 112714 347134 113334 347218
rect 112714 346898 112746 347134
rect 112982 346898 113066 347134
rect 113302 346898 113334 347134
rect 112714 329454 113334 346898
rect 112714 329218 112746 329454
rect 112982 329218 113066 329454
rect 113302 329218 113334 329454
rect 112714 329134 113334 329218
rect 112714 328898 112746 329134
rect 112982 328898 113066 329134
rect 113302 328898 113334 329134
rect 112714 311454 113334 328898
rect 112714 311218 112746 311454
rect 112982 311218 113066 311454
rect 113302 311218 113334 311454
rect 112714 311134 113334 311218
rect 112714 310898 112746 311134
rect 112982 310898 113066 311134
rect 113302 310898 113334 311134
rect 112714 293454 113334 310898
rect 112714 293218 112746 293454
rect 112982 293218 113066 293454
rect 113302 293218 113334 293454
rect 112714 293134 113334 293218
rect 112714 292898 112746 293134
rect 112982 292898 113066 293134
rect 113302 292898 113334 293134
rect 112714 275454 113334 292898
rect 112714 275218 112746 275454
rect 112982 275218 113066 275454
rect 113302 275218 113334 275454
rect 112714 275134 113334 275218
rect 112714 274898 112746 275134
rect 112982 274898 113066 275134
rect 113302 274898 113334 275134
rect 112714 257454 113334 274898
rect 112714 257218 112746 257454
rect 112982 257218 113066 257454
rect 113302 257218 113334 257454
rect 112714 257134 113334 257218
rect 112714 256898 112746 257134
rect 112982 256898 113066 257134
rect 113302 256898 113334 257134
rect 112714 239454 113334 256898
rect 112714 239218 112746 239454
rect 112982 239218 113066 239454
rect 113302 239218 113334 239454
rect 112714 239134 113334 239218
rect 112714 238898 112746 239134
rect 112982 238898 113066 239134
rect 113302 238898 113334 239134
rect 112714 221454 113334 238898
rect 112714 221218 112746 221454
rect 112982 221218 113066 221454
rect 113302 221218 113334 221454
rect 112714 221134 113334 221218
rect 112714 220898 112746 221134
rect 112982 220898 113066 221134
rect 113302 220898 113334 221134
rect 112714 203454 113334 220898
rect 112714 203218 112746 203454
rect 112982 203218 113066 203454
rect 113302 203218 113334 203454
rect 112714 203134 113334 203218
rect 112714 202898 112746 203134
rect 112982 202898 113066 203134
rect 113302 202898 113334 203134
rect 112714 185454 113334 202898
rect 112714 185218 112746 185454
rect 112982 185218 113066 185454
rect 113302 185218 113334 185454
rect 112714 185134 113334 185218
rect 112714 184898 112746 185134
rect 112982 184898 113066 185134
rect 113302 184898 113334 185134
rect 112714 167454 113334 184898
rect 112714 167218 112746 167454
rect 112982 167218 113066 167454
rect 113302 167218 113334 167454
rect 112714 167134 113334 167218
rect 112714 166898 112746 167134
rect 112982 166898 113066 167134
rect 113302 166898 113334 167134
rect 112714 149454 113334 166898
rect 112714 149218 112746 149454
rect 112982 149218 113066 149454
rect 113302 149218 113334 149454
rect 112714 149134 113334 149218
rect 112714 148898 112746 149134
rect 112982 148898 113066 149134
rect 113302 148898 113334 149134
rect 112714 131454 113334 148898
rect 112714 131218 112746 131454
rect 112982 131218 113066 131454
rect 113302 131218 113334 131454
rect 112714 131134 113334 131218
rect 112714 130898 112746 131134
rect 112982 130898 113066 131134
rect 113302 130898 113334 131134
rect 112714 113454 113334 130898
rect 112714 113218 112746 113454
rect 112982 113218 113066 113454
rect 113302 113218 113334 113454
rect 112714 113134 113334 113218
rect 112714 112898 112746 113134
rect 112982 112898 113066 113134
rect 113302 112898 113334 113134
rect 112714 95454 113334 112898
rect 112714 95218 112746 95454
rect 112982 95218 113066 95454
rect 113302 95218 113334 95454
rect 112714 95134 113334 95218
rect 112714 94898 112746 95134
rect 112982 94898 113066 95134
rect 113302 94898 113334 95134
rect 112714 77454 113334 94898
rect 112714 77218 112746 77454
rect 112982 77218 113066 77454
rect 113302 77218 113334 77454
rect 112714 77134 113334 77218
rect 112714 76898 112746 77134
rect 112982 76898 113066 77134
rect 113302 76898 113334 77134
rect 112714 59454 113334 76898
rect 112714 59218 112746 59454
rect 112982 59218 113066 59454
rect 113302 59218 113334 59454
rect 112714 59134 113334 59218
rect 112714 58898 112746 59134
rect 112982 58898 113066 59134
rect 113302 58898 113334 59134
rect 112714 58629 113334 58898
rect 116434 462052 117054 464004
rect 116434 461816 116466 462052
rect 116702 461816 116786 462052
rect 117022 461816 117054 462052
rect 116434 461732 117054 461816
rect 116434 461496 116466 461732
rect 116702 461496 116786 461732
rect 117022 461496 117054 461732
rect 116434 441174 117054 461496
rect 116434 440938 116466 441174
rect 116702 440938 116786 441174
rect 117022 440938 117054 441174
rect 116434 440854 117054 440938
rect 116434 440618 116466 440854
rect 116702 440618 116786 440854
rect 117022 440618 117054 440854
rect 116434 423174 117054 440618
rect 116434 422938 116466 423174
rect 116702 422938 116786 423174
rect 117022 422938 117054 423174
rect 116434 422854 117054 422938
rect 116434 422618 116466 422854
rect 116702 422618 116786 422854
rect 117022 422618 117054 422854
rect 116434 405174 117054 422618
rect 116434 404938 116466 405174
rect 116702 404938 116786 405174
rect 117022 404938 117054 405174
rect 116434 404854 117054 404938
rect 116434 404618 116466 404854
rect 116702 404618 116786 404854
rect 117022 404618 117054 404854
rect 116434 387174 117054 404618
rect 116434 386938 116466 387174
rect 116702 386938 116786 387174
rect 117022 386938 117054 387174
rect 116434 386854 117054 386938
rect 116434 386618 116466 386854
rect 116702 386618 116786 386854
rect 117022 386618 117054 386854
rect 116434 369174 117054 386618
rect 116434 368938 116466 369174
rect 116702 368938 116786 369174
rect 117022 368938 117054 369174
rect 116434 368854 117054 368938
rect 116434 368618 116466 368854
rect 116702 368618 116786 368854
rect 117022 368618 117054 368854
rect 116434 351174 117054 368618
rect 116434 350938 116466 351174
rect 116702 350938 116786 351174
rect 117022 350938 117054 351174
rect 116434 350854 117054 350938
rect 116434 350618 116466 350854
rect 116702 350618 116786 350854
rect 117022 350618 117054 350854
rect 116434 333174 117054 350618
rect 116434 332938 116466 333174
rect 116702 332938 116786 333174
rect 117022 332938 117054 333174
rect 116434 332854 117054 332938
rect 116434 332618 116466 332854
rect 116702 332618 116786 332854
rect 117022 332618 117054 332854
rect 116434 315174 117054 332618
rect 116434 314938 116466 315174
rect 116702 314938 116786 315174
rect 117022 314938 117054 315174
rect 116434 314854 117054 314938
rect 116434 314618 116466 314854
rect 116702 314618 116786 314854
rect 117022 314618 117054 314854
rect 116434 297174 117054 314618
rect 116434 296938 116466 297174
rect 116702 296938 116786 297174
rect 117022 296938 117054 297174
rect 116434 296854 117054 296938
rect 116434 296618 116466 296854
rect 116702 296618 116786 296854
rect 117022 296618 117054 296854
rect 116434 279174 117054 296618
rect 116434 278938 116466 279174
rect 116702 278938 116786 279174
rect 117022 278938 117054 279174
rect 116434 278854 117054 278938
rect 116434 278618 116466 278854
rect 116702 278618 116786 278854
rect 117022 278618 117054 278854
rect 116434 261174 117054 278618
rect 116434 260938 116466 261174
rect 116702 260938 116786 261174
rect 117022 260938 117054 261174
rect 116434 260854 117054 260938
rect 116434 260618 116466 260854
rect 116702 260618 116786 260854
rect 117022 260618 117054 260854
rect 116434 243174 117054 260618
rect 116434 242938 116466 243174
rect 116702 242938 116786 243174
rect 117022 242938 117054 243174
rect 116434 242854 117054 242938
rect 116434 242618 116466 242854
rect 116702 242618 116786 242854
rect 117022 242618 117054 242854
rect 116434 225174 117054 242618
rect 116434 224938 116466 225174
rect 116702 224938 116786 225174
rect 117022 224938 117054 225174
rect 116434 224854 117054 224938
rect 116434 224618 116466 224854
rect 116702 224618 116786 224854
rect 117022 224618 117054 224854
rect 116434 207174 117054 224618
rect 116434 206938 116466 207174
rect 116702 206938 116786 207174
rect 117022 206938 117054 207174
rect 116434 206854 117054 206938
rect 116434 206618 116466 206854
rect 116702 206618 116786 206854
rect 117022 206618 117054 206854
rect 116434 189174 117054 206618
rect 116434 188938 116466 189174
rect 116702 188938 116786 189174
rect 117022 188938 117054 189174
rect 116434 188854 117054 188938
rect 116434 188618 116466 188854
rect 116702 188618 116786 188854
rect 117022 188618 117054 188854
rect 116434 171174 117054 188618
rect 116434 170938 116466 171174
rect 116702 170938 116786 171174
rect 117022 170938 117054 171174
rect 116434 170854 117054 170938
rect 116434 170618 116466 170854
rect 116702 170618 116786 170854
rect 117022 170618 117054 170854
rect 116434 153174 117054 170618
rect 116434 152938 116466 153174
rect 116702 152938 116786 153174
rect 117022 152938 117054 153174
rect 116434 152854 117054 152938
rect 116434 152618 116466 152854
rect 116702 152618 116786 152854
rect 117022 152618 117054 152854
rect 116434 135174 117054 152618
rect 116434 134938 116466 135174
rect 116702 134938 116786 135174
rect 117022 134938 117054 135174
rect 116434 134854 117054 134938
rect 116434 134618 116466 134854
rect 116702 134618 116786 134854
rect 117022 134618 117054 134854
rect 116434 117174 117054 134618
rect 116434 116938 116466 117174
rect 116702 116938 116786 117174
rect 117022 116938 117054 117174
rect 116434 116854 117054 116938
rect 116434 116618 116466 116854
rect 116702 116618 116786 116854
rect 117022 116618 117054 116854
rect 116434 99174 117054 116618
rect 116434 98938 116466 99174
rect 116702 98938 116786 99174
rect 117022 98938 117054 99174
rect 116434 98854 117054 98938
rect 116434 98618 116466 98854
rect 116702 98618 116786 98854
rect 117022 98618 117054 98854
rect 116434 81174 117054 98618
rect 116434 80938 116466 81174
rect 116702 80938 116786 81174
rect 117022 80938 117054 81174
rect 116434 80854 117054 80938
rect 116434 80618 116466 80854
rect 116702 80618 116786 80854
rect 117022 80618 117054 80854
rect 116434 63174 117054 80618
rect 116434 62938 116466 63174
rect 116702 62938 116786 63174
rect 117022 62938 117054 63174
rect 116434 62854 117054 62938
rect 116434 62618 116466 62854
rect 116702 62618 116786 62854
rect 117022 62618 117054 62854
rect 116434 58629 117054 62618
rect 120154 463012 120774 464004
rect 120154 462776 120186 463012
rect 120422 462776 120506 463012
rect 120742 462776 120774 463012
rect 120154 462692 120774 462776
rect 120154 462456 120186 462692
rect 120422 462456 120506 462692
rect 120742 462456 120774 462692
rect 120154 444894 120774 462456
rect 120154 444658 120186 444894
rect 120422 444658 120506 444894
rect 120742 444658 120774 444894
rect 120154 444574 120774 444658
rect 120154 444338 120186 444574
rect 120422 444338 120506 444574
rect 120742 444338 120774 444574
rect 120154 426894 120774 444338
rect 120154 426658 120186 426894
rect 120422 426658 120506 426894
rect 120742 426658 120774 426894
rect 120154 426574 120774 426658
rect 120154 426338 120186 426574
rect 120422 426338 120506 426574
rect 120742 426338 120774 426574
rect 120154 408894 120774 426338
rect 120154 408658 120186 408894
rect 120422 408658 120506 408894
rect 120742 408658 120774 408894
rect 120154 408574 120774 408658
rect 120154 408338 120186 408574
rect 120422 408338 120506 408574
rect 120742 408338 120774 408574
rect 120154 390894 120774 408338
rect 120154 390658 120186 390894
rect 120422 390658 120506 390894
rect 120742 390658 120774 390894
rect 120154 390574 120774 390658
rect 120154 390338 120186 390574
rect 120422 390338 120506 390574
rect 120742 390338 120774 390574
rect 120154 372894 120774 390338
rect 120154 372658 120186 372894
rect 120422 372658 120506 372894
rect 120742 372658 120774 372894
rect 120154 372574 120774 372658
rect 120154 372338 120186 372574
rect 120422 372338 120506 372574
rect 120742 372338 120774 372574
rect 120154 354894 120774 372338
rect 120154 354658 120186 354894
rect 120422 354658 120506 354894
rect 120742 354658 120774 354894
rect 120154 354574 120774 354658
rect 120154 354338 120186 354574
rect 120422 354338 120506 354574
rect 120742 354338 120774 354574
rect 120154 336894 120774 354338
rect 120154 336658 120186 336894
rect 120422 336658 120506 336894
rect 120742 336658 120774 336894
rect 120154 336574 120774 336658
rect 120154 336338 120186 336574
rect 120422 336338 120506 336574
rect 120742 336338 120774 336574
rect 120154 318894 120774 336338
rect 120154 318658 120186 318894
rect 120422 318658 120506 318894
rect 120742 318658 120774 318894
rect 120154 318574 120774 318658
rect 120154 318338 120186 318574
rect 120422 318338 120506 318574
rect 120742 318338 120774 318574
rect 120154 300894 120774 318338
rect 120154 300658 120186 300894
rect 120422 300658 120506 300894
rect 120742 300658 120774 300894
rect 120154 300574 120774 300658
rect 120154 300338 120186 300574
rect 120422 300338 120506 300574
rect 120742 300338 120774 300574
rect 120154 282894 120774 300338
rect 120154 282658 120186 282894
rect 120422 282658 120506 282894
rect 120742 282658 120774 282894
rect 120154 282574 120774 282658
rect 120154 282338 120186 282574
rect 120422 282338 120506 282574
rect 120742 282338 120774 282574
rect 120154 264894 120774 282338
rect 120154 264658 120186 264894
rect 120422 264658 120506 264894
rect 120742 264658 120774 264894
rect 120154 264574 120774 264658
rect 120154 264338 120186 264574
rect 120422 264338 120506 264574
rect 120742 264338 120774 264574
rect 120154 246894 120774 264338
rect 120154 246658 120186 246894
rect 120422 246658 120506 246894
rect 120742 246658 120774 246894
rect 120154 246574 120774 246658
rect 120154 246338 120186 246574
rect 120422 246338 120506 246574
rect 120742 246338 120774 246574
rect 120154 228894 120774 246338
rect 120154 228658 120186 228894
rect 120422 228658 120506 228894
rect 120742 228658 120774 228894
rect 120154 228574 120774 228658
rect 120154 228338 120186 228574
rect 120422 228338 120506 228574
rect 120742 228338 120774 228574
rect 120154 210894 120774 228338
rect 120154 210658 120186 210894
rect 120422 210658 120506 210894
rect 120742 210658 120774 210894
rect 120154 210574 120774 210658
rect 120154 210338 120186 210574
rect 120422 210338 120506 210574
rect 120742 210338 120774 210574
rect 120154 192894 120774 210338
rect 120154 192658 120186 192894
rect 120422 192658 120506 192894
rect 120742 192658 120774 192894
rect 120154 192574 120774 192658
rect 120154 192338 120186 192574
rect 120422 192338 120506 192574
rect 120742 192338 120774 192574
rect 120154 174894 120774 192338
rect 120154 174658 120186 174894
rect 120422 174658 120506 174894
rect 120742 174658 120774 174894
rect 120154 174574 120774 174658
rect 120154 174338 120186 174574
rect 120422 174338 120506 174574
rect 120742 174338 120774 174574
rect 120154 156894 120774 174338
rect 120154 156658 120186 156894
rect 120422 156658 120506 156894
rect 120742 156658 120774 156894
rect 120154 156574 120774 156658
rect 120154 156338 120186 156574
rect 120422 156338 120506 156574
rect 120742 156338 120774 156574
rect 120154 138894 120774 156338
rect 120154 138658 120186 138894
rect 120422 138658 120506 138894
rect 120742 138658 120774 138894
rect 120154 138574 120774 138658
rect 120154 138338 120186 138574
rect 120422 138338 120506 138574
rect 120742 138338 120774 138574
rect 120154 120894 120774 138338
rect 120154 120658 120186 120894
rect 120422 120658 120506 120894
rect 120742 120658 120774 120894
rect 120154 120574 120774 120658
rect 120154 120338 120186 120574
rect 120422 120338 120506 120574
rect 120742 120338 120774 120574
rect 120154 102894 120774 120338
rect 120154 102658 120186 102894
rect 120422 102658 120506 102894
rect 120742 102658 120774 102894
rect 120154 102574 120774 102658
rect 120154 102338 120186 102574
rect 120422 102338 120506 102574
rect 120742 102338 120774 102574
rect 120154 84894 120774 102338
rect 120154 84658 120186 84894
rect 120422 84658 120506 84894
rect 120742 84658 120774 84894
rect 120154 84574 120774 84658
rect 120154 84338 120186 84574
rect 120422 84338 120506 84574
rect 120742 84338 120774 84574
rect 120154 66894 120774 84338
rect 120154 66658 120186 66894
rect 120422 66658 120506 66894
rect 120742 66658 120774 66894
rect 120154 66574 120774 66658
rect 120154 66338 120186 66574
rect 120422 66338 120506 66574
rect 120742 66338 120774 66574
rect 120154 58629 120774 66338
rect 123874 463972 124494 464004
rect 123874 463736 123906 463972
rect 124142 463736 124226 463972
rect 124462 463736 124494 463972
rect 123874 463652 124494 463736
rect 123874 463416 123906 463652
rect 124142 463416 124226 463652
rect 124462 463416 124494 463652
rect 123874 448614 124494 463416
rect 123874 448378 123906 448614
rect 124142 448378 124226 448614
rect 124462 448378 124494 448614
rect 123874 448294 124494 448378
rect 123874 448058 123906 448294
rect 124142 448058 124226 448294
rect 124462 448058 124494 448294
rect 123874 430614 124494 448058
rect 123874 430378 123906 430614
rect 124142 430378 124226 430614
rect 124462 430378 124494 430614
rect 123874 430294 124494 430378
rect 123874 430058 123906 430294
rect 124142 430058 124226 430294
rect 124462 430058 124494 430294
rect 123874 412614 124494 430058
rect 123874 412378 123906 412614
rect 124142 412378 124226 412614
rect 124462 412378 124494 412614
rect 123874 412294 124494 412378
rect 123874 412058 123906 412294
rect 124142 412058 124226 412294
rect 124462 412058 124494 412294
rect 123874 394614 124494 412058
rect 123874 394378 123906 394614
rect 124142 394378 124226 394614
rect 124462 394378 124494 394614
rect 123874 394294 124494 394378
rect 123874 394058 123906 394294
rect 124142 394058 124226 394294
rect 124462 394058 124494 394294
rect 123874 376614 124494 394058
rect 123874 376378 123906 376614
rect 124142 376378 124226 376614
rect 124462 376378 124494 376614
rect 123874 376294 124494 376378
rect 123874 376058 123906 376294
rect 124142 376058 124226 376294
rect 124462 376058 124494 376294
rect 123874 358614 124494 376058
rect 123874 358378 123906 358614
rect 124142 358378 124226 358614
rect 124462 358378 124494 358614
rect 123874 358294 124494 358378
rect 123874 358058 123906 358294
rect 124142 358058 124226 358294
rect 124462 358058 124494 358294
rect 123874 340614 124494 358058
rect 123874 340378 123906 340614
rect 124142 340378 124226 340614
rect 124462 340378 124494 340614
rect 123874 340294 124494 340378
rect 123874 340058 123906 340294
rect 124142 340058 124226 340294
rect 124462 340058 124494 340294
rect 123874 322614 124494 340058
rect 123874 322378 123906 322614
rect 124142 322378 124226 322614
rect 124462 322378 124494 322614
rect 123874 322294 124494 322378
rect 123874 322058 123906 322294
rect 124142 322058 124226 322294
rect 124462 322058 124494 322294
rect 123874 304614 124494 322058
rect 123874 304378 123906 304614
rect 124142 304378 124226 304614
rect 124462 304378 124494 304614
rect 123874 304294 124494 304378
rect 123874 304058 123906 304294
rect 124142 304058 124226 304294
rect 124462 304058 124494 304294
rect 123874 286614 124494 304058
rect 123874 286378 123906 286614
rect 124142 286378 124226 286614
rect 124462 286378 124494 286614
rect 123874 286294 124494 286378
rect 123874 286058 123906 286294
rect 124142 286058 124226 286294
rect 124462 286058 124494 286294
rect 123874 268614 124494 286058
rect 123874 268378 123906 268614
rect 124142 268378 124226 268614
rect 124462 268378 124494 268614
rect 123874 268294 124494 268378
rect 123874 268058 123906 268294
rect 124142 268058 124226 268294
rect 124462 268058 124494 268294
rect 123874 250614 124494 268058
rect 123874 250378 123906 250614
rect 124142 250378 124226 250614
rect 124462 250378 124494 250614
rect 123874 250294 124494 250378
rect 123874 250058 123906 250294
rect 124142 250058 124226 250294
rect 124462 250058 124494 250294
rect 123874 232614 124494 250058
rect 123874 232378 123906 232614
rect 124142 232378 124226 232614
rect 124462 232378 124494 232614
rect 123874 232294 124494 232378
rect 123874 232058 123906 232294
rect 124142 232058 124226 232294
rect 124462 232058 124494 232294
rect 123874 214614 124494 232058
rect 123874 214378 123906 214614
rect 124142 214378 124226 214614
rect 124462 214378 124494 214614
rect 123874 214294 124494 214378
rect 123874 214058 123906 214294
rect 124142 214058 124226 214294
rect 124462 214058 124494 214294
rect 123874 196614 124494 214058
rect 123874 196378 123906 196614
rect 124142 196378 124226 196614
rect 124462 196378 124494 196614
rect 123874 196294 124494 196378
rect 123874 196058 123906 196294
rect 124142 196058 124226 196294
rect 124462 196058 124494 196294
rect 123874 178614 124494 196058
rect 123874 178378 123906 178614
rect 124142 178378 124226 178614
rect 124462 178378 124494 178614
rect 123874 178294 124494 178378
rect 123874 178058 123906 178294
rect 124142 178058 124226 178294
rect 124462 178058 124494 178294
rect 123874 160614 124494 178058
rect 123874 160378 123906 160614
rect 124142 160378 124226 160614
rect 124462 160378 124494 160614
rect 123874 160294 124494 160378
rect 123874 160058 123906 160294
rect 124142 160058 124226 160294
rect 124462 160058 124494 160294
rect 123874 142614 124494 160058
rect 123874 142378 123906 142614
rect 124142 142378 124226 142614
rect 124462 142378 124494 142614
rect 123874 142294 124494 142378
rect 123874 142058 123906 142294
rect 124142 142058 124226 142294
rect 124462 142058 124494 142294
rect 123874 124614 124494 142058
rect 123874 124378 123906 124614
rect 124142 124378 124226 124614
rect 124462 124378 124494 124614
rect 123874 124294 124494 124378
rect 123874 124058 123906 124294
rect 124142 124058 124226 124294
rect 124462 124058 124494 124294
rect 123874 106614 124494 124058
rect 123874 106378 123906 106614
rect 124142 106378 124226 106614
rect 124462 106378 124494 106614
rect 123874 106294 124494 106378
rect 123874 106058 123906 106294
rect 124142 106058 124226 106294
rect 124462 106058 124494 106294
rect 123874 88614 124494 106058
rect 123874 88378 123906 88614
rect 124142 88378 124226 88614
rect 124462 88378 124494 88614
rect 123874 88294 124494 88378
rect 123874 88058 123906 88294
rect 124142 88058 124226 88294
rect 124462 88058 124494 88294
rect 123874 70614 124494 88058
rect 123874 70378 123906 70614
rect 124142 70378 124226 70614
rect 124462 70378 124494 70614
rect 123874 70294 124494 70378
rect 123874 70058 123906 70294
rect 124142 70058 124226 70294
rect 124462 70058 124494 70294
rect 123874 58629 124494 70058
rect 130714 461092 131334 464004
rect 130714 460856 130746 461092
rect 130982 460856 131066 461092
rect 131302 460856 131334 461092
rect 130714 460772 131334 460856
rect 130714 460536 130746 460772
rect 130982 460536 131066 460772
rect 131302 460536 131334 460772
rect 130714 455454 131334 460536
rect 130714 455218 130746 455454
rect 130982 455218 131066 455454
rect 131302 455218 131334 455454
rect 130714 455134 131334 455218
rect 130714 454898 130746 455134
rect 130982 454898 131066 455134
rect 131302 454898 131334 455134
rect 130714 437454 131334 454898
rect 130714 437218 130746 437454
rect 130982 437218 131066 437454
rect 131302 437218 131334 437454
rect 130714 437134 131334 437218
rect 130714 436898 130746 437134
rect 130982 436898 131066 437134
rect 131302 436898 131334 437134
rect 130714 419454 131334 436898
rect 130714 419218 130746 419454
rect 130982 419218 131066 419454
rect 131302 419218 131334 419454
rect 130714 419134 131334 419218
rect 130714 418898 130746 419134
rect 130982 418898 131066 419134
rect 131302 418898 131334 419134
rect 130714 401454 131334 418898
rect 130714 401218 130746 401454
rect 130982 401218 131066 401454
rect 131302 401218 131334 401454
rect 130714 401134 131334 401218
rect 130714 400898 130746 401134
rect 130982 400898 131066 401134
rect 131302 400898 131334 401134
rect 130714 383454 131334 400898
rect 130714 383218 130746 383454
rect 130982 383218 131066 383454
rect 131302 383218 131334 383454
rect 130714 383134 131334 383218
rect 130714 382898 130746 383134
rect 130982 382898 131066 383134
rect 131302 382898 131334 383134
rect 130714 365454 131334 382898
rect 130714 365218 130746 365454
rect 130982 365218 131066 365454
rect 131302 365218 131334 365454
rect 130714 365134 131334 365218
rect 130714 364898 130746 365134
rect 130982 364898 131066 365134
rect 131302 364898 131334 365134
rect 130714 347454 131334 364898
rect 130714 347218 130746 347454
rect 130982 347218 131066 347454
rect 131302 347218 131334 347454
rect 130714 347134 131334 347218
rect 130714 346898 130746 347134
rect 130982 346898 131066 347134
rect 131302 346898 131334 347134
rect 130714 329454 131334 346898
rect 130714 329218 130746 329454
rect 130982 329218 131066 329454
rect 131302 329218 131334 329454
rect 130714 329134 131334 329218
rect 130714 328898 130746 329134
rect 130982 328898 131066 329134
rect 131302 328898 131334 329134
rect 130714 311454 131334 328898
rect 130714 311218 130746 311454
rect 130982 311218 131066 311454
rect 131302 311218 131334 311454
rect 130714 311134 131334 311218
rect 130714 310898 130746 311134
rect 130982 310898 131066 311134
rect 131302 310898 131334 311134
rect 130714 293454 131334 310898
rect 130714 293218 130746 293454
rect 130982 293218 131066 293454
rect 131302 293218 131334 293454
rect 130714 293134 131334 293218
rect 130714 292898 130746 293134
rect 130982 292898 131066 293134
rect 131302 292898 131334 293134
rect 130714 275454 131334 292898
rect 130714 275218 130746 275454
rect 130982 275218 131066 275454
rect 131302 275218 131334 275454
rect 130714 275134 131334 275218
rect 130714 274898 130746 275134
rect 130982 274898 131066 275134
rect 131302 274898 131334 275134
rect 130714 257454 131334 274898
rect 130714 257218 130746 257454
rect 130982 257218 131066 257454
rect 131302 257218 131334 257454
rect 130714 257134 131334 257218
rect 130714 256898 130746 257134
rect 130982 256898 131066 257134
rect 131302 256898 131334 257134
rect 130714 239454 131334 256898
rect 130714 239218 130746 239454
rect 130982 239218 131066 239454
rect 131302 239218 131334 239454
rect 130714 239134 131334 239218
rect 130714 238898 130746 239134
rect 130982 238898 131066 239134
rect 131302 238898 131334 239134
rect 130714 221454 131334 238898
rect 130714 221218 130746 221454
rect 130982 221218 131066 221454
rect 131302 221218 131334 221454
rect 130714 221134 131334 221218
rect 130714 220898 130746 221134
rect 130982 220898 131066 221134
rect 131302 220898 131334 221134
rect 130714 203454 131334 220898
rect 130714 203218 130746 203454
rect 130982 203218 131066 203454
rect 131302 203218 131334 203454
rect 130714 203134 131334 203218
rect 130714 202898 130746 203134
rect 130982 202898 131066 203134
rect 131302 202898 131334 203134
rect 130714 185454 131334 202898
rect 130714 185218 130746 185454
rect 130982 185218 131066 185454
rect 131302 185218 131334 185454
rect 130714 185134 131334 185218
rect 130714 184898 130746 185134
rect 130982 184898 131066 185134
rect 131302 184898 131334 185134
rect 130714 167454 131334 184898
rect 130714 167218 130746 167454
rect 130982 167218 131066 167454
rect 131302 167218 131334 167454
rect 130714 167134 131334 167218
rect 130714 166898 130746 167134
rect 130982 166898 131066 167134
rect 131302 166898 131334 167134
rect 130714 149454 131334 166898
rect 130714 149218 130746 149454
rect 130982 149218 131066 149454
rect 131302 149218 131334 149454
rect 130714 149134 131334 149218
rect 130714 148898 130746 149134
rect 130982 148898 131066 149134
rect 131302 148898 131334 149134
rect 130714 131454 131334 148898
rect 130714 131218 130746 131454
rect 130982 131218 131066 131454
rect 131302 131218 131334 131454
rect 130714 131134 131334 131218
rect 130714 130898 130746 131134
rect 130982 130898 131066 131134
rect 131302 130898 131334 131134
rect 130714 113454 131334 130898
rect 130714 113218 130746 113454
rect 130982 113218 131066 113454
rect 131302 113218 131334 113454
rect 130714 113134 131334 113218
rect 130714 112898 130746 113134
rect 130982 112898 131066 113134
rect 131302 112898 131334 113134
rect 130714 95454 131334 112898
rect 130714 95218 130746 95454
rect 130982 95218 131066 95454
rect 131302 95218 131334 95454
rect 130714 95134 131334 95218
rect 130714 94898 130746 95134
rect 130982 94898 131066 95134
rect 131302 94898 131334 95134
rect 130714 77454 131334 94898
rect 130714 77218 130746 77454
rect 130982 77218 131066 77454
rect 131302 77218 131334 77454
rect 130714 77134 131334 77218
rect 130714 76898 130746 77134
rect 130982 76898 131066 77134
rect 131302 76898 131334 77134
rect 130714 59454 131334 76898
rect 130714 59218 130746 59454
rect 130982 59218 131066 59454
rect 131302 59218 131334 59454
rect 130714 59134 131334 59218
rect 130714 58898 130746 59134
rect 130982 58898 131066 59134
rect 131302 58898 131334 59134
rect 130714 58629 131334 58898
rect 134434 462052 135054 464004
rect 134434 461816 134466 462052
rect 134702 461816 134786 462052
rect 135022 461816 135054 462052
rect 134434 461732 135054 461816
rect 134434 461496 134466 461732
rect 134702 461496 134786 461732
rect 135022 461496 135054 461732
rect 134434 441174 135054 461496
rect 134434 440938 134466 441174
rect 134702 440938 134786 441174
rect 135022 440938 135054 441174
rect 134434 440854 135054 440938
rect 134434 440618 134466 440854
rect 134702 440618 134786 440854
rect 135022 440618 135054 440854
rect 134434 423174 135054 440618
rect 134434 422938 134466 423174
rect 134702 422938 134786 423174
rect 135022 422938 135054 423174
rect 134434 422854 135054 422938
rect 134434 422618 134466 422854
rect 134702 422618 134786 422854
rect 135022 422618 135054 422854
rect 134434 405174 135054 422618
rect 134434 404938 134466 405174
rect 134702 404938 134786 405174
rect 135022 404938 135054 405174
rect 134434 404854 135054 404938
rect 134434 404618 134466 404854
rect 134702 404618 134786 404854
rect 135022 404618 135054 404854
rect 134434 387174 135054 404618
rect 134434 386938 134466 387174
rect 134702 386938 134786 387174
rect 135022 386938 135054 387174
rect 134434 386854 135054 386938
rect 134434 386618 134466 386854
rect 134702 386618 134786 386854
rect 135022 386618 135054 386854
rect 134434 369174 135054 386618
rect 134434 368938 134466 369174
rect 134702 368938 134786 369174
rect 135022 368938 135054 369174
rect 134434 368854 135054 368938
rect 134434 368618 134466 368854
rect 134702 368618 134786 368854
rect 135022 368618 135054 368854
rect 134434 351174 135054 368618
rect 134434 350938 134466 351174
rect 134702 350938 134786 351174
rect 135022 350938 135054 351174
rect 134434 350854 135054 350938
rect 134434 350618 134466 350854
rect 134702 350618 134786 350854
rect 135022 350618 135054 350854
rect 134434 333174 135054 350618
rect 134434 332938 134466 333174
rect 134702 332938 134786 333174
rect 135022 332938 135054 333174
rect 134434 332854 135054 332938
rect 134434 332618 134466 332854
rect 134702 332618 134786 332854
rect 135022 332618 135054 332854
rect 134434 315174 135054 332618
rect 134434 314938 134466 315174
rect 134702 314938 134786 315174
rect 135022 314938 135054 315174
rect 134434 314854 135054 314938
rect 134434 314618 134466 314854
rect 134702 314618 134786 314854
rect 135022 314618 135054 314854
rect 134434 297174 135054 314618
rect 134434 296938 134466 297174
rect 134702 296938 134786 297174
rect 135022 296938 135054 297174
rect 134434 296854 135054 296938
rect 134434 296618 134466 296854
rect 134702 296618 134786 296854
rect 135022 296618 135054 296854
rect 134434 279174 135054 296618
rect 134434 278938 134466 279174
rect 134702 278938 134786 279174
rect 135022 278938 135054 279174
rect 134434 278854 135054 278938
rect 134434 278618 134466 278854
rect 134702 278618 134786 278854
rect 135022 278618 135054 278854
rect 134434 261174 135054 278618
rect 134434 260938 134466 261174
rect 134702 260938 134786 261174
rect 135022 260938 135054 261174
rect 134434 260854 135054 260938
rect 134434 260618 134466 260854
rect 134702 260618 134786 260854
rect 135022 260618 135054 260854
rect 134434 243174 135054 260618
rect 134434 242938 134466 243174
rect 134702 242938 134786 243174
rect 135022 242938 135054 243174
rect 134434 242854 135054 242938
rect 134434 242618 134466 242854
rect 134702 242618 134786 242854
rect 135022 242618 135054 242854
rect 134434 225174 135054 242618
rect 134434 224938 134466 225174
rect 134702 224938 134786 225174
rect 135022 224938 135054 225174
rect 134434 224854 135054 224938
rect 134434 224618 134466 224854
rect 134702 224618 134786 224854
rect 135022 224618 135054 224854
rect 134434 207174 135054 224618
rect 134434 206938 134466 207174
rect 134702 206938 134786 207174
rect 135022 206938 135054 207174
rect 134434 206854 135054 206938
rect 134434 206618 134466 206854
rect 134702 206618 134786 206854
rect 135022 206618 135054 206854
rect 134434 189174 135054 206618
rect 134434 188938 134466 189174
rect 134702 188938 134786 189174
rect 135022 188938 135054 189174
rect 134434 188854 135054 188938
rect 134434 188618 134466 188854
rect 134702 188618 134786 188854
rect 135022 188618 135054 188854
rect 134434 171174 135054 188618
rect 134434 170938 134466 171174
rect 134702 170938 134786 171174
rect 135022 170938 135054 171174
rect 134434 170854 135054 170938
rect 134434 170618 134466 170854
rect 134702 170618 134786 170854
rect 135022 170618 135054 170854
rect 134434 153174 135054 170618
rect 134434 152938 134466 153174
rect 134702 152938 134786 153174
rect 135022 152938 135054 153174
rect 134434 152854 135054 152938
rect 134434 152618 134466 152854
rect 134702 152618 134786 152854
rect 135022 152618 135054 152854
rect 134434 135174 135054 152618
rect 134434 134938 134466 135174
rect 134702 134938 134786 135174
rect 135022 134938 135054 135174
rect 134434 134854 135054 134938
rect 134434 134618 134466 134854
rect 134702 134618 134786 134854
rect 135022 134618 135054 134854
rect 134434 117174 135054 134618
rect 134434 116938 134466 117174
rect 134702 116938 134786 117174
rect 135022 116938 135054 117174
rect 134434 116854 135054 116938
rect 134434 116618 134466 116854
rect 134702 116618 134786 116854
rect 135022 116618 135054 116854
rect 134434 99174 135054 116618
rect 134434 98938 134466 99174
rect 134702 98938 134786 99174
rect 135022 98938 135054 99174
rect 134434 98854 135054 98938
rect 134434 98618 134466 98854
rect 134702 98618 134786 98854
rect 135022 98618 135054 98854
rect 134434 81174 135054 98618
rect 134434 80938 134466 81174
rect 134702 80938 134786 81174
rect 135022 80938 135054 81174
rect 134434 80854 135054 80938
rect 134434 80618 134466 80854
rect 134702 80618 134786 80854
rect 135022 80618 135054 80854
rect 134434 63174 135054 80618
rect 134434 62938 134466 63174
rect 134702 62938 134786 63174
rect 135022 62938 135054 63174
rect 134434 62854 135054 62938
rect 134434 62618 134466 62854
rect 134702 62618 134786 62854
rect 135022 62618 135054 62854
rect 87874 52378 87906 52614
rect 88142 52378 88226 52614
rect 88462 52378 88494 52614
rect 87874 52294 88494 52378
rect 87874 52058 87906 52294
rect 88142 52058 88226 52294
rect 88462 52058 88494 52294
rect 87874 34614 88494 52058
rect 95788 45174 96108 45206
rect 95788 44938 95830 45174
rect 96066 44938 96108 45174
rect 95788 44854 96108 44938
rect 95788 44618 95830 44854
rect 96066 44618 96108 44854
rect 95788 44586 96108 44618
rect 126508 45174 126828 45206
rect 126508 44938 126550 45174
rect 126786 44938 126828 45174
rect 126508 44854 126828 44938
rect 126508 44618 126550 44854
rect 126786 44618 126828 44854
rect 126508 44586 126828 44618
rect 134434 45174 135054 62618
rect 134434 44938 134466 45174
rect 134702 44938 134786 45174
rect 135022 44938 135054 45174
rect 134434 44854 135054 44938
rect 134434 44618 134466 44854
rect 134702 44618 134786 44854
rect 135022 44618 135054 44854
rect 95128 41454 95448 41486
rect 95128 41218 95170 41454
rect 95406 41218 95448 41454
rect 95128 41134 95448 41218
rect 95128 40898 95170 41134
rect 95406 40898 95448 41134
rect 95128 40866 95448 40898
rect 125848 41454 126168 41486
rect 125848 41218 125890 41454
rect 126126 41218 126168 41454
rect 125848 41134 126168 41218
rect 125848 40898 125890 41134
rect 126126 40898 126168 41134
rect 125848 40866 126168 40898
rect 87874 34378 87906 34614
rect 88142 34378 88226 34614
rect 88462 34378 88494 34614
rect 87874 34294 88494 34378
rect 87874 34058 87906 34294
rect 88142 34058 88226 34294
rect 88462 34058 88494 34294
rect 87874 16614 88494 34058
rect 95788 27174 96108 27206
rect 95788 26938 95830 27174
rect 96066 26938 96108 27174
rect 95788 26854 96108 26938
rect 95788 26618 95830 26854
rect 96066 26618 96108 26854
rect 95788 26586 96108 26618
rect 134434 27174 135054 44618
rect 134434 26938 134466 27174
rect 134702 26938 134786 27174
rect 135022 26938 135054 27174
rect 134434 26854 135054 26938
rect 134434 26618 134466 26854
rect 134702 26618 134786 26854
rect 135022 26618 135054 26854
rect 95128 23454 95448 23486
rect 95128 23218 95170 23454
rect 95406 23218 95448 23454
rect 95128 23134 95448 23218
rect 95128 22898 95170 23134
rect 95406 22898 95448 23134
rect 95128 22866 95448 22898
rect 87874 16378 87906 16614
rect 88142 16378 88226 16614
rect 88462 16378 88494 16614
rect 87874 16294 88494 16378
rect 87874 16058 87906 16294
rect 88142 16058 88226 16294
rect 88462 16058 88494 16294
rect 87874 -3736 88494 16058
rect 87874 -3972 87906 -3736
rect 88142 -3972 88226 -3736
rect 88462 -3972 88494 -3736
rect 87874 -4056 88494 -3972
rect 87874 -4292 87906 -4056
rect 88142 -4292 88226 -4056
rect 88462 -4292 88494 -4056
rect 87874 -4324 88494 -4292
rect 94714 5454 95334 19988
rect 100339 19412 100405 19413
rect 100339 19348 100340 19412
rect 100404 19348 100405 19412
rect 100339 19347 100405 19348
rect 108435 19412 108501 19413
rect 108435 19348 108436 19412
rect 108500 19348 108501 19412
rect 108435 19347 108501 19348
rect 94714 5218 94746 5454
rect 94982 5218 95066 5454
rect 95302 5218 95334 5454
rect 94714 5134 95334 5218
rect 94714 4898 94746 5134
rect 94982 4898 95066 5134
rect 95302 4898 95334 5134
rect 94714 -856 95334 4898
rect 94714 -1092 94746 -856
rect 94982 -1092 95066 -856
rect 95302 -1092 95334 -856
rect 94714 -1176 95334 -1092
rect 94714 -1412 94746 -1176
rect 94982 -1412 95066 -1176
rect 95302 -1412 95334 -1176
rect 94714 -4324 95334 -1412
rect 98434 9174 99054 17955
rect 98434 8938 98466 9174
rect 98702 8938 98786 9174
rect 99022 8938 99054 9174
rect 98434 8854 99054 8938
rect 98434 8618 98466 8854
rect 98702 8618 98786 8854
rect 99022 8618 99054 8854
rect 98434 -1816 99054 8618
rect 100342 1138 100402 19347
rect 102154 12894 102774 17955
rect 102154 12658 102186 12894
rect 102422 12658 102506 12894
rect 102742 12658 102774 12894
rect 102154 12574 102774 12658
rect 102154 12338 102186 12574
rect 102422 12338 102506 12574
rect 102742 12338 102774 12574
rect 98434 -2052 98466 -1816
rect 98702 -2052 98786 -1816
rect 99022 -2052 99054 -1816
rect 98434 -2136 99054 -2052
rect 98434 -2372 98466 -2136
rect 98702 -2372 98786 -2136
rect 99022 -2372 99054 -2136
rect 98434 -4324 99054 -2372
rect 102154 -2776 102774 12338
rect 102154 -3012 102186 -2776
rect 102422 -3012 102506 -2776
rect 102742 -3012 102774 -2776
rect 102154 -3096 102774 -3012
rect 102154 -3332 102186 -3096
rect 102422 -3332 102506 -3096
rect 102742 -3332 102774 -3096
rect 102154 -4324 102774 -3332
rect 105874 16614 106494 17955
rect 105874 16378 105906 16614
rect 106142 16378 106226 16614
rect 106462 16378 106494 16614
rect 108438 16590 108498 19347
rect 108438 16530 109050 16590
rect 105874 16294 106494 16378
rect 105874 16058 105906 16294
rect 106142 16058 106226 16294
rect 106462 16058 106494 16294
rect 105874 -3736 106494 16058
rect 108990 1138 109050 16530
rect 112714 5454 113334 17955
rect 112714 5218 112746 5454
rect 112982 5218 113066 5454
rect 113302 5218 113334 5454
rect 112714 5134 113334 5218
rect 112714 4898 112746 5134
rect 112982 4898 113066 5134
rect 113302 4898 113334 5134
rect 105874 -3972 105906 -3736
rect 106142 -3972 106226 -3736
rect 106462 -3972 106494 -3736
rect 105874 -4056 106494 -3972
rect 105874 -4292 105906 -4056
rect 106142 -4292 106226 -4056
rect 106462 -4292 106494 -4056
rect 105874 -4324 106494 -4292
rect 112714 -856 113334 4898
rect 112714 -1092 112746 -856
rect 112982 -1092 113066 -856
rect 113302 -1092 113334 -856
rect 112714 -1176 113334 -1092
rect 112714 -1412 112746 -1176
rect 112982 -1412 113066 -1176
rect 113302 -1412 113334 -1176
rect 112714 -4324 113334 -1412
rect 116434 9174 117054 17955
rect 116434 8938 116466 9174
rect 116702 8938 116786 9174
rect 117022 8938 117054 9174
rect 116434 8854 117054 8938
rect 116434 8618 116466 8854
rect 116702 8618 116786 8854
rect 117022 8618 117054 8854
rect 116434 -1816 117054 8618
rect 116434 -2052 116466 -1816
rect 116702 -2052 116786 -1816
rect 117022 -2052 117054 -1816
rect 116434 -2136 117054 -2052
rect 116434 -2372 116466 -2136
rect 116702 -2372 116786 -2136
rect 117022 -2372 117054 -2136
rect 116434 -4324 117054 -2372
rect 120154 12894 120774 17955
rect 120154 12658 120186 12894
rect 120422 12658 120506 12894
rect 120742 12658 120774 12894
rect 120154 12574 120774 12658
rect 120154 12338 120186 12574
rect 120422 12338 120506 12574
rect 120742 12338 120774 12574
rect 120154 -2776 120774 12338
rect 120154 -3012 120186 -2776
rect 120422 -3012 120506 -2776
rect 120742 -3012 120774 -2776
rect 120154 -3096 120774 -3012
rect 120154 -3332 120186 -3096
rect 120422 -3332 120506 -3096
rect 120742 -3332 120774 -3096
rect 120154 -4324 120774 -3332
rect 123874 16614 124494 17955
rect 123874 16378 123906 16614
rect 124142 16378 124226 16614
rect 124462 16378 124494 16614
rect 123874 16294 124494 16378
rect 123874 16058 123906 16294
rect 124142 16058 124226 16294
rect 124462 16058 124494 16294
rect 123874 -3736 124494 16058
rect 123874 -3972 123906 -3736
rect 124142 -3972 124226 -3736
rect 124462 -3972 124494 -3736
rect 123874 -4056 124494 -3972
rect 123874 -4292 123906 -4056
rect 124142 -4292 124226 -4056
rect 124462 -4292 124494 -4056
rect 123874 -4324 124494 -4292
rect 130714 5454 131334 17955
rect 130714 5218 130746 5454
rect 130982 5218 131066 5454
rect 131302 5218 131334 5454
rect 130714 5134 131334 5218
rect 130714 4898 130746 5134
rect 130982 4898 131066 5134
rect 131302 4898 131334 5134
rect 130714 -856 131334 4898
rect 130714 -1092 130746 -856
rect 130982 -1092 131066 -856
rect 131302 -1092 131334 -856
rect 130714 -1176 131334 -1092
rect 130714 -1412 130746 -1176
rect 130982 -1412 131066 -1176
rect 131302 -1412 131334 -1176
rect 130714 -4324 131334 -1412
rect 134434 9174 135054 26618
rect 134434 8938 134466 9174
rect 134702 8938 134786 9174
rect 135022 8938 135054 9174
rect 134434 8854 135054 8938
rect 134434 8618 134466 8854
rect 134702 8618 134786 8854
rect 135022 8618 135054 8854
rect 134434 -1816 135054 8618
rect 138154 463012 138774 464004
rect 138154 462776 138186 463012
rect 138422 462776 138506 463012
rect 138742 462776 138774 463012
rect 138154 462692 138774 462776
rect 138154 462456 138186 462692
rect 138422 462456 138506 462692
rect 138742 462456 138774 462692
rect 138154 444894 138774 462456
rect 138154 444658 138186 444894
rect 138422 444658 138506 444894
rect 138742 444658 138774 444894
rect 138154 444574 138774 444658
rect 138154 444338 138186 444574
rect 138422 444338 138506 444574
rect 138742 444338 138774 444574
rect 138154 426894 138774 444338
rect 138154 426658 138186 426894
rect 138422 426658 138506 426894
rect 138742 426658 138774 426894
rect 138154 426574 138774 426658
rect 138154 426338 138186 426574
rect 138422 426338 138506 426574
rect 138742 426338 138774 426574
rect 138154 408894 138774 426338
rect 138154 408658 138186 408894
rect 138422 408658 138506 408894
rect 138742 408658 138774 408894
rect 138154 408574 138774 408658
rect 138154 408338 138186 408574
rect 138422 408338 138506 408574
rect 138742 408338 138774 408574
rect 138154 390894 138774 408338
rect 138154 390658 138186 390894
rect 138422 390658 138506 390894
rect 138742 390658 138774 390894
rect 138154 390574 138774 390658
rect 138154 390338 138186 390574
rect 138422 390338 138506 390574
rect 138742 390338 138774 390574
rect 138154 372894 138774 390338
rect 138154 372658 138186 372894
rect 138422 372658 138506 372894
rect 138742 372658 138774 372894
rect 138154 372574 138774 372658
rect 138154 372338 138186 372574
rect 138422 372338 138506 372574
rect 138742 372338 138774 372574
rect 138154 354894 138774 372338
rect 138154 354658 138186 354894
rect 138422 354658 138506 354894
rect 138742 354658 138774 354894
rect 138154 354574 138774 354658
rect 138154 354338 138186 354574
rect 138422 354338 138506 354574
rect 138742 354338 138774 354574
rect 138154 336894 138774 354338
rect 138154 336658 138186 336894
rect 138422 336658 138506 336894
rect 138742 336658 138774 336894
rect 138154 336574 138774 336658
rect 138154 336338 138186 336574
rect 138422 336338 138506 336574
rect 138742 336338 138774 336574
rect 138154 318894 138774 336338
rect 138154 318658 138186 318894
rect 138422 318658 138506 318894
rect 138742 318658 138774 318894
rect 138154 318574 138774 318658
rect 138154 318338 138186 318574
rect 138422 318338 138506 318574
rect 138742 318338 138774 318574
rect 138154 300894 138774 318338
rect 138154 300658 138186 300894
rect 138422 300658 138506 300894
rect 138742 300658 138774 300894
rect 138154 300574 138774 300658
rect 138154 300338 138186 300574
rect 138422 300338 138506 300574
rect 138742 300338 138774 300574
rect 138154 282894 138774 300338
rect 138154 282658 138186 282894
rect 138422 282658 138506 282894
rect 138742 282658 138774 282894
rect 138154 282574 138774 282658
rect 138154 282338 138186 282574
rect 138422 282338 138506 282574
rect 138742 282338 138774 282574
rect 138154 264894 138774 282338
rect 138154 264658 138186 264894
rect 138422 264658 138506 264894
rect 138742 264658 138774 264894
rect 138154 264574 138774 264658
rect 138154 264338 138186 264574
rect 138422 264338 138506 264574
rect 138742 264338 138774 264574
rect 138154 246894 138774 264338
rect 138154 246658 138186 246894
rect 138422 246658 138506 246894
rect 138742 246658 138774 246894
rect 138154 246574 138774 246658
rect 138154 246338 138186 246574
rect 138422 246338 138506 246574
rect 138742 246338 138774 246574
rect 138154 228894 138774 246338
rect 138154 228658 138186 228894
rect 138422 228658 138506 228894
rect 138742 228658 138774 228894
rect 138154 228574 138774 228658
rect 138154 228338 138186 228574
rect 138422 228338 138506 228574
rect 138742 228338 138774 228574
rect 138154 210894 138774 228338
rect 138154 210658 138186 210894
rect 138422 210658 138506 210894
rect 138742 210658 138774 210894
rect 138154 210574 138774 210658
rect 138154 210338 138186 210574
rect 138422 210338 138506 210574
rect 138742 210338 138774 210574
rect 138154 192894 138774 210338
rect 138154 192658 138186 192894
rect 138422 192658 138506 192894
rect 138742 192658 138774 192894
rect 138154 192574 138774 192658
rect 138154 192338 138186 192574
rect 138422 192338 138506 192574
rect 138742 192338 138774 192574
rect 138154 174894 138774 192338
rect 138154 174658 138186 174894
rect 138422 174658 138506 174894
rect 138742 174658 138774 174894
rect 138154 174574 138774 174658
rect 138154 174338 138186 174574
rect 138422 174338 138506 174574
rect 138742 174338 138774 174574
rect 138154 156894 138774 174338
rect 138154 156658 138186 156894
rect 138422 156658 138506 156894
rect 138742 156658 138774 156894
rect 138154 156574 138774 156658
rect 138154 156338 138186 156574
rect 138422 156338 138506 156574
rect 138742 156338 138774 156574
rect 138154 138894 138774 156338
rect 138154 138658 138186 138894
rect 138422 138658 138506 138894
rect 138742 138658 138774 138894
rect 138154 138574 138774 138658
rect 138154 138338 138186 138574
rect 138422 138338 138506 138574
rect 138742 138338 138774 138574
rect 138154 120894 138774 138338
rect 138154 120658 138186 120894
rect 138422 120658 138506 120894
rect 138742 120658 138774 120894
rect 138154 120574 138774 120658
rect 138154 120338 138186 120574
rect 138422 120338 138506 120574
rect 138742 120338 138774 120574
rect 138154 102894 138774 120338
rect 138154 102658 138186 102894
rect 138422 102658 138506 102894
rect 138742 102658 138774 102894
rect 138154 102574 138774 102658
rect 138154 102338 138186 102574
rect 138422 102338 138506 102574
rect 138742 102338 138774 102574
rect 138154 84894 138774 102338
rect 138154 84658 138186 84894
rect 138422 84658 138506 84894
rect 138742 84658 138774 84894
rect 138154 84574 138774 84658
rect 138154 84338 138186 84574
rect 138422 84338 138506 84574
rect 138742 84338 138774 84574
rect 138154 66894 138774 84338
rect 138154 66658 138186 66894
rect 138422 66658 138506 66894
rect 138742 66658 138774 66894
rect 138154 66574 138774 66658
rect 138154 66338 138186 66574
rect 138422 66338 138506 66574
rect 138742 66338 138774 66574
rect 138154 48894 138774 66338
rect 138154 48658 138186 48894
rect 138422 48658 138506 48894
rect 138742 48658 138774 48894
rect 138154 48574 138774 48658
rect 138154 48338 138186 48574
rect 138422 48338 138506 48574
rect 138742 48338 138774 48574
rect 138154 30894 138774 48338
rect 138154 30658 138186 30894
rect 138422 30658 138506 30894
rect 138742 30658 138774 30894
rect 138154 30574 138774 30658
rect 138154 30338 138186 30574
rect 138422 30338 138506 30574
rect 138742 30338 138774 30574
rect 138154 12894 138774 30338
rect 138154 12658 138186 12894
rect 138422 12658 138506 12894
rect 138742 12658 138774 12894
rect 138154 12574 138774 12658
rect 138154 12338 138186 12574
rect 138422 12338 138506 12574
rect 138742 12338 138774 12574
rect 137875 916 137941 917
rect 137875 852 137876 916
rect 137940 852 137941 916
rect 137875 851 137941 852
rect 137878 458 137938 851
rect 134434 -2052 134466 -1816
rect 134702 -2052 134786 -1816
rect 135022 -2052 135054 -1816
rect 134434 -2136 135054 -2052
rect 134434 -2372 134466 -2136
rect 134702 -2372 134786 -2136
rect 135022 -2372 135054 -2136
rect 134434 -4324 135054 -2372
rect 138154 -2776 138774 12338
rect 138154 -3012 138186 -2776
rect 138422 -3012 138506 -2776
rect 138742 -3012 138774 -2776
rect 138154 -3096 138774 -3012
rect 138154 -3332 138186 -3096
rect 138422 -3332 138506 -3096
rect 138742 -3332 138774 -3096
rect 138154 -4324 138774 -3332
rect 141874 463972 142494 464004
rect 141874 463736 141906 463972
rect 142142 463736 142226 463972
rect 142462 463736 142494 463972
rect 141874 463652 142494 463736
rect 141874 463416 141906 463652
rect 142142 463416 142226 463652
rect 142462 463416 142494 463652
rect 141874 448614 142494 463416
rect 141874 448378 141906 448614
rect 142142 448378 142226 448614
rect 142462 448378 142494 448614
rect 141874 448294 142494 448378
rect 141874 448058 141906 448294
rect 142142 448058 142226 448294
rect 142462 448058 142494 448294
rect 141874 430614 142494 448058
rect 141874 430378 141906 430614
rect 142142 430378 142226 430614
rect 142462 430378 142494 430614
rect 141874 430294 142494 430378
rect 141874 430058 141906 430294
rect 142142 430058 142226 430294
rect 142462 430058 142494 430294
rect 141874 412614 142494 430058
rect 141874 412378 141906 412614
rect 142142 412378 142226 412614
rect 142462 412378 142494 412614
rect 141874 412294 142494 412378
rect 141874 412058 141906 412294
rect 142142 412058 142226 412294
rect 142462 412058 142494 412294
rect 141874 394614 142494 412058
rect 141874 394378 141906 394614
rect 142142 394378 142226 394614
rect 142462 394378 142494 394614
rect 141874 394294 142494 394378
rect 141874 394058 141906 394294
rect 142142 394058 142226 394294
rect 142462 394058 142494 394294
rect 141874 376614 142494 394058
rect 141874 376378 141906 376614
rect 142142 376378 142226 376614
rect 142462 376378 142494 376614
rect 141874 376294 142494 376378
rect 141874 376058 141906 376294
rect 142142 376058 142226 376294
rect 142462 376058 142494 376294
rect 141874 358614 142494 376058
rect 141874 358378 141906 358614
rect 142142 358378 142226 358614
rect 142462 358378 142494 358614
rect 141874 358294 142494 358378
rect 141874 358058 141906 358294
rect 142142 358058 142226 358294
rect 142462 358058 142494 358294
rect 141874 340614 142494 358058
rect 141874 340378 141906 340614
rect 142142 340378 142226 340614
rect 142462 340378 142494 340614
rect 141874 340294 142494 340378
rect 141874 340058 141906 340294
rect 142142 340058 142226 340294
rect 142462 340058 142494 340294
rect 141874 322614 142494 340058
rect 141874 322378 141906 322614
rect 142142 322378 142226 322614
rect 142462 322378 142494 322614
rect 141874 322294 142494 322378
rect 141874 322058 141906 322294
rect 142142 322058 142226 322294
rect 142462 322058 142494 322294
rect 141874 304614 142494 322058
rect 141874 304378 141906 304614
rect 142142 304378 142226 304614
rect 142462 304378 142494 304614
rect 141874 304294 142494 304378
rect 141874 304058 141906 304294
rect 142142 304058 142226 304294
rect 142462 304058 142494 304294
rect 141874 286614 142494 304058
rect 141874 286378 141906 286614
rect 142142 286378 142226 286614
rect 142462 286378 142494 286614
rect 141874 286294 142494 286378
rect 141874 286058 141906 286294
rect 142142 286058 142226 286294
rect 142462 286058 142494 286294
rect 141874 268614 142494 286058
rect 141874 268378 141906 268614
rect 142142 268378 142226 268614
rect 142462 268378 142494 268614
rect 141874 268294 142494 268378
rect 141874 268058 141906 268294
rect 142142 268058 142226 268294
rect 142462 268058 142494 268294
rect 141874 250614 142494 268058
rect 141874 250378 141906 250614
rect 142142 250378 142226 250614
rect 142462 250378 142494 250614
rect 141874 250294 142494 250378
rect 141874 250058 141906 250294
rect 142142 250058 142226 250294
rect 142462 250058 142494 250294
rect 141874 232614 142494 250058
rect 141874 232378 141906 232614
rect 142142 232378 142226 232614
rect 142462 232378 142494 232614
rect 141874 232294 142494 232378
rect 141874 232058 141906 232294
rect 142142 232058 142226 232294
rect 142462 232058 142494 232294
rect 141874 214614 142494 232058
rect 141874 214378 141906 214614
rect 142142 214378 142226 214614
rect 142462 214378 142494 214614
rect 141874 214294 142494 214378
rect 141874 214058 141906 214294
rect 142142 214058 142226 214294
rect 142462 214058 142494 214294
rect 141874 196614 142494 214058
rect 141874 196378 141906 196614
rect 142142 196378 142226 196614
rect 142462 196378 142494 196614
rect 141874 196294 142494 196378
rect 141874 196058 141906 196294
rect 142142 196058 142226 196294
rect 142462 196058 142494 196294
rect 141874 178614 142494 196058
rect 141874 178378 141906 178614
rect 142142 178378 142226 178614
rect 142462 178378 142494 178614
rect 141874 178294 142494 178378
rect 141874 178058 141906 178294
rect 142142 178058 142226 178294
rect 142462 178058 142494 178294
rect 141874 160614 142494 178058
rect 141874 160378 141906 160614
rect 142142 160378 142226 160614
rect 142462 160378 142494 160614
rect 141874 160294 142494 160378
rect 141874 160058 141906 160294
rect 142142 160058 142226 160294
rect 142462 160058 142494 160294
rect 141874 142614 142494 160058
rect 141874 142378 141906 142614
rect 142142 142378 142226 142614
rect 142462 142378 142494 142614
rect 141874 142294 142494 142378
rect 141874 142058 141906 142294
rect 142142 142058 142226 142294
rect 142462 142058 142494 142294
rect 141874 124614 142494 142058
rect 141874 124378 141906 124614
rect 142142 124378 142226 124614
rect 142462 124378 142494 124614
rect 141874 124294 142494 124378
rect 141874 124058 141906 124294
rect 142142 124058 142226 124294
rect 142462 124058 142494 124294
rect 141874 106614 142494 124058
rect 141874 106378 141906 106614
rect 142142 106378 142226 106614
rect 142462 106378 142494 106614
rect 141874 106294 142494 106378
rect 141874 106058 141906 106294
rect 142142 106058 142226 106294
rect 142462 106058 142494 106294
rect 141874 88614 142494 106058
rect 141874 88378 141906 88614
rect 142142 88378 142226 88614
rect 142462 88378 142494 88614
rect 141874 88294 142494 88378
rect 141874 88058 141906 88294
rect 142142 88058 142226 88294
rect 142462 88058 142494 88294
rect 141874 70614 142494 88058
rect 141874 70378 141906 70614
rect 142142 70378 142226 70614
rect 142462 70378 142494 70614
rect 141874 70294 142494 70378
rect 141874 70058 141906 70294
rect 142142 70058 142226 70294
rect 142462 70058 142494 70294
rect 141874 52614 142494 70058
rect 141874 52378 141906 52614
rect 142142 52378 142226 52614
rect 142462 52378 142494 52614
rect 141874 52294 142494 52378
rect 141874 52058 141906 52294
rect 142142 52058 142226 52294
rect 142462 52058 142494 52294
rect 141874 34614 142494 52058
rect 141874 34378 141906 34614
rect 142142 34378 142226 34614
rect 142462 34378 142494 34614
rect 141874 34294 142494 34378
rect 141874 34058 141906 34294
rect 142142 34058 142226 34294
rect 142462 34058 142494 34294
rect 141874 16614 142494 34058
rect 141874 16378 141906 16614
rect 142142 16378 142226 16614
rect 142462 16378 142494 16614
rect 141874 16294 142494 16378
rect 141874 16058 141906 16294
rect 142142 16058 142226 16294
rect 142462 16058 142494 16294
rect 141874 -3736 142494 16058
rect 141874 -3972 141906 -3736
rect 142142 -3972 142226 -3736
rect 142462 -3972 142494 -3736
rect 141874 -4056 142494 -3972
rect 141874 -4292 141906 -4056
rect 142142 -4292 142226 -4056
rect 142462 -4292 142494 -4056
rect 141874 -4324 142494 -4292
rect 148714 461092 149334 464004
rect 148714 460856 148746 461092
rect 148982 460856 149066 461092
rect 149302 460856 149334 461092
rect 148714 460772 149334 460856
rect 148714 460536 148746 460772
rect 148982 460536 149066 460772
rect 149302 460536 149334 460772
rect 148714 455454 149334 460536
rect 148714 455218 148746 455454
rect 148982 455218 149066 455454
rect 149302 455218 149334 455454
rect 148714 455134 149334 455218
rect 148714 454898 148746 455134
rect 148982 454898 149066 455134
rect 149302 454898 149334 455134
rect 148714 437454 149334 454898
rect 148714 437218 148746 437454
rect 148982 437218 149066 437454
rect 149302 437218 149334 437454
rect 148714 437134 149334 437218
rect 148714 436898 148746 437134
rect 148982 436898 149066 437134
rect 149302 436898 149334 437134
rect 148714 419454 149334 436898
rect 148714 419218 148746 419454
rect 148982 419218 149066 419454
rect 149302 419218 149334 419454
rect 148714 419134 149334 419218
rect 148714 418898 148746 419134
rect 148982 418898 149066 419134
rect 149302 418898 149334 419134
rect 148714 401454 149334 418898
rect 148714 401218 148746 401454
rect 148982 401218 149066 401454
rect 149302 401218 149334 401454
rect 148714 401134 149334 401218
rect 148714 400898 148746 401134
rect 148982 400898 149066 401134
rect 149302 400898 149334 401134
rect 148714 383454 149334 400898
rect 148714 383218 148746 383454
rect 148982 383218 149066 383454
rect 149302 383218 149334 383454
rect 148714 383134 149334 383218
rect 148714 382898 148746 383134
rect 148982 382898 149066 383134
rect 149302 382898 149334 383134
rect 148714 365454 149334 382898
rect 148714 365218 148746 365454
rect 148982 365218 149066 365454
rect 149302 365218 149334 365454
rect 148714 365134 149334 365218
rect 148714 364898 148746 365134
rect 148982 364898 149066 365134
rect 149302 364898 149334 365134
rect 148714 347454 149334 364898
rect 148714 347218 148746 347454
rect 148982 347218 149066 347454
rect 149302 347218 149334 347454
rect 148714 347134 149334 347218
rect 148714 346898 148746 347134
rect 148982 346898 149066 347134
rect 149302 346898 149334 347134
rect 148714 329454 149334 346898
rect 148714 329218 148746 329454
rect 148982 329218 149066 329454
rect 149302 329218 149334 329454
rect 148714 329134 149334 329218
rect 148714 328898 148746 329134
rect 148982 328898 149066 329134
rect 149302 328898 149334 329134
rect 148714 311454 149334 328898
rect 148714 311218 148746 311454
rect 148982 311218 149066 311454
rect 149302 311218 149334 311454
rect 148714 311134 149334 311218
rect 148714 310898 148746 311134
rect 148982 310898 149066 311134
rect 149302 310898 149334 311134
rect 148714 293454 149334 310898
rect 148714 293218 148746 293454
rect 148982 293218 149066 293454
rect 149302 293218 149334 293454
rect 148714 293134 149334 293218
rect 148714 292898 148746 293134
rect 148982 292898 149066 293134
rect 149302 292898 149334 293134
rect 148714 275454 149334 292898
rect 148714 275218 148746 275454
rect 148982 275218 149066 275454
rect 149302 275218 149334 275454
rect 148714 275134 149334 275218
rect 148714 274898 148746 275134
rect 148982 274898 149066 275134
rect 149302 274898 149334 275134
rect 148714 257454 149334 274898
rect 148714 257218 148746 257454
rect 148982 257218 149066 257454
rect 149302 257218 149334 257454
rect 148714 257134 149334 257218
rect 148714 256898 148746 257134
rect 148982 256898 149066 257134
rect 149302 256898 149334 257134
rect 148714 239454 149334 256898
rect 148714 239218 148746 239454
rect 148982 239218 149066 239454
rect 149302 239218 149334 239454
rect 148714 239134 149334 239218
rect 148714 238898 148746 239134
rect 148982 238898 149066 239134
rect 149302 238898 149334 239134
rect 148714 221454 149334 238898
rect 148714 221218 148746 221454
rect 148982 221218 149066 221454
rect 149302 221218 149334 221454
rect 148714 221134 149334 221218
rect 148714 220898 148746 221134
rect 148982 220898 149066 221134
rect 149302 220898 149334 221134
rect 148714 203454 149334 220898
rect 148714 203218 148746 203454
rect 148982 203218 149066 203454
rect 149302 203218 149334 203454
rect 148714 203134 149334 203218
rect 148714 202898 148746 203134
rect 148982 202898 149066 203134
rect 149302 202898 149334 203134
rect 148714 185454 149334 202898
rect 148714 185218 148746 185454
rect 148982 185218 149066 185454
rect 149302 185218 149334 185454
rect 148714 185134 149334 185218
rect 148714 184898 148746 185134
rect 148982 184898 149066 185134
rect 149302 184898 149334 185134
rect 148714 167454 149334 184898
rect 148714 167218 148746 167454
rect 148982 167218 149066 167454
rect 149302 167218 149334 167454
rect 148714 167134 149334 167218
rect 148714 166898 148746 167134
rect 148982 166898 149066 167134
rect 149302 166898 149334 167134
rect 148714 149454 149334 166898
rect 148714 149218 148746 149454
rect 148982 149218 149066 149454
rect 149302 149218 149334 149454
rect 148714 149134 149334 149218
rect 148714 148898 148746 149134
rect 148982 148898 149066 149134
rect 149302 148898 149334 149134
rect 148714 131454 149334 148898
rect 148714 131218 148746 131454
rect 148982 131218 149066 131454
rect 149302 131218 149334 131454
rect 148714 131134 149334 131218
rect 148714 130898 148746 131134
rect 148982 130898 149066 131134
rect 149302 130898 149334 131134
rect 148714 113454 149334 130898
rect 148714 113218 148746 113454
rect 148982 113218 149066 113454
rect 149302 113218 149334 113454
rect 148714 113134 149334 113218
rect 148714 112898 148746 113134
rect 148982 112898 149066 113134
rect 149302 112898 149334 113134
rect 148714 95454 149334 112898
rect 148714 95218 148746 95454
rect 148982 95218 149066 95454
rect 149302 95218 149334 95454
rect 148714 95134 149334 95218
rect 148714 94898 148746 95134
rect 148982 94898 149066 95134
rect 149302 94898 149334 95134
rect 148714 77454 149334 94898
rect 148714 77218 148746 77454
rect 148982 77218 149066 77454
rect 149302 77218 149334 77454
rect 148714 77134 149334 77218
rect 148714 76898 148746 77134
rect 148982 76898 149066 77134
rect 149302 76898 149334 77134
rect 148714 59454 149334 76898
rect 148714 59218 148746 59454
rect 148982 59218 149066 59454
rect 149302 59218 149334 59454
rect 148714 59134 149334 59218
rect 148714 58898 148746 59134
rect 148982 58898 149066 59134
rect 149302 58898 149334 59134
rect 148714 41454 149334 58898
rect 148714 41218 148746 41454
rect 148982 41218 149066 41454
rect 149302 41218 149334 41454
rect 148714 41134 149334 41218
rect 148714 40898 148746 41134
rect 148982 40898 149066 41134
rect 149302 40898 149334 41134
rect 148714 23454 149334 40898
rect 148714 23218 148746 23454
rect 148982 23218 149066 23454
rect 149302 23218 149334 23454
rect 148714 23134 149334 23218
rect 148714 22898 148746 23134
rect 148982 22898 149066 23134
rect 149302 22898 149334 23134
rect 148714 5454 149334 22898
rect 152434 462052 153054 464004
rect 152434 461816 152466 462052
rect 152702 461816 152786 462052
rect 153022 461816 153054 462052
rect 152434 461732 153054 461816
rect 152434 461496 152466 461732
rect 152702 461496 152786 461732
rect 153022 461496 153054 461732
rect 152434 441174 153054 461496
rect 152434 440938 152466 441174
rect 152702 440938 152786 441174
rect 153022 440938 153054 441174
rect 152434 440854 153054 440938
rect 152434 440618 152466 440854
rect 152702 440618 152786 440854
rect 153022 440618 153054 440854
rect 152434 423174 153054 440618
rect 152434 422938 152466 423174
rect 152702 422938 152786 423174
rect 153022 422938 153054 423174
rect 152434 422854 153054 422938
rect 152434 422618 152466 422854
rect 152702 422618 152786 422854
rect 153022 422618 153054 422854
rect 152434 405174 153054 422618
rect 152434 404938 152466 405174
rect 152702 404938 152786 405174
rect 153022 404938 153054 405174
rect 152434 404854 153054 404938
rect 152434 404618 152466 404854
rect 152702 404618 152786 404854
rect 153022 404618 153054 404854
rect 152434 387174 153054 404618
rect 152434 386938 152466 387174
rect 152702 386938 152786 387174
rect 153022 386938 153054 387174
rect 152434 386854 153054 386938
rect 152434 386618 152466 386854
rect 152702 386618 152786 386854
rect 153022 386618 153054 386854
rect 152434 369174 153054 386618
rect 152434 368938 152466 369174
rect 152702 368938 152786 369174
rect 153022 368938 153054 369174
rect 152434 368854 153054 368938
rect 152434 368618 152466 368854
rect 152702 368618 152786 368854
rect 153022 368618 153054 368854
rect 152434 351174 153054 368618
rect 152434 350938 152466 351174
rect 152702 350938 152786 351174
rect 153022 350938 153054 351174
rect 152434 350854 153054 350938
rect 152434 350618 152466 350854
rect 152702 350618 152786 350854
rect 153022 350618 153054 350854
rect 152434 333174 153054 350618
rect 152434 332938 152466 333174
rect 152702 332938 152786 333174
rect 153022 332938 153054 333174
rect 152434 332854 153054 332938
rect 152434 332618 152466 332854
rect 152702 332618 152786 332854
rect 153022 332618 153054 332854
rect 152434 315174 153054 332618
rect 152434 314938 152466 315174
rect 152702 314938 152786 315174
rect 153022 314938 153054 315174
rect 152434 314854 153054 314938
rect 152434 314618 152466 314854
rect 152702 314618 152786 314854
rect 153022 314618 153054 314854
rect 152434 297174 153054 314618
rect 152434 296938 152466 297174
rect 152702 296938 152786 297174
rect 153022 296938 153054 297174
rect 152434 296854 153054 296938
rect 152434 296618 152466 296854
rect 152702 296618 152786 296854
rect 153022 296618 153054 296854
rect 152434 279174 153054 296618
rect 152434 278938 152466 279174
rect 152702 278938 152786 279174
rect 153022 278938 153054 279174
rect 152434 278854 153054 278938
rect 152434 278618 152466 278854
rect 152702 278618 152786 278854
rect 153022 278618 153054 278854
rect 152434 261174 153054 278618
rect 152434 260938 152466 261174
rect 152702 260938 152786 261174
rect 153022 260938 153054 261174
rect 152434 260854 153054 260938
rect 152434 260618 152466 260854
rect 152702 260618 152786 260854
rect 153022 260618 153054 260854
rect 152434 243174 153054 260618
rect 152434 242938 152466 243174
rect 152702 242938 152786 243174
rect 153022 242938 153054 243174
rect 152434 242854 153054 242938
rect 152434 242618 152466 242854
rect 152702 242618 152786 242854
rect 153022 242618 153054 242854
rect 152434 225174 153054 242618
rect 152434 224938 152466 225174
rect 152702 224938 152786 225174
rect 153022 224938 153054 225174
rect 152434 224854 153054 224938
rect 152434 224618 152466 224854
rect 152702 224618 152786 224854
rect 153022 224618 153054 224854
rect 152434 207174 153054 224618
rect 152434 206938 152466 207174
rect 152702 206938 152786 207174
rect 153022 206938 153054 207174
rect 152434 206854 153054 206938
rect 152434 206618 152466 206854
rect 152702 206618 152786 206854
rect 153022 206618 153054 206854
rect 152434 189174 153054 206618
rect 152434 188938 152466 189174
rect 152702 188938 152786 189174
rect 153022 188938 153054 189174
rect 152434 188854 153054 188938
rect 152434 188618 152466 188854
rect 152702 188618 152786 188854
rect 153022 188618 153054 188854
rect 152434 171174 153054 188618
rect 152434 170938 152466 171174
rect 152702 170938 152786 171174
rect 153022 170938 153054 171174
rect 152434 170854 153054 170938
rect 152434 170618 152466 170854
rect 152702 170618 152786 170854
rect 153022 170618 153054 170854
rect 152434 153174 153054 170618
rect 152434 152938 152466 153174
rect 152702 152938 152786 153174
rect 153022 152938 153054 153174
rect 152434 152854 153054 152938
rect 152434 152618 152466 152854
rect 152702 152618 152786 152854
rect 153022 152618 153054 152854
rect 152434 135174 153054 152618
rect 152434 134938 152466 135174
rect 152702 134938 152786 135174
rect 153022 134938 153054 135174
rect 152434 134854 153054 134938
rect 152434 134618 152466 134854
rect 152702 134618 152786 134854
rect 153022 134618 153054 134854
rect 152434 117174 153054 134618
rect 152434 116938 152466 117174
rect 152702 116938 152786 117174
rect 153022 116938 153054 117174
rect 152434 116854 153054 116938
rect 152434 116618 152466 116854
rect 152702 116618 152786 116854
rect 153022 116618 153054 116854
rect 152434 99174 153054 116618
rect 152434 98938 152466 99174
rect 152702 98938 152786 99174
rect 153022 98938 153054 99174
rect 152434 98854 153054 98938
rect 152434 98618 152466 98854
rect 152702 98618 152786 98854
rect 153022 98618 153054 98854
rect 152434 81174 153054 98618
rect 152434 80938 152466 81174
rect 152702 80938 152786 81174
rect 153022 80938 153054 81174
rect 152434 80854 153054 80938
rect 152434 80618 152466 80854
rect 152702 80618 152786 80854
rect 153022 80618 153054 80854
rect 152434 63174 153054 80618
rect 152434 62938 152466 63174
rect 152702 62938 152786 63174
rect 153022 62938 153054 63174
rect 152434 62854 153054 62938
rect 152434 62618 152466 62854
rect 152702 62618 152786 62854
rect 153022 62618 153054 62854
rect 152434 45174 153054 62618
rect 156154 463012 156774 464004
rect 156154 462776 156186 463012
rect 156422 462776 156506 463012
rect 156742 462776 156774 463012
rect 156154 462692 156774 462776
rect 156154 462456 156186 462692
rect 156422 462456 156506 462692
rect 156742 462456 156774 462692
rect 156154 444894 156774 462456
rect 156154 444658 156186 444894
rect 156422 444658 156506 444894
rect 156742 444658 156774 444894
rect 156154 444574 156774 444658
rect 156154 444338 156186 444574
rect 156422 444338 156506 444574
rect 156742 444338 156774 444574
rect 156154 426894 156774 444338
rect 156154 426658 156186 426894
rect 156422 426658 156506 426894
rect 156742 426658 156774 426894
rect 156154 426574 156774 426658
rect 156154 426338 156186 426574
rect 156422 426338 156506 426574
rect 156742 426338 156774 426574
rect 156154 408894 156774 426338
rect 156154 408658 156186 408894
rect 156422 408658 156506 408894
rect 156742 408658 156774 408894
rect 156154 408574 156774 408658
rect 156154 408338 156186 408574
rect 156422 408338 156506 408574
rect 156742 408338 156774 408574
rect 156154 390894 156774 408338
rect 156154 390658 156186 390894
rect 156422 390658 156506 390894
rect 156742 390658 156774 390894
rect 156154 390574 156774 390658
rect 156154 390338 156186 390574
rect 156422 390338 156506 390574
rect 156742 390338 156774 390574
rect 156154 372894 156774 390338
rect 156154 372658 156186 372894
rect 156422 372658 156506 372894
rect 156742 372658 156774 372894
rect 156154 372574 156774 372658
rect 156154 372338 156186 372574
rect 156422 372338 156506 372574
rect 156742 372338 156774 372574
rect 156154 354894 156774 372338
rect 156154 354658 156186 354894
rect 156422 354658 156506 354894
rect 156742 354658 156774 354894
rect 156154 354574 156774 354658
rect 156154 354338 156186 354574
rect 156422 354338 156506 354574
rect 156742 354338 156774 354574
rect 156154 336894 156774 354338
rect 156154 336658 156186 336894
rect 156422 336658 156506 336894
rect 156742 336658 156774 336894
rect 156154 336574 156774 336658
rect 156154 336338 156186 336574
rect 156422 336338 156506 336574
rect 156742 336338 156774 336574
rect 156154 318894 156774 336338
rect 156154 318658 156186 318894
rect 156422 318658 156506 318894
rect 156742 318658 156774 318894
rect 156154 318574 156774 318658
rect 156154 318338 156186 318574
rect 156422 318338 156506 318574
rect 156742 318338 156774 318574
rect 156154 300894 156774 318338
rect 156154 300658 156186 300894
rect 156422 300658 156506 300894
rect 156742 300658 156774 300894
rect 156154 300574 156774 300658
rect 156154 300338 156186 300574
rect 156422 300338 156506 300574
rect 156742 300338 156774 300574
rect 156154 282894 156774 300338
rect 156154 282658 156186 282894
rect 156422 282658 156506 282894
rect 156742 282658 156774 282894
rect 156154 282574 156774 282658
rect 156154 282338 156186 282574
rect 156422 282338 156506 282574
rect 156742 282338 156774 282574
rect 156154 264894 156774 282338
rect 156154 264658 156186 264894
rect 156422 264658 156506 264894
rect 156742 264658 156774 264894
rect 156154 264574 156774 264658
rect 156154 264338 156186 264574
rect 156422 264338 156506 264574
rect 156742 264338 156774 264574
rect 156154 246894 156774 264338
rect 156154 246658 156186 246894
rect 156422 246658 156506 246894
rect 156742 246658 156774 246894
rect 156154 246574 156774 246658
rect 156154 246338 156186 246574
rect 156422 246338 156506 246574
rect 156742 246338 156774 246574
rect 156154 228894 156774 246338
rect 156154 228658 156186 228894
rect 156422 228658 156506 228894
rect 156742 228658 156774 228894
rect 156154 228574 156774 228658
rect 156154 228338 156186 228574
rect 156422 228338 156506 228574
rect 156742 228338 156774 228574
rect 156154 210894 156774 228338
rect 156154 210658 156186 210894
rect 156422 210658 156506 210894
rect 156742 210658 156774 210894
rect 156154 210574 156774 210658
rect 156154 210338 156186 210574
rect 156422 210338 156506 210574
rect 156742 210338 156774 210574
rect 156154 192894 156774 210338
rect 156154 192658 156186 192894
rect 156422 192658 156506 192894
rect 156742 192658 156774 192894
rect 156154 192574 156774 192658
rect 156154 192338 156186 192574
rect 156422 192338 156506 192574
rect 156742 192338 156774 192574
rect 156154 174894 156774 192338
rect 156154 174658 156186 174894
rect 156422 174658 156506 174894
rect 156742 174658 156774 174894
rect 156154 174574 156774 174658
rect 156154 174338 156186 174574
rect 156422 174338 156506 174574
rect 156742 174338 156774 174574
rect 156154 156894 156774 174338
rect 156154 156658 156186 156894
rect 156422 156658 156506 156894
rect 156742 156658 156774 156894
rect 156154 156574 156774 156658
rect 156154 156338 156186 156574
rect 156422 156338 156506 156574
rect 156742 156338 156774 156574
rect 156154 138894 156774 156338
rect 156154 138658 156186 138894
rect 156422 138658 156506 138894
rect 156742 138658 156774 138894
rect 156154 138574 156774 138658
rect 156154 138338 156186 138574
rect 156422 138338 156506 138574
rect 156742 138338 156774 138574
rect 156154 120894 156774 138338
rect 156154 120658 156186 120894
rect 156422 120658 156506 120894
rect 156742 120658 156774 120894
rect 156154 120574 156774 120658
rect 156154 120338 156186 120574
rect 156422 120338 156506 120574
rect 156742 120338 156774 120574
rect 156154 102894 156774 120338
rect 156154 102658 156186 102894
rect 156422 102658 156506 102894
rect 156742 102658 156774 102894
rect 156154 102574 156774 102658
rect 156154 102338 156186 102574
rect 156422 102338 156506 102574
rect 156742 102338 156774 102574
rect 156154 84894 156774 102338
rect 156154 84658 156186 84894
rect 156422 84658 156506 84894
rect 156742 84658 156774 84894
rect 156154 84574 156774 84658
rect 156154 84338 156186 84574
rect 156422 84338 156506 84574
rect 156742 84338 156774 84574
rect 156154 66894 156774 84338
rect 156154 66658 156186 66894
rect 156422 66658 156506 66894
rect 156742 66658 156774 66894
rect 156154 66574 156774 66658
rect 156154 66338 156186 66574
rect 156422 66338 156506 66574
rect 156742 66338 156774 66574
rect 156154 59724 156774 66338
rect 159874 463972 160494 464004
rect 159874 463736 159906 463972
rect 160142 463736 160226 463972
rect 160462 463736 160494 463972
rect 159874 463652 160494 463736
rect 159874 463416 159906 463652
rect 160142 463416 160226 463652
rect 160462 463416 160494 463652
rect 159874 448614 160494 463416
rect 159874 448378 159906 448614
rect 160142 448378 160226 448614
rect 160462 448378 160494 448614
rect 159874 448294 160494 448378
rect 159874 448058 159906 448294
rect 160142 448058 160226 448294
rect 160462 448058 160494 448294
rect 159874 430614 160494 448058
rect 159874 430378 159906 430614
rect 160142 430378 160226 430614
rect 160462 430378 160494 430614
rect 159874 430294 160494 430378
rect 159874 430058 159906 430294
rect 160142 430058 160226 430294
rect 160462 430058 160494 430294
rect 159874 412614 160494 430058
rect 159874 412378 159906 412614
rect 160142 412378 160226 412614
rect 160462 412378 160494 412614
rect 159874 412294 160494 412378
rect 159874 412058 159906 412294
rect 160142 412058 160226 412294
rect 160462 412058 160494 412294
rect 159874 394614 160494 412058
rect 159874 394378 159906 394614
rect 160142 394378 160226 394614
rect 160462 394378 160494 394614
rect 159874 394294 160494 394378
rect 159874 394058 159906 394294
rect 160142 394058 160226 394294
rect 160462 394058 160494 394294
rect 159874 376614 160494 394058
rect 159874 376378 159906 376614
rect 160142 376378 160226 376614
rect 160462 376378 160494 376614
rect 159874 376294 160494 376378
rect 159874 376058 159906 376294
rect 160142 376058 160226 376294
rect 160462 376058 160494 376294
rect 159874 358614 160494 376058
rect 159874 358378 159906 358614
rect 160142 358378 160226 358614
rect 160462 358378 160494 358614
rect 159874 358294 160494 358378
rect 159874 358058 159906 358294
rect 160142 358058 160226 358294
rect 160462 358058 160494 358294
rect 159874 340614 160494 358058
rect 159874 340378 159906 340614
rect 160142 340378 160226 340614
rect 160462 340378 160494 340614
rect 159874 340294 160494 340378
rect 159874 340058 159906 340294
rect 160142 340058 160226 340294
rect 160462 340058 160494 340294
rect 159874 322614 160494 340058
rect 159874 322378 159906 322614
rect 160142 322378 160226 322614
rect 160462 322378 160494 322614
rect 159874 322294 160494 322378
rect 159874 322058 159906 322294
rect 160142 322058 160226 322294
rect 160462 322058 160494 322294
rect 159874 304614 160494 322058
rect 159874 304378 159906 304614
rect 160142 304378 160226 304614
rect 160462 304378 160494 304614
rect 159874 304294 160494 304378
rect 159874 304058 159906 304294
rect 160142 304058 160226 304294
rect 160462 304058 160494 304294
rect 159874 286614 160494 304058
rect 159874 286378 159906 286614
rect 160142 286378 160226 286614
rect 160462 286378 160494 286614
rect 159874 286294 160494 286378
rect 159874 286058 159906 286294
rect 160142 286058 160226 286294
rect 160462 286058 160494 286294
rect 159874 268614 160494 286058
rect 159874 268378 159906 268614
rect 160142 268378 160226 268614
rect 160462 268378 160494 268614
rect 159874 268294 160494 268378
rect 159874 268058 159906 268294
rect 160142 268058 160226 268294
rect 160462 268058 160494 268294
rect 159874 250614 160494 268058
rect 159874 250378 159906 250614
rect 160142 250378 160226 250614
rect 160462 250378 160494 250614
rect 159874 250294 160494 250378
rect 159874 250058 159906 250294
rect 160142 250058 160226 250294
rect 160462 250058 160494 250294
rect 159874 232614 160494 250058
rect 159874 232378 159906 232614
rect 160142 232378 160226 232614
rect 160462 232378 160494 232614
rect 159874 232294 160494 232378
rect 159874 232058 159906 232294
rect 160142 232058 160226 232294
rect 160462 232058 160494 232294
rect 159874 214614 160494 232058
rect 159874 214378 159906 214614
rect 160142 214378 160226 214614
rect 160462 214378 160494 214614
rect 159874 214294 160494 214378
rect 159874 214058 159906 214294
rect 160142 214058 160226 214294
rect 160462 214058 160494 214294
rect 159874 196614 160494 214058
rect 159874 196378 159906 196614
rect 160142 196378 160226 196614
rect 160462 196378 160494 196614
rect 159874 196294 160494 196378
rect 159874 196058 159906 196294
rect 160142 196058 160226 196294
rect 160462 196058 160494 196294
rect 159874 178614 160494 196058
rect 159874 178378 159906 178614
rect 160142 178378 160226 178614
rect 160462 178378 160494 178614
rect 159874 178294 160494 178378
rect 159874 178058 159906 178294
rect 160142 178058 160226 178294
rect 160462 178058 160494 178294
rect 159874 160614 160494 178058
rect 159874 160378 159906 160614
rect 160142 160378 160226 160614
rect 160462 160378 160494 160614
rect 159874 160294 160494 160378
rect 159874 160058 159906 160294
rect 160142 160058 160226 160294
rect 160462 160058 160494 160294
rect 159874 142614 160494 160058
rect 159874 142378 159906 142614
rect 160142 142378 160226 142614
rect 160462 142378 160494 142614
rect 159874 142294 160494 142378
rect 159874 142058 159906 142294
rect 160142 142058 160226 142294
rect 160462 142058 160494 142294
rect 159874 124614 160494 142058
rect 159874 124378 159906 124614
rect 160142 124378 160226 124614
rect 160462 124378 160494 124614
rect 159874 124294 160494 124378
rect 159874 124058 159906 124294
rect 160142 124058 160226 124294
rect 160462 124058 160494 124294
rect 159874 106614 160494 124058
rect 159874 106378 159906 106614
rect 160142 106378 160226 106614
rect 160462 106378 160494 106614
rect 159874 106294 160494 106378
rect 159874 106058 159906 106294
rect 160142 106058 160226 106294
rect 160462 106058 160494 106294
rect 159874 88614 160494 106058
rect 159874 88378 159906 88614
rect 160142 88378 160226 88614
rect 160462 88378 160494 88614
rect 159874 88294 160494 88378
rect 159874 88058 159906 88294
rect 160142 88058 160226 88294
rect 160462 88058 160494 88294
rect 159874 70614 160494 88058
rect 159874 70378 159906 70614
rect 160142 70378 160226 70614
rect 160462 70378 160494 70614
rect 159874 70294 160494 70378
rect 159874 70058 159906 70294
rect 160142 70058 160226 70294
rect 160462 70058 160494 70294
rect 159874 52614 160494 70058
rect 159874 52378 159906 52614
rect 160142 52378 160226 52614
rect 160462 52378 160494 52614
rect 159874 52294 160494 52378
rect 159874 52058 159906 52294
rect 160142 52058 160226 52294
rect 160462 52058 160494 52294
rect 152434 44938 152466 45174
rect 152702 44938 152786 45174
rect 153022 44938 153054 45174
rect 152434 44854 153054 44938
rect 152434 44618 152466 44854
rect 152702 44618 152786 44854
rect 153022 44618 153054 44854
rect 152434 27174 153054 44618
rect 157228 45174 157548 45206
rect 157228 44938 157270 45174
rect 157506 44938 157548 45174
rect 157228 44854 157548 44938
rect 157228 44618 157270 44854
rect 157506 44618 157548 44854
rect 157228 44586 157548 44618
rect 156568 41454 156888 41486
rect 156568 41218 156610 41454
rect 156846 41218 156888 41454
rect 156568 41134 156888 41218
rect 156568 40898 156610 41134
rect 156846 40898 156888 41134
rect 156568 40866 156888 40898
rect 159874 34614 160494 52058
rect 159874 34378 159906 34614
rect 160142 34378 160226 34614
rect 160462 34378 160494 34614
rect 159874 34294 160494 34378
rect 159874 34058 159906 34294
rect 160142 34058 160226 34294
rect 160462 34058 160494 34294
rect 152434 26938 152466 27174
rect 152702 26938 152786 27174
rect 153022 26938 153054 27174
rect 152434 26854 153054 26938
rect 152434 26618 152466 26854
rect 152702 26618 152786 26854
rect 153022 26618 153054 26854
rect 151859 19412 151925 19413
rect 151859 19348 151860 19412
rect 151924 19348 151925 19412
rect 151859 19347 151925 19348
rect 148714 5218 148746 5454
rect 148982 5218 149066 5454
rect 149302 5218 149334 5454
rect 148714 5134 149334 5218
rect 148714 4898 148746 5134
rect 148982 4898 149066 5134
rect 149302 4898 149334 5134
rect 148714 -856 149334 4898
rect 151862 458 151922 19347
rect 152434 9174 153054 26618
rect 157228 27174 157548 27206
rect 157228 26938 157270 27174
rect 157506 26938 157548 27174
rect 157228 26854 157548 26938
rect 157228 26618 157270 26854
rect 157506 26618 157548 26854
rect 157228 26586 157548 26618
rect 156568 23454 156888 23486
rect 156568 23218 156610 23454
rect 156846 23218 156888 23454
rect 156568 23134 156888 23218
rect 156568 22898 156610 23134
rect 156846 22898 156888 23134
rect 156568 22866 156888 22898
rect 152434 8938 152466 9174
rect 152702 8938 152786 9174
rect 153022 8938 153054 9174
rect 152434 8854 153054 8938
rect 152434 8618 152466 8854
rect 152702 8618 152786 8854
rect 153022 8618 153054 8854
rect 148714 -1092 148746 -856
rect 148982 -1092 149066 -856
rect 149302 -1092 149334 -856
rect 148714 -1176 149334 -1092
rect 148714 -1412 148746 -1176
rect 148982 -1412 149066 -1176
rect 149302 -1412 149334 -1176
rect 148714 -4324 149334 -1412
rect 152434 -1816 153054 8618
rect 152434 -2052 152466 -1816
rect 152702 -2052 152786 -1816
rect 153022 -2052 153054 -1816
rect 152434 -2136 153054 -2052
rect 152434 -2372 152466 -2136
rect 152702 -2372 152786 -2136
rect 153022 -2372 153054 -2136
rect 152434 -4324 153054 -2372
rect 156154 12894 156774 19988
rect 156154 12658 156186 12894
rect 156422 12658 156506 12894
rect 156742 12658 156774 12894
rect 156154 12574 156774 12658
rect 156154 12338 156186 12574
rect 156422 12338 156506 12574
rect 156742 12338 156774 12574
rect 156154 -2776 156774 12338
rect 156154 -3012 156186 -2776
rect 156422 -3012 156506 -2776
rect 156742 -3012 156774 -2776
rect 156154 -3096 156774 -3012
rect 156154 -3332 156186 -3096
rect 156422 -3332 156506 -3096
rect 156742 -3332 156774 -3096
rect 156154 -4324 156774 -3332
rect 159874 16614 160494 34058
rect 159874 16378 159906 16614
rect 160142 16378 160226 16614
rect 160462 16378 160494 16614
rect 159874 16294 160494 16378
rect 159874 16058 159906 16294
rect 160142 16058 160226 16294
rect 160462 16058 160494 16294
rect 159874 -3736 160494 16058
rect 159874 -3972 159906 -3736
rect 160142 -3972 160226 -3736
rect 160462 -3972 160494 -3736
rect 159874 -4056 160494 -3972
rect 159874 -4292 159906 -4056
rect 160142 -4292 160226 -4056
rect 160462 -4292 160494 -4056
rect 159874 -4324 160494 -4292
rect 166714 461092 167334 464004
rect 166714 460856 166746 461092
rect 166982 460856 167066 461092
rect 167302 460856 167334 461092
rect 166714 460772 167334 460856
rect 166714 460536 166746 460772
rect 166982 460536 167066 460772
rect 167302 460536 167334 460772
rect 166714 455454 167334 460536
rect 166714 455218 166746 455454
rect 166982 455218 167066 455454
rect 167302 455218 167334 455454
rect 166714 455134 167334 455218
rect 166714 454898 166746 455134
rect 166982 454898 167066 455134
rect 167302 454898 167334 455134
rect 166714 437454 167334 454898
rect 166714 437218 166746 437454
rect 166982 437218 167066 437454
rect 167302 437218 167334 437454
rect 166714 437134 167334 437218
rect 166714 436898 166746 437134
rect 166982 436898 167066 437134
rect 167302 436898 167334 437134
rect 166714 419454 167334 436898
rect 166714 419218 166746 419454
rect 166982 419218 167066 419454
rect 167302 419218 167334 419454
rect 166714 419134 167334 419218
rect 166714 418898 166746 419134
rect 166982 418898 167066 419134
rect 167302 418898 167334 419134
rect 166714 401454 167334 418898
rect 166714 401218 166746 401454
rect 166982 401218 167066 401454
rect 167302 401218 167334 401454
rect 166714 401134 167334 401218
rect 166714 400898 166746 401134
rect 166982 400898 167066 401134
rect 167302 400898 167334 401134
rect 166714 383454 167334 400898
rect 166714 383218 166746 383454
rect 166982 383218 167066 383454
rect 167302 383218 167334 383454
rect 166714 383134 167334 383218
rect 166714 382898 166746 383134
rect 166982 382898 167066 383134
rect 167302 382898 167334 383134
rect 166714 365454 167334 382898
rect 166714 365218 166746 365454
rect 166982 365218 167066 365454
rect 167302 365218 167334 365454
rect 166714 365134 167334 365218
rect 166714 364898 166746 365134
rect 166982 364898 167066 365134
rect 167302 364898 167334 365134
rect 166714 347454 167334 364898
rect 166714 347218 166746 347454
rect 166982 347218 167066 347454
rect 167302 347218 167334 347454
rect 166714 347134 167334 347218
rect 166714 346898 166746 347134
rect 166982 346898 167066 347134
rect 167302 346898 167334 347134
rect 166714 329454 167334 346898
rect 166714 329218 166746 329454
rect 166982 329218 167066 329454
rect 167302 329218 167334 329454
rect 166714 329134 167334 329218
rect 166714 328898 166746 329134
rect 166982 328898 167066 329134
rect 167302 328898 167334 329134
rect 166714 311454 167334 328898
rect 166714 311218 166746 311454
rect 166982 311218 167066 311454
rect 167302 311218 167334 311454
rect 166714 311134 167334 311218
rect 166714 310898 166746 311134
rect 166982 310898 167066 311134
rect 167302 310898 167334 311134
rect 166714 293454 167334 310898
rect 166714 293218 166746 293454
rect 166982 293218 167066 293454
rect 167302 293218 167334 293454
rect 166714 293134 167334 293218
rect 166714 292898 166746 293134
rect 166982 292898 167066 293134
rect 167302 292898 167334 293134
rect 166714 275454 167334 292898
rect 166714 275218 166746 275454
rect 166982 275218 167066 275454
rect 167302 275218 167334 275454
rect 166714 275134 167334 275218
rect 166714 274898 166746 275134
rect 166982 274898 167066 275134
rect 167302 274898 167334 275134
rect 166714 257454 167334 274898
rect 166714 257218 166746 257454
rect 166982 257218 167066 257454
rect 167302 257218 167334 257454
rect 166714 257134 167334 257218
rect 166714 256898 166746 257134
rect 166982 256898 167066 257134
rect 167302 256898 167334 257134
rect 166714 239454 167334 256898
rect 166714 239218 166746 239454
rect 166982 239218 167066 239454
rect 167302 239218 167334 239454
rect 166714 239134 167334 239218
rect 166714 238898 166746 239134
rect 166982 238898 167066 239134
rect 167302 238898 167334 239134
rect 166714 221454 167334 238898
rect 166714 221218 166746 221454
rect 166982 221218 167066 221454
rect 167302 221218 167334 221454
rect 166714 221134 167334 221218
rect 166714 220898 166746 221134
rect 166982 220898 167066 221134
rect 167302 220898 167334 221134
rect 166714 203454 167334 220898
rect 166714 203218 166746 203454
rect 166982 203218 167066 203454
rect 167302 203218 167334 203454
rect 166714 203134 167334 203218
rect 166714 202898 166746 203134
rect 166982 202898 167066 203134
rect 167302 202898 167334 203134
rect 166714 185454 167334 202898
rect 166714 185218 166746 185454
rect 166982 185218 167066 185454
rect 167302 185218 167334 185454
rect 166714 185134 167334 185218
rect 166714 184898 166746 185134
rect 166982 184898 167066 185134
rect 167302 184898 167334 185134
rect 166714 167454 167334 184898
rect 166714 167218 166746 167454
rect 166982 167218 167066 167454
rect 167302 167218 167334 167454
rect 166714 167134 167334 167218
rect 166714 166898 166746 167134
rect 166982 166898 167066 167134
rect 167302 166898 167334 167134
rect 166714 149454 167334 166898
rect 166714 149218 166746 149454
rect 166982 149218 167066 149454
rect 167302 149218 167334 149454
rect 166714 149134 167334 149218
rect 166714 148898 166746 149134
rect 166982 148898 167066 149134
rect 167302 148898 167334 149134
rect 166714 131454 167334 148898
rect 166714 131218 166746 131454
rect 166982 131218 167066 131454
rect 167302 131218 167334 131454
rect 166714 131134 167334 131218
rect 166714 130898 166746 131134
rect 166982 130898 167066 131134
rect 167302 130898 167334 131134
rect 166714 113454 167334 130898
rect 166714 113218 166746 113454
rect 166982 113218 167066 113454
rect 167302 113218 167334 113454
rect 166714 113134 167334 113218
rect 166714 112898 166746 113134
rect 166982 112898 167066 113134
rect 167302 112898 167334 113134
rect 166714 95454 167334 112898
rect 166714 95218 166746 95454
rect 166982 95218 167066 95454
rect 167302 95218 167334 95454
rect 166714 95134 167334 95218
rect 166714 94898 166746 95134
rect 166982 94898 167066 95134
rect 167302 94898 167334 95134
rect 166714 77454 167334 94898
rect 166714 77218 166746 77454
rect 166982 77218 167066 77454
rect 167302 77218 167334 77454
rect 166714 77134 167334 77218
rect 166714 76898 166746 77134
rect 166982 76898 167066 77134
rect 167302 76898 167334 77134
rect 166714 59454 167334 76898
rect 166714 59218 166746 59454
rect 166982 59218 167066 59454
rect 167302 59218 167334 59454
rect 166714 59134 167334 59218
rect 166714 58898 166746 59134
rect 166982 58898 167066 59134
rect 167302 58898 167334 59134
rect 166714 41454 167334 58898
rect 166714 41218 166746 41454
rect 166982 41218 167066 41454
rect 167302 41218 167334 41454
rect 166714 41134 167334 41218
rect 166714 40898 166746 41134
rect 166982 40898 167066 41134
rect 167302 40898 167334 41134
rect 166714 23454 167334 40898
rect 166714 23218 166746 23454
rect 166982 23218 167066 23454
rect 167302 23218 167334 23454
rect 166714 23134 167334 23218
rect 166714 22898 166746 23134
rect 166982 22898 167066 23134
rect 167302 22898 167334 23134
rect 166714 5454 167334 22898
rect 166714 5218 166746 5454
rect 166982 5218 167066 5454
rect 167302 5218 167334 5454
rect 166714 5134 167334 5218
rect 166714 4898 166746 5134
rect 166982 4898 167066 5134
rect 167302 4898 167334 5134
rect 166714 -856 167334 4898
rect 166714 -1092 166746 -856
rect 166982 -1092 167066 -856
rect 167302 -1092 167334 -856
rect 166714 -1176 167334 -1092
rect 166714 -1412 166746 -1176
rect 166982 -1412 167066 -1176
rect 167302 -1412 167334 -1176
rect 166714 -4324 167334 -1412
rect 170434 462052 171054 464004
rect 170434 461816 170466 462052
rect 170702 461816 170786 462052
rect 171022 461816 171054 462052
rect 170434 461732 171054 461816
rect 170434 461496 170466 461732
rect 170702 461496 170786 461732
rect 171022 461496 171054 461732
rect 170434 441174 171054 461496
rect 170434 440938 170466 441174
rect 170702 440938 170786 441174
rect 171022 440938 171054 441174
rect 170434 440854 171054 440938
rect 170434 440618 170466 440854
rect 170702 440618 170786 440854
rect 171022 440618 171054 440854
rect 170434 423174 171054 440618
rect 170434 422938 170466 423174
rect 170702 422938 170786 423174
rect 171022 422938 171054 423174
rect 170434 422854 171054 422938
rect 170434 422618 170466 422854
rect 170702 422618 170786 422854
rect 171022 422618 171054 422854
rect 170434 405174 171054 422618
rect 170434 404938 170466 405174
rect 170702 404938 170786 405174
rect 171022 404938 171054 405174
rect 170434 404854 171054 404938
rect 170434 404618 170466 404854
rect 170702 404618 170786 404854
rect 171022 404618 171054 404854
rect 170434 387174 171054 404618
rect 170434 386938 170466 387174
rect 170702 386938 170786 387174
rect 171022 386938 171054 387174
rect 170434 386854 171054 386938
rect 170434 386618 170466 386854
rect 170702 386618 170786 386854
rect 171022 386618 171054 386854
rect 170434 369174 171054 386618
rect 170434 368938 170466 369174
rect 170702 368938 170786 369174
rect 171022 368938 171054 369174
rect 170434 368854 171054 368938
rect 170434 368618 170466 368854
rect 170702 368618 170786 368854
rect 171022 368618 171054 368854
rect 170434 351174 171054 368618
rect 170434 350938 170466 351174
rect 170702 350938 170786 351174
rect 171022 350938 171054 351174
rect 170434 350854 171054 350938
rect 170434 350618 170466 350854
rect 170702 350618 170786 350854
rect 171022 350618 171054 350854
rect 170434 333174 171054 350618
rect 170434 332938 170466 333174
rect 170702 332938 170786 333174
rect 171022 332938 171054 333174
rect 170434 332854 171054 332938
rect 170434 332618 170466 332854
rect 170702 332618 170786 332854
rect 171022 332618 171054 332854
rect 170434 315174 171054 332618
rect 170434 314938 170466 315174
rect 170702 314938 170786 315174
rect 171022 314938 171054 315174
rect 170434 314854 171054 314938
rect 170434 314618 170466 314854
rect 170702 314618 170786 314854
rect 171022 314618 171054 314854
rect 170434 297174 171054 314618
rect 170434 296938 170466 297174
rect 170702 296938 170786 297174
rect 171022 296938 171054 297174
rect 170434 296854 171054 296938
rect 170434 296618 170466 296854
rect 170702 296618 170786 296854
rect 171022 296618 171054 296854
rect 170434 279174 171054 296618
rect 170434 278938 170466 279174
rect 170702 278938 170786 279174
rect 171022 278938 171054 279174
rect 170434 278854 171054 278938
rect 170434 278618 170466 278854
rect 170702 278618 170786 278854
rect 171022 278618 171054 278854
rect 170434 261174 171054 278618
rect 170434 260938 170466 261174
rect 170702 260938 170786 261174
rect 171022 260938 171054 261174
rect 170434 260854 171054 260938
rect 170434 260618 170466 260854
rect 170702 260618 170786 260854
rect 171022 260618 171054 260854
rect 170434 243174 171054 260618
rect 170434 242938 170466 243174
rect 170702 242938 170786 243174
rect 171022 242938 171054 243174
rect 170434 242854 171054 242938
rect 170434 242618 170466 242854
rect 170702 242618 170786 242854
rect 171022 242618 171054 242854
rect 170434 225174 171054 242618
rect 170434 224938 170466 225174
rect 170702 224938 170786 225174
rect 171022 224938 171054 225174
rect 170434 224854 171054 224938
rect 170434 224618 170466 224854
rect 170702 224618 170786 224854
rect 171022 224618 171054 224854
rect 170434 207174 171054 224618
rect 170434 206938 170466 207174
rect 170702 206938 170786 207174
rect 171022 206938 171054 207174
rect 170434 206854 171054 206938
rect 170434 206618 170466 206854
rect 170702 206618 170786 206854
rect 171022 206618 171054 206854
rect 170434 189174 171054 206618
rect 170434 188938 170466 189174
rect 170702 188938 170786 189174
rect 171022 188938 171054 189174
rect 170434 188854 171054 188938
rect 170434 188618 170466 188854
rect 170702 188618 170786 188854
rect 171022 188618 171054 188854
rect 170434 171174 171054 188618
rect 170434 170938 170466 171174
rect 170702 170938 170786 171174
rect 171022 170938 171054 171174
rect 170434 170854 171054 170938
rect 170434 170618 170466 170854
rect 170702 170618 170786 170854
rect 171022 170618 171054 170854
rect 170434 153174 171054 170618
rect 170434 152938 170466 153174
rect 170702 152938 170786 153174
rect 171022 152938 171054 153174
rect 170434 152854 171054 152938
rect 170434 152618 170466 152854
rect 170702 152618 170786 152854
rect 171022 152618 171054 152854
rect 170434 135174 171054 152618
rect 170434 134938 170466 135174
rect 170702 134938 170786 135174
rect 171022 134938 171054 135174
rect 170434 134854 171054 134938
rect 170434 134618 170466 134854
rect 170702 134618 170786 134854
rect 171022 134618 171054 134854
rect 170434 117174 171054 134618
rect 170434 116938 170466 117174
rect 170702 116938 170786 117174
rect 171022 116938 171054 117174
rect 170434 116854 171054 116938
rect 170434 116618 170466 116854
rect 170702 116618 170786 116854
rect 171022 116618 171054 116854
rect 170434 99174 171054 116618
rect 170434 98938 170466 99174
rect 170702 98938 170786 99174
rect 171022 98938 171054 99174
rect 170434 98854 171054 98938
rect 170434 98618 170466 98854
rect 170702 98618 170786 98854
rect 171022 98618 171054 98854
rect 170434 81174 171054 98618
rect 170434 80938 170466 81174
rect 170702 80938 170786 81174
rect 171022 80938 171054 81174
rect 170434 80854 171054 80938
rect 170434 80618 170466 80854
rect 170702 80618 170786 80854
rect 171022 80618 171054 80854
rect 170434 63174 171054 80618
rect 170434 62938 170466 63174
rect 170702 62938 170786 63174
rect 171022 62938 171054 63174
rect 170434 62854 171054 62938
rect 170434 62618 170466 62854
rect 170702 62618 170786 62854
rect 171022 62618 171054 62854
rect 170434 45174 171054 62618
rect 170434 44938 170466 45174
rect 170702 44938 170786 45174
rect 171022 44938 171054 45174
rect 170434 44854 171054 44938
rect 170434 44618 170466 44854
rect 170702 44618 170786 44854
rect 171022 44618 171054 44854
rect 170434 27174 171054 44618
rect 170434 26938 170466 27174
rect 170702 26938 170786 27174
rect 171022 26938 171054 27174
rect 170434 26854 171054 26938
rect 170434 26618 170466 26854
rect 170702 26618 170786 26854
rect 171022 26618 171054 26854
rect 170434 9174 171054 26618
rect 170434 8938 170466 9174
rect 170702 8938 170786 9174
rect 171022 8938 171054 9174
rect 170434 8854 171054 8938
rect 170434 8618 170466 8854
rect 170702 8618 170786 8854
rect 171022 8618 171054 8854
rect 170434 -1816 171054 8618
rect 170434 -2052 170466 -1816
rect 170702 -2052 170786 -1816
rect 171022 -2052 171054 -1816
rect 170434 -2136 171054 -2052
rect 170434 -2372 170466 -2136
rect 170702 -2372 170786 -2136
rect 171022 -2372 171054 -2136
rect 170434 -4324 171054 -2372
rect 174154 463012 174774 464004
rect 174154 462776 174186 463012
rect 174422 462776 174506 463012
rect 174742 462776 174774 463012
rect 174154 462692 174774 462776
rect 174154 462456 174186 462692
rect 174422 462456 174506 462692
rect 174742 462456 174774 462692
rect 174154 444894 174774 462456
rect 174154 444658 174186 444894
rect 174422 444658 174506 444894
rect 174742 444658 174774 444894
rect 174154 444574 174774 444658
rect 174154 444338 174186 444574
rect 174422 444338 174506 444574
rect 174742 444338 174774 444574
rect 174154 426894 174774 444338
rect 174154 426658 174186 426894
rect 174422 426658 174506 426894
rect 174742 426658 174774 426894
rect 174154 426574 174774 426658
rect 174154 426338 174186 426574
rect 174422 426338 174506 426574
rect 174742 426338 174774 426574
rect 174154 408894 174774 426338
rect 174154 408658 174186 408894
rect 174422 408658 174506 408894
rect 174742 408658 174774 408894
rect 174154 408574 174774 408658
rect 174154 408338 174186 408574
rect 174422 408338 174506 408574
rect 174742 408338 174774 408574
rect 174154 390894 174774 408338
rect 174154 390658 174186 390894
rect 174422 390658 174506 390894
rect 174742 390658 174774 390894
rect 174154 390574 174774 390658
rect 174154 390338 174186 390574
rect 174422 390338 174506 390574
rect 174742 390338 174774 390574
rect 174154 372894 174774 390338
rect 174154 372658 174186 372894
rect 174422 372658 174506 372894
rect 174742 372658 174774 372894
rect 174154 372574 174774 372658
rect 174154 372338 174186 372574
rect 174422 372338 174506 372574
rect 174742 372338 174774 372574
rect 174154 354894 174774 372338
rect 174154 354658 174186 354894
rect 174422 354658 174506 354894
rect 174742 354658 174774 354894
rect 174154 354574 174774 354658
rect 174154 354338 174186 354574
rect 174422 354338 174506 354574
rect 174742 354338 174774 354574
rect 174154 336894 174774 354338
rect 174154 336658 174186 336894
rect 174422 336658 174506 336894
rect 174742 336658 174774 336894
rect 174154 336574 174774 336658
rect 174154 336338 174186 336574
rect 174422 336338 174506 336574
rect 174742 336338 174774 336574
rect 174154 318894 174774 336338
rect 174154 318658 174186 318894
rect 174422 318658 174506 318894
rect 174742 318658 174774 318894
rect 174154 318574 174774 318658
rect 174154 318338 174186 318574
rect 174422 318338 174506 318574
rect 174742 318338 174774 318574
rect 174154 300894 174774 318338
rect 174154 300658 174186 300894
rect 174422 300658 174506 300894
rect 174742 300658 174774 300894
rect 174154 300574 174774 300658
rect 174154 300338 174186 300574
rect 174422 300338 174506 300574
rect 174742 300338 174774 300574
rect 174154 282894 174774 300338
rect 174154 282658 174186 282894
rect 174422 282658 174506 282894
rect 174742 282658 174774 282894
rect 174154 282574 174774 282658
rect 174154 282338 174186 282574
rect 174422 282338 174506 282574
rect 174742 282338 174774 282574
rect 174154 264894 174774 282338
rect 174154 264658 174186 264894
rect 174422 264658 174506 264894
rect 174742 264658 174774 264894
rect 174154 264574 174774 264658
rect 174154 264338 174186 264574
rect 174422 264338 174506 264574
rect 174742 264338 174774 264574
rect 174154 246894 174774 264338
rect 174154 246658 174186 246894
rect 174422 246658 174506 246894
rect 174742 246658 174774 246894
rect 174154 246574 174774 246658
rect 174154 246338 174186 246574
rect 174422 246338 174506 246574
rect 174742 246338 174774 246574
rect 174154 228894 174774 246338
rect 174154 228658 174186 228894
rect 174422 228658 174506 228894
rect 174742 228658 174774 228894
rect 174154 228574 174774 228658
rect 174154 228338 174186 228574
rect 174422 228338 174506 228574
rect 174742 228338 174774 228574
rect 174154 210894 174774 228338
rect 174154 210658 174186 210894
rect 174422 210658 174506 210894
rect 174742 210658 174774 210894
rect 174154 210574 174774 210658
rect 174154 210338 174186 210574
rect 174422 210338 174506 210574
rect 174742 210338 174774 210574
rect 174154 192894 174774 210338
rect 174154 192658 174186 192894
rect 174422 192658 174506 192894
rect 174742 192658 174774 192894
rect 174154 192574 174774 192658
rect 174154 192338 174186 192574
rect 174422 192338 174506 192574
rect 174742 192338 174774 192574
rect 174154 174894 174774 192338
rect 174154 174658 174186 174894
rect 174422 174658 174506 174894
rect 174742 174658 174774 174894
rect 174154 174574 174774 174658
rect 174154 174338 174186 174574
rect 174422 174338 174506 174574
rect 174742 174338 174774 174574
rect 174154 156894 174774 174338
rect 174154 156658 174186 156894
rect 174422 156658 174506 156894
rect 174742 156658 174774 156894
rect 174154 156574 174774 156658
rect 174154 156338 174186 156574
rect 174422 156338 174506 156574
rect 174742 156338 174774 156574
rect 174154 138894 174774 156338
rect 174154 138658 174186 138894
rect 174422 138658 174506 138894
rect 174742 138658 174774 138894
rect 174154 138574 174774 138658
rect 174154 138338 174186 138574
rect 174422 138338 174506 138574
rect 174742 138338 174774 138574
rect 174154 120894 174774 138338
rect 174154 120658 174186 120894
rect 174422 120658 174506 120894
rect 174742 120658 174774 120894
rect 174154 120574 174774 120658
rect 174154 120338 174186 120574
rect 174422 120338 174506 120574
rect 174742 120338 174774 120574
rect 174154 102894 174774 120338
rect 174154 102658 174186 102894
rect 174422 102658 174506 102894
rect 174742 102658 174774 102894
rect 174154 102574 174774 102658
rect 174154 102338 174186 102574
rect 174422 102338 174506 102574
rect 174742 102338 174774 102574
rect 174154 84894 174774 102338
rect 174154 84658 174186 84894
rect 174422 84658 174506 84894
rect 174742 84658 174774 84894
rect 174154 84574 174774 84658
rect 174154 84338 174186 84574
rect 174422 84338 174506 84574
rect 174742 84338 174774 84574
rect 174154 66894 174774 84338
rect 174154 66658 174186 66894
rect 174422 66658 174506 66894
rect 174742 66658 174774 66894
rect 174154 66574 174774 66658
rect 174154 66338 174186 66574
rect 174422 66338 174506 66574
rect 174742 66338 174774 66574
rect 174154 48894 174774 66338
rect 174154 48658 174186 48894
rect 174422 48658 174506 48894
rect 174742 48658 174774 48894
rect 174154 48574 174774 48658
rect 174154 48338 174186 48574
rect 174422 48338 174506 48574
rect 174742 48338 174774 48574
rect 174154 30894 174774 48338
rect 174154 30658 174186 30894
rect 174422 30658 174506 30894
rect 174742 30658 174774 30894
rect 174154 30574 174774 30658
rect 174154 30338 174186 30574
rect 174422 30338 174506 30574
rect 174742 30338 174774 30574
rect 174154 12894 174774 30338
rect 174154 12658 174186 12894
rect 174422 12658 174506 12894
rect 174742 12658 174774 12894
rect 174154 12574 174774 12658
rect 174154 12338 174186 12574
rect 174422 12338 174506 12574
rect 174742 12338 174774 12574
rect 174154 -2776 174774 12338
rect 174154 -3012 174186 -2776
rect 174422 -3012 174506 -2776
rect 174742 -3012 174774 -2776
rect 174154 -3096 174774 -3012
rect 174154 -3332 174186 -3096
rect 174422 -3332 174506 -3096
rect 174742 -3332 174774 -3096
rect 174154 -4324 174774 -3332
rect 177874 463972 178494 464004
rect 177874 463736 177906 463972
rect 178142 463736 178226 463972
rect 178462 463736 178494 463972
rect 177874 463652 178494 463736
rect 177874 463416 177906 463652
rect 178142 463416 178226 463652
rect 178462 463416 178494 463652
rect 177874 448614 178494 463416
rect 177874 448378 177906 448614
rect 178142 448378 178226 448614
rect 178462 448378 178494 448614
rect 177874 448294 178494 448378
rect 177874 448058 177906 448294
rect 178142 448058 178226 448294
rect 178462 448058 178494 448294
rect 177874 430614 178494 448058
rect 177874 430378 177906 430614
rect 178142 430378 178226 430614
rect 178462 430378 178494 430614
rect 177874 430294 178494 430378
rect 177874 430058 177906 430294
rect 178142 430058 178226 430294
rect 178462 430058 178494 430294
rect 177874 412614 178494 430058
rect 177874 412378 177906 412614
rect 178142 412378 178226 412614
rect 178462 412378 178494 412614
rect 177874 412294 178494 412378
rect 177874 412058 177906 412294
rect 178142 412058 178226 412294
rect 178462 412058 178494 412294
rect 177874 394614 178494 412058
rect 177874 394378 177906 394614
rect 178142 394378 178226 394614
rect 178462 394378 178494 394614
rect 177874 394294 178494 394378
rect 177874 394058 177906 394294
rect 178142 394058 178226 394294
rect 178462 394058 178494 394294
rect 177874 376614 178494 394058
rect 177874 376378 177906 376614
rect 178142 376378 178226 376614
rect 178462 376378 178494 376614
rect 177874 376294 178494 376378
rect 177874 376058 177906 376294
rect 178142 376058 178226 376294
rect 178462 376058 178494 376294
rect 177874 358614 178494 376058
rect 177874 358378 177906 358614
rect 178142 358378 178226 358614
rect 178462 358378 178494 358614
rect 177874 358294 178494 358378
rect 177874 358058 177906 358294
rect 178142 358058 178226 358294
rect 178462 358058 178494 358294
rect 177874 340614 178494 358058
rect 177874 340378 177906 340614
rect 178142 340378 178226 340614
rect 178462 340378 178494 340614
rect 177874 340294 178494 340378
rect 177874 340058 177906 340294
rect 178142 340058 178226 340294
rect 178462 340058 178494 340294
rect 177874 322614 178494 340058
rect 177874 322378 177906 322614
rect 178142 322378 178226 322614
rect 178462 322378 178494 322614
rect 177874 322294 178494 322378
rect 177874 322058 177906 322294
rect 178142 322058 178226 322294
rect 178462 322058 178494 322294
rect 177874 304614 178494 322058
rect 177874 304378 177906 304614
rect 178142 304378 178226 304614
rect 178462 304378 178494 304614
rect 177874 304294 178494 304378
rect 177874 304058 177906 304294
rect 178142 304058 178226 304294
rect 178462 304058 178494 304294
rect 177874 286614 178494 304058
rect 177874 286378 177906 286614
rect 178142 286378 178226 286614
rect 178462 286378 178494 286614
rect 177874 286294 178494 286378
rect 177874 286058 177906 286294
rect 178142 286058 178226 286294
rect 178462 286058 178494 286294
rect 177874 268614 178494 286058
rect 177874 268378 177906 268614
rect 178142 268378 178226 268614
rect 178462 268378 178494 268614
rect 177874 268294 178494 268378
rect 177874 268058 177906 268294
rect 178142 268058 178226 268294
rect 178462 268058 178494 268294
rect 177874 250614 178494 268058
rect 177874 250378 177906 250614
rect 178142 250378 178226 250614
rect 178462 250378 178494 250614
rect 177874 250294 178494 250378
rect 177874 250058 177906 250294
rect 178142 250058 178226 250294
rect 178462 250058 178494 250294
rect 177874 232614 178494 250058
rect 177874 232378 177906 232614
rect 178142 232378 178226 232614
rect 178462 232378 178494 232614
rect 177874 232294 178494 232378
rect 177874 232058 177906 232294
rect 178142 232058 178226 232294
rect 178462 232058 178494 232294
rect 177874 214614 178494 232058
rect 177874 214378 177906 214614
rect 178142 214378 178226 214614
rect 178462 214378 178494 214614
rect 177874 214294 178494 214378
rect 177874 214058 177906 214294
rect 178142 214058 178226 214294
rect 178462 214058 178494 214294
rect 177874 196614 178494 214058
rect 177874 196378 177906 196614
rect 178142 196378 178226 196614
rect 178462 196378 178494 196614
rect 177874 196294 178494 196378
rect 177874 196058 177906 196294
rect 178142 196058 178226 196294
rect 178462 196058 178494 196294
rect 177874 178614 178494 196058
rect 177874 178378 177906 178614
rect 178142 178378 178226 178614
rect 178462 178378 178494 178614
rect 177874 178294 178494 178378
rect 177874 178058 177906 178294
rect 178142 178058 178226 178294
rect 178462 178058 178494 178294
rect 177874 160614 178494 178058
rect 177874 160378 177906 160614
rect 178142 160378 178226 160614
rect 178462 160378 178494 160614
rect 177874 160294 178494 160378
rect 177874 160058 177906 160294
rect 178142 160058 178226 160294
rect 178462 160058 178494 160294
rect 177874 142614 178494 160058
rect 177874 142378 177906 142614
rect 178142 142378 178226 142614
rect 178462 142378 178494 142614
rect 177874 142294 178494 142378
rect 177874 142058 177906 142294
rect 178142 142058 178226 142294
rect 178462 142058 178494 142294
rect 177874 124614 178494 142058
rect 177874 124378 177906 124614
rect 178142 124378 178226 124614
rect 178462 124378 178494 124614
rect 177874 124294 178494 124378
rect 177874 124058 177906 124294
rect 178142 124058 178226 124294
rect 178462 124058 178494 124294
rect 177874 106614 178494 124058
rect 177874 106378 177906 106614
rect 178142 106378 178226 106614
rect 178462 106378 178494 106614
rect 177874 106294 178494 106378
rect 177874 106058 177906 106294
rect 178142 106058 178226 106294
rect 178462 106058 178494 106294
rect 177874 88614 178494 106058
rect 177874 88378 177906 88614
rect 178142 88378 178226 88614
rect 178462 88378 178494 88614
rect 177874 88294 178494 88378
rect 177874 88058 177906 88294
rect 178142 88058 178226 88294
rect 178462 88058 178494 88294
rect 177874 70614 178494 88058
rect 177874 70378 177906 70614
rect 178142 70378 178226 70614
rect 178462 70378 178494 70614
rect 177874 70294 178494 70378
rect 177874 70058 177906 70294
rect 178142 70058 178226 70294
rect 178462 70058 178494 70294
rect 177874 52614 178494 70058
rect 177874 52378 177906 52614
rect 178142 52378 178226 52614
rect 178462 52378 178494 52614
rect 177874 52294 178494 52378
rect 177874 52058 177906 52294
rect 178142 52058 178226 52294
rect 178462 52058 178494 52294
rect 177874 34614 178494 52058
rect 177874 34378 177906 34614
rect 178142 34378 178226 34614
rect 178462 34378 178494 34614
rect 177874 34294 178494 34378
rect 177874 34058 177906 34294
rect 178142 34058 178226 34294
rect 178462 34058 178494 34294
rect 177874 16614 178494 34058
rect 177874 16378 177906 16614
rect 178142 16378 178226 16614
rect 178462 16378 178494 16614
rect 177874 16294 178494 16378
rect 177874 16058 177906 16294
rect 178142 16058 178226 16294
rect 178462 16058 178494 16294
rect 177874 -3736 178494 16058
rect 177874 -3972 177906 -3736
rect 178142 -3972 178226 -3736
rect 178462 -3972 178494 -3736
rect 177874 -4056 178494 -3972
rect 177874 -4292 177906 -4056
rect 178142 -4292 178226 -4056
rect 178462 -4292 178494 -4056
rect 177874 -4324 178494 -4292
rect 184714 461092 185334 464004
rect 184714 460856 184746 461092
rect 184982 460856 185066 461092
rect 185302 460856 185334 461092
rect 184714 460772 185334 460856
rect 184714 460536 184746 460772
rect 184982 460536 185066 460772
rect 185302 460536 185334 460772
rect 184714 455454 185334 460536
rect 184714 455218 184746 455454
rect 184982 455218 185066 455454
rect 185302 455218 185334 455454
rect 184714 455134 185334 455218
rect 184714 454898 184746 455134
rect 184982 454898 185066 455134
rect 185302 454898 185334 455134
rect 184714 437454 185334 454898
rect 184714 437218 184746 437454
rect 184982 437218 185066 437454
rect 185302 437218 185334 437454
rect 184714 437134 185334 437218
rect 184714 436898 184746 437134
rect 184982 436898 185066 437134
rect 185302 436898 185334 437134
rect 184714 419454 185334 436898
rect 184714 419218 184746 419454
rect 184982 419218 185066 419454
rect 185302 419218 185334 419454
rect 184714 419134 185334 419218
rect 184714 418898 184746 419134
rect 184982 418898 185066 419134
rect 185302 418898 185334 419134
rect 184714 401454 185334 418898
rect 184714 401218 184746 401454
rect 184982 401218 185066 401454
rect 185302 401218 185334 401454
rect 184714 401134 185334 401218
rect 184714 400898 184746 401134
rect 184982 400898 185066 401134
rect 185302 400898 185334 401134
rect 184714 383454 185334 400898
rect 184714 383218 184746 383454
rect 184982 383218 185066 383454
rect 185302 383218 185334 383454
rect 184714 383134 185334 383218
rect 184714 382898 184746 383134
rect 184982 382898 185066 383134
rect 185302 382898 185334 383134
rect 184714 365454 185334 382898
rect 184714 365218 184746 365454
rect 184982 365218 185066 365454
rect 185302 365218 185334 365454
rect 184714 365134 185334 365218
rect 184714 364898 184746 365134
rect 184982 364898 185066 365134
rect 185302 364898 185334 365134
rect 184714 347454 185334 364898
rect 184714 347218 184746 347454
rect 184982 347218 185066 347454
rect 185302 347218 185334 347454
rect 184714 347134 185334 347218
rect 184714 346898 184746 347134
rect 184982 346898 185066 347134
rect 185302 346898 185334 347134
rect 184714 329454 185334 346898
rect 184714 329218 184746 329454
rect 184982 329218 185066 329454
rect 185302 329218 185334 329454
rect 184714 329134 185334 329218
rect 184714 328898 184746 329134
rect 184982 328898 185066 329134
rect 185302 328898 185334 329134
rect 184714 311454 185334 328898
rect 184714 311218 184746 311454
rect 184982 311218 185066 311454
rect 185302 311218 185334 311454
rect 184714 311134 185334 311218
rect 184714 310898 184746 311134
rect 184982 310898 185066 311134
rect 185302 310898 185334 311134
rect 184714 293454 185334 310898
rect 184714 293218 184746 293454
rect 184982 293218 185066 293454
rect 185302 293218 185334 293454
rect 184714 293134 185334 293218
rect 184714 292898 184746 293134
rect 184982 292898 185066 293134
rect 185302 292898 185334 293134
rect 184714 275454 185334 292898
rect 184714 275218 184746 275454
rect 184982 275218 185066 275454
rect 185302 275218 185334 275454
rect 184714 275134 185334 275218
rect 184714 274898 184746 275134
rect 184982 274898 185066 275134
rect 185302 274898 185334 275134
rect 184714 257454 185334 274898
rect 184714 257218 184746 257454
rect 184982 257218 185066 257454
rect 185302 257218 185334 257454
rect 184714 257134 185334 257218
rect 184714 256898 184746 257134
rect 184982 256898 185066 257134
rect 185302 256898 185334 257134
rect 184714 239454 185334 256898
rect 184714 239218 184746 239454
rect 184982 239218 185066 239454
rect 185302 239218 185334 239454
rect 184714 239134 185334 239218
rect 184714 238898 184746 239134
rect 184982 238898 185066 239134
rect 185302 238898 185334 239134
rect 184714 221454 185334 238898
rect 184714 221218 184746 221454
rect 184982 221218 185066 221454
rect 185302 221218 185334 221454
rect 184714 221134 185334 221218
rect 184714 220898 184746 221134
rect 184982 220898 185066 221134
rect 185302 220898 185334 221134
rect 184714 203454 185334 220898
rect 184714 203218 184746 203454
rect 184982 203218 185066 203454
rect 185302 203218 185334 203454
rect 184714 203134 185334 203218
rect 184714 202898 184746 203134
rect 184982 202898 185066 203134
rect 185302 202898 185334 203134
rect 184714 185454 185334 202898
rect 184714 185218 184746 185454
rect 184982 185218 185066 185454
rect 185302 185218 185334 185454
rect 184714 185134 185334 185218
rect 184714 184898 184746 185134
rect 184982 184898 185066 185134
rect 185302 184898 185334 185134
rect 184714 167454 185334 184898
rect 184714 167218 184746 167454
rect 184982 167218 185066 167454
rect 185302 167218 185334 167454
rect 184714 167134 185334 167218
rect 184714 166898 184746 167134
rect 184982 166898 185066 167134
rect 185302 166898 185334 167134
rect 184714 149454 185334 166898
rect 184714 149218 184746 149454
rect 184982 149218 185066 149454
rect 185302 149218 185334 149454
rect 184714 149134 185334 149218
rect 184714 148898 184746 149134
rect 184982 148898 185066 149134
rect 185302 148898 185334 149134
rect 184714 131454 185334 148898
rect 184714 131218 184746 131454
rect 184982 131218 185066 131454
rect 185302 131218 185334 131454
rect 184714 131134 185334 131218
rect 184714 130898 184746 131134
rect 184982 130898 185066 131134
rect 185302 130898 185334 131134
rect 184714 113454 185334 130898
rect 184714 113218 184746 113454
rect 184982 113218 185066 113454
rect 185302 113218 185334 113454
rect 184714 113134 185334 113218
rect 184714 112898 184746 113134
rect 184982 112898 185066 113134
rect 185302 112898 185334 113134
rect 184714 95454 185334 112898
rect 184714 95218 184746 95454
rect 184982 95218 185066 95454
rect 185302 95218 185334 95454
rect 184714 95134 185334 95218
rect 184714 94898 184746 95134
rect 184982 94898 185066 95134
rect 185302 94898 185334 95134
rect 184714 77454 185334 94898
rect 184714 77218 184746 77454
rect 184982 77218 185066 77454
rect 185302 77218 185334 77454
rect 184714 77134 185334 77218
rect 184714 76898 184746 77134
rect 184982 76898 185066 77134
rect 185302 76898 185334 77134
rect 184714 59454 185334 76898
rect 184714 59218 184746 59454
rect 184982 59218 185066 59454
rect 185302 59218 185334 59454
rect 184714 59134 185334 59218
rect 184714 58898 184746 59134
rect 184982 58898 185066 59134
rect 185302 58898 185334 59134
rect 184714 41454 185334 58898
rect 184714 41218 184746 41454
rect 184982 41218 185066 41454
rect 185302 41218 185334 41454
rect 184714 41134 185334 41218
rect 184714 40898 184746 41134
rect 184982 40898 185066 41134
rect 185302 40898 185334 41134
rect 184714 23454 185334 40898
rect 184714 23218 184746 23454
rect 184982 23218 185066 23454
rect 185302 23218 185334 23454
rect 184714 23134 185334 23218
rect 184714 22898 184746 23134
rect 184982 22898 185066 23134
rect 185302 22898 185334 23134
rect 184714 5454 185334 22898
rect 184714 5218 184746 5454
rect 184982 5218 185066 5454
rect 185302 5218 185334 5454
rect 184714 5134 185334 5218
rect 184714 4898 184746 5134
rect 184982 4898 185066 5134
rect 185302 4898 185334 5134
rect 184714 -856 185334 4898
rect 184714 -1092 184746 -856
rect 184982 -1092 185066 -856
rect 185302 -1092 185334 -856
rect 184714 -1176 185334 -1092
rect 184714 -1412 184746 -1176
rect 184982 -1412 185066 -1176
rect 185302 -1412 185334 -1176
rect 184714 -4324 185334 -1412
rect 188434 462052 189054 464004
rect 188434 461816 188466 462052
rect 188702 461816 188786 462052
rect 189022 461816 189054 462052
rect 188434 461732 189054 461816
rect 188434 461496 188466 461732
rect 188702 461496 188786 461732
rect 189022 461496 189054 461732
rect 188434 441174 189054 461496
rect 188434 440938 188466 441174
rect 188702 440938 188786 441174
rect 189022 440938 189054 441174
rect 188434 440854 189054 440938
rect 188434 440618 188466 440854
rect 188702 440618 188786 440854
rect 189022 440618 189054 440854
rect 188434 423174 189054 440618
rect 188434 422938 188466 423174
rect 188702 422938 188786 423174
rect 189022 422938 189054 423174
rect 188434 422854 189054 422938
rect 188434 422618 188466 422854
rect 188702 422618 188786 422854
rect 189022 422618 189054 422854
rect 188434 405174 189054 422618
rect 188434 404938 188466 405174
rect 188702 404938 188786 405174
rect 189022 404938 189054 405174
rect 188434 404854 189054 404938
rect 188434 404618 188466 404854
rect 188702 404618 188786 404854
rect 189022 404618 189054 404854
rect 188434 387174 189054 404618
rect 188434 386938 188466 387174
rect 188702 386938 188786 387174
rect 189022 386938 189054 387174
rect 188434 386854 189054 386938
rect 188434 386618 188466 386854
rect 188702 386618 188786 386854
rect 189022 386618 189054 386854
rect 188434 369174 189054 386618
rect 188434 368938 188466 369174
rect 188702 368938 188786 369174
rect 189022 368938 189054 369174
rect 188434 368854 189054 368938
rect 188434 368618 188466 368854
rect 188702 368618 188786 368854
rect 189022 368618 189054 368854
rect 188434 351174 189054 368618
rect 188434 350938 188466 351174
rect 188702 350938 188786 351174
rect 189022 350938 189054 351174
rect 188434 350854 189054 350938
rect 188434 350618 188466 350854
rect 188702 350618 188786 350854
rect 189022 350618 189054 350854
rect 188434 333174 189054 350618
rect 188434 332938 188466 333174
rect 188702 332938 188786 333174
rect 189022 332938 189054 333174
rect 188434 332854 189054 332938
rect 188434 332618 188466 332854
rect 188702 332618 188786 332854
rect 189022 332618 189054 332854
rect 188434 315174 189054 332618
rect 188434 314938 188466 315174
rect 188702 314938 188786 315174
rect 189022 314938 189054 315174
rect 188434 314854 189054 314938
rect 188434 314618 188466 314854
rect 188702 314618 188786 314854
rect 189022 314618 189054 314854
rect 188434 297174 189054 314618
rect 188434 296938 188466 297174
rect 188702 296938 188786 297174
rect 189022 296938 189054 297174
rect 188434 296854 189054 296938
rect 188434 296618 188466 296854
rect 188702 296618 188786 296854
rect 189022 296618 189054 296854
rect 188434 279174 189054 296618
rect 188434 278938 188466 279174
rect 188702 278938 188786 279174
rect 189022 278938 189054 279174
rect 188434 278854 189054 278938
rect 188434 278618 188466 278854
rect 188702 278618 188786 278854
rect 189022 278618 189054 278854
rect 188434 261174 189054 278618
rect 188434 260938 188466 261174
rect 188702 260938 188786 261174
rect 189022 260938 189054 261174
rect 188434 260854 189054 260938
rect 188434 260618 188466 260854
rect 188702 260618 188786 260854
rect 189022 260618 189054 260854
rect 188434 243174 189054 260618
rect 188434 242938 188466 243174
rect 188702 242938 188786 243174
rect 189022 242938 189054 243174
rect 188434 242854 189054 242938
rect 188434 242618 188466 242854
rect 188702 242618 188786 242854
rect 189022 242618 189054 242854
rect 188434 225174 189054 242618
rect 188434 224938 188466 225174
rect 188702 224938 188786 225174
rect 189022 224938 189054 225174
rect 188434 224854 189054 224938
rect 188434 224618 188466 224854
rect 188702 224618 188786 224854
rect 189022 224618 189054 224854
rect 188434 207174 189054 224618
rect 188434 206938 188466 207174
rect 188702 206938 188786 207174
rect 189022 206938 189054 207174
rect 188434 206854 189054 206938
rect 188434 206618 188466 206854
rect 188702 206618 188786 206854
rect 189022 206618 189054 206854
rect 188434 189174 189054 206618
rect 188434 188938 188466 189174
rect 188702 188938 188786 189174
rect 189022 188938 189054 189174
rect 188434 188854 189054 188938
rect 188434 188618 188466 188854
rect 188702 188618 188786 188854
rect 189022 188618 189054 188854
rect 188434 171174 189054 188618
rect 188434 170938 188466 171174
rect 188702 170938 188786 171174
rect 189022 170938 189054 171174
rect 188434 170854 189054 170938
rect 188434 170618 188466 170854
rect 188702 170618 188786 170854
rect 189022 170618 189054 170854
rect 188434 153174 189054 170618
rect 188434 152938 188466 153174
rect 188702 152938 188786 153174
rect 189022 152938 189054 153174
rect 188434 152854 189054 152938
rect 188434 152618 188466 152854
rect 188702 152618 188786 152854
rect 189022 152618 189054 152854
rect 188434 135174 189054 152618
rect 188434 134938 188466 135174
rect 188702 134938 188786 135174
rect 189022 134938 189054 135174
rect 188434 134854 189054 134938
rect 188434 134618 188466 134854
rect 188702 134618 188786 134854
rect 189022 134618 189054 134854
rect 188434 117174 189054 134618
rect 188434 116938 188466 117174
rect 188702 116938 188786 117174
rect 189022 116938 189054 117174
rect 188434 116854 189054 116938
rect 188434 116618 188466 116854
rect 188702 116618 188786 116854
rect 189022 116618 189054 116854
rect 188434 99174 189054 116618
rect 188434 98938 188466 99174
rect 188702 98938 188786 99174
rect 189022 98938 189054 99174
rect 188434 98854 189054 98938
rect 188434 98618 188466 98854
rect 188702 98618 188786 98854
rect 189022 98618 189054 98854
rect 188434 81174 189054 98618
rect 188434 80938 188466 81174
rect 188702 80938 188786 81174
rect 189022 80938 189054 81174
rect 188434 80854 189054 80938
rect 188434 80618 188466 80854
rect 188702 80618 188786 80854
rect 189022 80618 189054 80854
rect 188434 63174 189054 80618
rect 188434 62938 188466 63174
rect 188702 62938 188786 63174
rect 189022 62938 189054 63174
rect 188434 62854 189054 62938
rect 188434 62618 188466 62854
rect 188702 62618 188786 62854
rect 189022 62618 189054 62854
rect 188434 45174 189054 62618
rect 188434 44938 188466 45174
rect 188702 44938 188786 45174
rect 189022 44938 189054 45174
rect 188434 44854 189054 44938
rect 188434 44618 188466 44854
rect 188702 44618 188786 44854
rect 189022 44618 189054 44854
rect 188434 27174 189054 44618
rect 188434 26938 188466 27174
rect 188702 26938 188786 27174
rect 189022 26938 189054 27174
rect 188434 26854 189054 26938
rect 188434 26618 188466 26854
rect 188702 26618 188786 26854
rect 189022 26618 189054 26854
rect 188434 9174 189054 26618
rect 188434 8938 188466 9174
rect 188702 8938 188786 9174
rect 189022 8938 189054 9174
rect 188434 8854 189054 8938
rect 188434 8618 188466 8854
rect 188702 8618 188786 8854
rect 189022 8618 189054 8854
rect 188434 -1816 189054 8618
rect 188434 -2052 188466 -1816
rect 188702 -2052 188786 -1816
rect 189022 -2052 189054 -1816
rect 188434 -2136 189054 -2052
rect 188434 -2372 188466 -2136
rect 188702 -2372 188786 -2136
rect 189022 -2372 189054 -2136
rect 188434 -4324 189054 -2372
rect 192154 463012 192774 464004
rect 192154 462776 192186 463012
rect 192422 462776 192506 463012
rect 192742 462776 192774 463012
rect 192154 462692 192774 462776
rect 192154 462456 192186 462692
rect 192422 462456 192506 462692
rect 192742 462456 192774 462692
rect 192154 444894 192774 462456
rect 192154 444658 192186 444894
rect 192422 444658 192506 444894
rect 192742 444658 192774 444894
rect 192154 444574 192774 444658
rect 192154 444338 192186 444574
rect 192422 444338 192506 444574
rect 192742 444338 192774 444574
rect 192154 426894 192774 444338
rect 192154 426658 192186 426894
rect 192422 426658 192506 426894
rect 192742 426658 192774 426894
rect 192154 426574 192774 426658
rect 192154 426338 192186 426574
rect 192422 426338 192506 426574
rect 192742 426338 192774 426574
rect 192154 408894 192774 426338
rect 192154 408658 192186 408894
rect 192422 408658 192506 408894
rect 192742 408658 192774 408894
rect 192154 408574 192774 408658
rect 192154 408338 192186 408574
rect 192422 408338 192506 408574
rect 192742 408338 192774 408574
rect 192154 390894 192774 408338
rect 192154 390658 192186 390894
rect 192422 390658 192506 390894
rect 192742 390658 192774 390894
rect 192154 390574 192774 390658
rect 192154 390338 192186 390574
rect 192422 390338 192506 390574
rect 192742 390338 192774 390574
rect 192154 372894 192774 390338
rect 192154 372658 192186 372894
rect 192422 372658 192506 372894
rect 192742 372658 192774 372894
rect 192154 372574 192774 372658
rect 192154 372338 192186 372574
rect 192422 372338 192506 372574
rect 192742 372338 192774 372574
rect 192154 354894 192774 372338
rect 192154 354658 192186 354894
rect 192422 354658 192506 354894
rect 192742 354658 192774 354894
rect 192154 354574 192774 354658
rect 192154 354338 192186 354574
rect 192422 354338 192506 354574
rect 192742 354338 192774 354574
rect 192154 336894 192774 354338
rect 192154 336658 192186 336894
rect 192422 336658 192506 336894
rect 192742 336658 192774 336894
rect 192154 336574 192774 336658
rect 192154 336338 192186 336574
rect 192422 336338 192506 336574
rect 192742 336338 192774 336574
rect 192154 318894 192774 336338
rect 192154 318658 192186 318894
rect 192422 318658 192506 318894
rect 192742 318658 192774 318894
rect 192154 318574 192774 318658
rect 192154 318338 192186 318574
rect 192422 318338 192506 318574
rect 192742 318338 192774 318574
rect 192154 300894 192774 318338
rect 192154 300658 192186 300894
rect 192422 300658 192506 300894
rect 192742 300658 192774 300894
rect 192154 300574 192774 300658
rect 192154 300338 192186 300574
rect 192422 300338 192506 300574
rect 192742 300338 192774 300574
rect 192154 282894 192774 300338
rect 192154 282658 192186 282894
rect 192422 282658 192506 282894
rect 192742 282658 192774 282894
rect 192154 282574 192774 282658
rect 192154 282338 192186 282574
rect 192422 282338 192506 282574
rect 192742 282338 192774 282574
rect 192154 264894 192774 282338
rect 192154 264658 192186 264894
rect 192422 264658 192506 264894
rect 192742 264658 192774 264894
rect 192154 264574 192774 264658
rect 192154 264338 192186 264574
rect 192422 264338 192506 264574
rect 192742 264338 192774 264574
rect 192154 246894 192774 264338
rect 192154 246658 192186 246894
rect 192422 246658 192506 246894
rect 192742 246658 192774 246894
rect 192154 246574 192774 246658
rect 192154 246338 192186 246574
rect 192422 246338 192506 246574
rect 192742 246338 192774 246574
rect 192154 228894 192774 246338
rect 192154 228658 192186 228894
rect 192422 228658 192506 228894
rect 192742 228658 192774 228894
rect 192154 228574 192774 228658
rect 192154 228338 192186 228574
rect 192422 228338 192506 228574
rect 192742 228338 192774 228574
rect 192154 210894 192774 228338
rect 192154 210658 192186 210894
rect 192422 210658 192506 210894
rect 192742 210658 192774 210894
rect 192154 210574 192774 210658
rect 192154 210338 192186 210574
rect 192422 210338 192506 210574
rect 192742 210338 192774 210574
rect 192154 192894 192774 210338
rect 192154 192658 192186 192894
rect 192422 192658 192506 192894
rect 192742 192658 192774 192894
rect 192154 192574 192774 192658
rect 192154 192338 192186 192574
rect 192422 192338 192506 192574
rect 192742 192338 192774 192574
rect 192154 174894 192774 192338
rect 192154 174658 192186 174894
rect 192422 174658 192506 174894
rect 192742 174658 192774 174894
rect 192154 174574 192774 174658
rect 192154 174338 192186 174574
rect 192422 174338 192506 174574
rect 192742 174338 192774 174574
rect 192154 156894 192774 174338
rect 192154 156658 192186 156894
rect 192422 156658 192506 156894
rect 192742 156658 192774 156894
rect 192154 156574 192774 156658
rect 192154 156338 192186 156574
rect 192422 156338 192506 156574
rect 192742 156338 192774 156574
rect 192154 138894 192774 156338
rect 192154 138658 192186 138894
rect 192422 138658 192506 138894
rect 192742 138658 192774 138894
rect 192154 138574 192774 138658
rect 192154 138338 192186 138574
rect 192422 138338 192506 138574
rect 192742 138338 192774 138574
rect 192154 120894 192774 138338
rect 192154 120658 192186 120894
rect 192422 120658 192506 120894
rect 192742 120658 192774 120894
rect 192154 120574 192774 120658
rect 192154 120338 192186 120574
rect 192422 120338 192506 120574
rect 192742 120338 192774 120574
rect 192154 102894 192774 120338
rect 192154 102658 192186 102894
rect 192422 102658 192506 102894
rect 192742 102658 192774 102894
rect 192154 102574 192774 102658
rect 192154 102338 192186 102574
rect 192422 102338 192506 102574
rect 192742 102338 192774 102574
rect 192154 84894 192774 102338
rect 192154 84658 192186 84894
rect 192422 84658 192506 84894
rect 192742 84658 192774 84894
rect 192154 84574 192774 84658
rect 192154 84338 192186 84574
rect 192422 84338 192506 84574
rect 192742 84338 192774 84574
rect 192154 66894 192774 84338
rect 192154 66658 192186 66894
rect 192422 66658 192506 66894
rect 192742 66658 192774 66894
rect 192154 66574 192774 66658
rect 192154 66338 192186 66574
rect 192422 66338 192506 66574
rect 192742 66338 192774 66574
rect 192154 48894 192774 66338
rect 192154 48658 192186 48894
rect 192422 48658 192506 48894
rect 192742 48658 192774 48894
rect 192154 48574 192774 48658
rect 192154 48338 192186 48574
rect 192422 48338 192506 48574
rect 192742 48338 192774 48574
rect 192154 30894 192774 48338
rect 192154 30658 192186 30894
rect 192422 30658 192506 30894
rect 192742 30658 192774 30894
rect 192154 30574 192774 30658
rect 192154 30338 192186 30574
rect 192422 30338 192506 30574
rect 192742 30338 192774 30574
rect 192154 12894 192774 30338
rect 192154 12658 192186 12894
rect 192422 12658 192506 12894
rect 192742 12658 192774 12894
rect 192154 12574 192774 12658
rect 192154 12338 192186 12574
rect 192422 12338 192506 12574
rect 192742 12338 192774 12574
rect 192154 -2776 192774 12338
rect 192154 -3012 192186 -2776
rect 192422 -3012 192506 -2776
rect 192742 -3012 192774 -2776
rect 192154 -3096 192774 -3012
rect 192154 -3332 192186 -3096
rect 192422 -3332 192506 -3096
rect 192742 -3332 192774 -3096
rect 192154 -4324 192774 -3332
rect 195874 463972 196494 464004
rect 195874 463736 195906 463972
rect 196142 463736 196226 463972
rect 196462 463736 196494 463972
rect 195874 463652 196494 463736
rect 195874 463416 195906 463652
rect 196142 463416 196226 463652
rect 196462 463416 196494 463652
rect 195874 448614 196494 463416
rect 195874 448378 195906 448614
rect 196142 448378 196226 448614
rect 196462 448378 196494 448614
rect 195874 448294 196494 448378
rect 195874 448058 195906 448294
rect 196142 448058 196226 448294
rect 196462 448058 196494 448294
rect 195874 430614 196494 448058
rect 195874 430378 195906 430614
rect 196142 430378 196226 430614
rect 196462 430378 196494 430614
rect 195874 430294 196494 430378
rect 195874 430058 195906 430294
rect 196142 430058 196226 430294
rect 196462 430058 196494 430294
rect 195874 412614 196494 430058
rect 195874 412378 195906 412614
rect 196142 412378 196226 412614
rect 196462 412378 196494 412614
rect 195874 412294 196494 412378
rect 195874 412058 195906 412294
rect 196142 412058 196226 412294
rect 196462 412058 196494 412294
rect 195874 394614 196494 412058
rect 195874 394378 195906 394614
rect 196142 394378 196226 394614
rect 196462 394378 196494 394614
rect 195874 394294 196494 394378
rect 195874 394058 195906 394294
rect 196142 394058 196226 394294
rect 196462 394058 196494 394294
rect 195874 376614 196494 394058
rect 195874 376378 195906 376614
rect 196142 376378 196226 376614
rect 196462 376378 196494 376614
rect 195874 376294 196494 376378
rect 195874 376058 195906 376294
rect 196142 376058 196226 376294
rect 196462 376058 196494 376294
rect 195874 358614 196494 376058
rect 195874 358378 195906 358614
rect 196142 358378 196226 358614
rect 196462 358378 196494 358614
rect 195874 358294 196494 358378
rect 195874 358058 195906 358294
rect 196142 358058 196226 358294
rect 196462 358058 196494 358294
rect 195874 340614 196494 358058
rect 195874 340378 195906 340614
rect 196142 340378 196226 340614
rect 196462 340378 196494 340614
rect 195874 340294 196494 340378
rect 195874 340058 195906 340294
rect 196142 340058 196226 340294
rect 196462 340058 196494 340294
rect 195874 322614 196494 340058
rect 195874 322378 195906 322614
rect 196142 322378 196226 322614
rect 196462 322378 196494 322614
rect 195874 322294 196494 322378
rect 195874 322058 195906 322294
rect 196142 322058 196226 322294
rect 196462 322058 196494 322294
rect 195874 304614 196494 322058
rect 195874 304378 195906 304614
rect 196142 304378 196226 304614
rect 196462 304378 196494 304614
rect 195874 304294 196494 304378
rect 195874 304058 195906 304294
rect 196142 304058 196226 304294
rect 196462 304058 196494 304294
rect 195874 286614 196494 304058
rect 195874 286378 195906 286614
rect 196142 286378 196226 286614
rect 196462 286378 196494 286614
rect 195874 286294 196494 286378
rect 195874 286058 195906 286294
rect 196142 286058 196226 286294
rect 196462 286058 196494 286294
rect 195874 268614 196494 286058
rect 195874 268378 195906 268614
rect 196142 268378 196226 268614
rect 196462 268378 196494 268614
rect 195874 268294 196494 268378
rect 195874 268058 195906 268294
rect 196142 268058 196226 268294
rect 196462 268058 196494 268294
rect 195874 250614 196494 268058
rect 195874 250378 195906 250614
rect 196142 250378 196226 250614
rect 196462 250378 196494 250614
rect 195874 250294 196494 250378
rect 195874 250058 195906 250294
rect 196142 250058 196226 250294
rect 196462 250058 196494 250294
rect 195874 232614 196494 250058
rect 195874 232378 195906 232614
rect 196142 232378 196226 232614
rect 196462 232378 196494 232614
rect 195874 232294 196494 232378
rect 195874 232058 195906 232294
rect 196142 232058 196226 232294
rect 196462 232058 196494 232294
rect 195874 214614 196494 232058
rect 195874 214378 195906 214614
rect 196142 214378 196226 214614
rect 196462 214378 196494 214614
rect 195874 214294 196494 214378
rect 195874 214058 195906 214294
rect 196142 214058 196226 214294
rect 196462 214058 196494 214294
rect 195874 196614 196494 214058
rect 195874 196378 195906 196614
rect 196142 196378 196226 196614
rect 196462 196378 196494 196614
rect 195874 196294 196494 196378
rect 195874 196058 195906 196294
rect 196142 196058 196226 196294
rect 196462 196058 196494 196294
rect 195874 178614 196494 196058
rect 195874 178378 195906 178614
rect 196142 178378 196226 178614
rect 196462 178378 196494 178614
rect 195874 178294 196494 178378
rect 195874 178058 195906 178294
rect 196142 178058 196226 178294
rect 196462 178058 196494 178294
rect 195874 160614 196494 178058
rect 195874 160378 195906 160614
rect 196142 160378 196226 160614
rect 196462 160378 196494 160614
rect 195874 160294 196494 160378
rect 195874 160058 195906 160294
rect 196142 160058 196226 160294
rect 196462 160058 196494 160294
rect 195874 142614 196494 160058
rect 195874 142378 195906 142614
rect 196142 142378 196226 142614
rect 196462 142378 196494 142614
rect 195874 142294 196494 142378
rect 195874 142058 195906 142294
rect 196142 142058 196226 142294
rect 196462 142058 196494 142294
rect 195874 124614 196494 142058
rect 195874 124378 195906 124614
rect 196142 124378 196226 124614
rect 196462 124378 196494 124614
rect 195874 124294 196494 124378
rect 195874 124058 195906 124294
rect 196142 124058 196226 124294
rect 196462 124058 196494 124294
rect 195874 106614 196494 124058
rect 195874 106378 195906 106614
rect 196142 106378 196226 106614
rect 196462 106378 196494 106614
rect 195874 106294 196494 106378
rect 195874 106058 195906 106294
rect 196142 106058 196226 106294
rect 196462 106058 196494 106294
rect 195874 88614 196494 106058
rect 195874 88378 195906 88614
rect 196142 88378 196226 88614
rect 196462 88378 196494 88614
rect 195874 88294 196494 88378
rect 195874 88058 195906 88294
rect 196142 88058 196226 88294
rect 196462 88058 196494 88294
rect 195874 70614 196494 88058
rect 195874 70378 195906 70614
rect 196142 70378 196226 70614
rect 196462 70378 196494 70614
rect 195874 70294 196494 70378
rect 195874 70058 195906 70294
rect 196142 70058 196226 70294
rect 196462 70058 196494 70294
rect 195874 52614 196494 70058
rect 195874 52378 195906 52614
rect 196142 52378 196226 52614
rect 196462 52378 196494 52614
rect 195874 52294 196494 52378
rect 195874 52058 195906 52294
rect 196142 52058 196226 52294
rect 196462 52058 196494 52294
rect 195874 34614 196494 52058
rect 195874 34378 195906 34614
rect 196142 34378 196226 34614
rect 196462 34378 196494 34614
rect 195874 34294 196494 34378
rect 195874 34058 195906 34294
rect 196142 34058 196226 34294
rect 196462 34058 196494 34294
rect 195874 16614 196494 34058
rect 195874 16378 195906 16614
rect 196142 16378 196226 16614
rect 196462 16378 196494 16614
rect 195874 16294 196494 16378
rect 195874 16058 195906 16294
rect 196142 16058 196226 16294
rect 196462 16058 196494 16294
rect 195874 -3736 196494 16058
rect 195874 -3972 195906 -3736
rect 196142 -3972 196226 -3736
rect 196462 -3972 196494 -3736
rect 195874 -4056 196494 -3972
rect 195874 -4292 195906 -4056
rect 196142 -4292 196226 -4056
rect 196462 -4292 196494 -4056
rect 195874 -4324 196494 -4292
rect 202714 461092 203334 464004
rect 202714 460856 202746 461092
rect 202982 460856 203066 461092
rect 203302 460856 203334 461092
rect 202714 460772 203334 460856
rect 202714 460536 202746 460772
rect 202982 460536 203066 460772
rect 203302 460536 203334 460772
rect 202714 455454 203334 460536
rect 202714 455218 202746 455454
rect 202982 455218 203066 455454
rect 203302 455218 203334 455454
rect 202714 455134 203334 455218
rect 202714 454898 202746 455134
rect 202982 454898 203066 455134
rect 203302 454898 203334 455134
rect 202714 437454 203334 454898
rect 202714 437218 202746 437454
rect 202982 437218 203066 437454
rect 203302 437218 203334 437454
rect 202714 437134 203334 437218
rect 202714 436898 202746 437134
rect 202982 436898 203066 437134
rect 203302 436898 203334 437134
rect 202714 419454 203334 436898
rect 202714 419218 202746 419454
rect 202982 419218 203066 419454
rect 203302 419218 203334 419454
rect 202714 419134 203334 419218
rect 202714 418898 202746 419134
rect 202982 418898 203066 419134
rect 203302 418898 203334 419134
rect 202714 401454 203334 418898
rect 202714 401218 202746 401454
rect 202982 401218 203066 401454
rect 203302 401218 203334 401454
rect 202714 401134 203334 401218
rect 202714 400898 202746 401134
rect 202982 400898 203066 401134
rect 203302 400898 203334 401134
rect 202714 383454 203334 400898
rect 202714 383218 202746 383454
rect 202982 383218 203066 383454
rect 203302 383218 203334 383454
rect 202714 383134 203334 383218
rect 202714 382898 202746 383134
rect 202982 382898 203066 383134
rect 203302 382898 203334 383134
rect 202714 365454 203334 382898
rect 202714 365218 202746 365454
rect 202982 365218 203066 365454
rect 203302 365218 203334 365454
rect 202714 365134 203334 365218
rect 202714 364898 202746 365134
rect 202982 364898 203066 365134
rect 203302 364898 203334 365134
rect 202714 347454 203334 364898
rect 202714 347218 202746 347454
rect 202982 347218 203066 347454
rect 203302 347218 203334 347454
rect 202714 347134 203334 347218
rect 202714 346898 202746 347134
rect 202982 346898 203066 347134
rect 203302 346898 203334 347134
rect 202714 329454 203334 346898
rect 202714 329218 202746 329454
rect 202982 329218 203066 329454
rect 203302 329218 203334 329454
rect 202714 329134 203334 329218
rect 202714 328898 202746 329134
rect 202982 328898 203066 329134
rect 203302 328898 203334 329134
rect 202714 311454 203334 328898
rect 202714 311218 202746 311454
rect 202982 311218 203066 311454
rect 203302 311218 203334 311454
rect 202714 311134 203334 311218
rect 202714 310898 202746 311134
rect 202982 310898 203066 311134
rect 203302 310898 203334 311134
rect 202714 293454 203334 310898
rect 202714 293218 202746 293454
rect 202982 293218 203066 293454
rect 203302 293218 203334 293454
rect 202714 293134 203334 293218
rect 202714 292898 202746 293134
rect 202982 292898 203066 293134
rect 203302 292898 203334 293134
rect 202714 275454 203334 292898
rect 202714 275218 202746 275454
rect 202982 275218 203066 275454
rect 203302 275218 203334 275454
rect 202714 275134 203334 275218
rect 202714 274898 202746 275134
rect 202982 274898 203066 275134
rect 203302 274898 203334 275134
rect 202714 257454 203334 274898
rect 202714 257218 202746 257454
rect 202982 257218 203066 257454
rect 203302 257218 203334 257454
rect 202714 257134 203334 257218
rect 202714 256898 202746 257134
rect 202982 256898 203066 257134
rect 203302 256898 203334 257134
rect 202714 239454 203334 256898
rect 202714 239218 202746 239454
rect 202982 239218 203066 239454
rect 203302 239218 203334 239454
rect 202714 239134 203334 239218
rect 202714 238898 202746 239134
rect 202982 238898 203066 239134
rect 203302 238898 203334 239134
rect 202714 221454 203334 238898
rect 202714 221218 202746 221454
rect 202982 221218 203066 221454
rect 203302 221218 203334 221454
rect 202714 221134 203334 221218
rect 202714 220898 202746 221134
rect 202982 220898 203066 221134
rect 203302 220898 203334 221134
rect 202714 203454 203334 220898
rect 202714 203218 202746 203454
rect 202982 203218 203066 203454
rect 203302 203218 203334 203454
rect 202714 203134 203334 203218
rect 202714 202898 202746 203134
rect 202982 202898 203066 203134
rect 203302 202898 203334 203134
rect 202714 185454 203334 202898
rect 202714 185218 202746 185454
rect 202982 185218 203066 185454
rect 203302 185218 203334 185454
rect 202714 185134 203334 185218
rect 202714 184898 202746 185134
rect 202982 184898 203066 185134
rect 203302 184898 203334 185134
rect 202714 167454 203334 184898
rect 202714 167218 202746 167454
rect 202982 167218 203066 167454
rect 203302 167218 203334 167454
rect 202714 167134 203334 167218
rect 202714 166898 202746 167134
rect 202982 166898 203066 167134
rect 203302 166898 203334 167134
rect 202714 149454 203334 166898
rect 202714 149218 202746 149454
rect 202982 149218 203066 149454
rect 203302 149218 203334 149454
rect 202714 149134 203334 149218
rect 202714 148898 202746 149134
rect 202982 148898 203066 149134
rect 203302 148898 203334 149134
rect 202714 131454 203334 148898
rect 202714 131218 202746 131454
rect 202982 131218 203066 131454
rect 203302 131218 203334 131454
rect 202714 131134 203334 131218
rect 202714 130898 202746 131134
rect 202982 130898 203066 131134
rect 203302 130898 203334 131134
rect 202714 113454 203334 130898
rect 202714 113218 202746 113454
rect 202982 113218 203066 113454
rect 203302 113218 203334 113454
rect 202714 113134 203334 113218
rect 202714 112898 202746 113134
rect 202982 112898 203066 113134
rect 203302 112898 203334 113134
rect 202714 95454 203334 112898
rect 202714 95218 202746 95454
rect 202982 95218 203066 95454
rect 203302 95218 203334 95454
rect 202714 95134 203334 95218
rect 202714 94898 202746 95134
rect 202982 94898 203066 95134
rect 203302 94898 203334 95134
rect 202714 77454 203334 94898
rect 202714 77218 202746 77454
rect 202982 77218 203066 77454
rect 203302 77218 203334 77454
rect 202714 77134 203334 77218
rect 202714 76898 202746 77134
rect 202982 76898 203066 77134
rect 203302 76898 203334 77134
rect 202714 59454 203334 76898
rect 202714 59218 202746 59454
rect 202982 59218 203066 59454
rect 203302 59218 203334 59454
rect 202714 59134 203334 59218
rect 202714 58898 202746 59134
rect 202982 58898 203066 59134
rect 203302 58898 203334 59134
rect 202714 41454 203334 58898
rect 202714 41218 202746 41454
rect 202982 41218 203066 41454
rect 203302 41218 203334 41454
rect 202714 41134 203334 41218
rect 202714 40898 202746 41134
rect 202982 40898 203066 41134
rect 203302 40898 203334 41134
rect 202714 23454 203334 40898
rect 202714 23218 202746 23454
rect 202982 23218 203066 23454
rect 203302 23218 203334 23454
rect 202714 23134 203334 23218
rect 202714 22898 202746 23134
rect 202982 22898 203066 23134
rect 203302 22898 203334 23134
rect 202714 5454 203334 22898
rect 202714 5218 202746 5454
rect 202982 5218 203066 5454
rect 203302 5218 203334 5454
rect 202714 5134 203334 5218
rect 202714 4898 202746 5134
rect 202982 4898 203066 5134
rect 203302 4898 203334 5134
rect 202714 -856 203334 4898
rect 202714 -1092 202746 -856
rect 202982 -1092 203066 -856
rect 203302 -1092 203334 -856
rect 202714 -1176 203334 -1092
rect 202714 -1412 202746 -1176
rect 202982 -1412 203066 -1176
rect 203302 -1412 203334 -1176
rect 202714 -4324 203334 -1412
rect 206434 462052 207054 464004
rect 206434 461816 206466 462052
rect 206702 461816 206786 462052
rect 207022 461816 207054 462052
rect 206434 461732 207054 461816
rect 206434 461496 206466 461732
rect 206702 461496 206786 461732
rect 207022 461496 207054 461732
rect 206434 441174 207054 461496
rect 206434 440938 206466 441174
rect 206702 440938 206786 441174
rect 207022 440938 207054 441174
rect 206434 440854 207054 440938
rect 206434 440618 206466 440854
rect 206702 440618 206786 440854
rect 207022 440618 207054 440854
rect 206434 423174 207054 440618
rect 206434 422938 206466 423174
rect 206702 422938 206786 423174
rect 207022 422938 207054 423174
rect 206434 422854 207054 422938
rect 206434 422618 206466 422854
rect 206702 422618 206786 422854
rect 207022 422618 207054 422854
rect 206434 405174 207054 422618
rect 206434 404938 206466 405174
rect 206702 404938 206786 405174
rect 207022 404938 207054 405174
rect 206434 404854 207054 404938
rect 206434 404618 206466 404854
rect 206702 404618 206786 404854
rect 207022 404618 207054 404854
rect 206434 387174 207054 404618
rect 206434 386938 206466 387174
rect 206702 386938 206786 387174
rect 207022 386938 207054 387174
rect 206434 386854 207054 386938
rect 206434 386618 206466 386854
rect 206702 386618 206786 386854
rect 207022 386618 207054 386854
rect 206434 369174 207054 386618
rect 206434 368938 206466 369174
rect 206702 368938 206786 369174
rect 207022 368938 207054 369174
rect 206434 368854 207054 368938
rect 206434 368618 206466 368854
rect 206702 368618 206786 368854
rect 207022 368618 207054 368854
rect 206434 351174 207054 368618
rect 206434 350938 206466 351174
rect 206702 350938 206786 351174
rect 207022 350938 207054 351174
rect 206434 350854 207054 350938
rect 206434 350618 206466 350854
rect 206702 350618 206786 350854
rect 207022 350618 207054 350854
rect 206434 333174 207054 350618
rect 206434 332938 206466 333174
rect 206702 332938 206786 333174
rect 207022 332938 207054 333174
rect 206434 332854 207054 332938
rect 206434 332618 206466 332854
rect 206702 332618 206786 332854
rect 207022 332618 207054 332854
rect 206434 315174 207054 332618
rect 206434 314938 206466 315174
rect 206702 314938 206786 315174
rect 207022 314938 207054 315174
rect 206434 314854 207054 314938
rect 206434 314618 206466 314854
rect 206702 314618 206786 314854
rect 207022 314618 207054 314854
rect 206434 297174 207054 314618
rect 206434 296938 206466 297174
rect 206702 296938 206786 297174
rect 207022 296938 207054 297174
rect 206434 296854 207054 296938
rect 206434 296618 206466 296854
rect 206702 296618 206786 296854
rect 207022 296618 207054 296854
rect 206434 279174 207054 296618
rect 206434 278938 206466 279174
rect 206702 278938 206786 279174
rect 207022 278938 207054 279174
rect 206434 278854 207054 278938
rect 206434 278618 206466 278854
rect 206702 278618 206786 278854
rect 207022 278618 207054 278854
rect 206434 261174 207054 278618
rect 206434 260938 206466 261174
rect 206702 260938 206786 261174
rect 207022 260938 207054 261174
rect 206434 260854 207054 260938
rect 206434 260618 206466 260854
rect 206702 260618 206786 260854
rect 207022 260618 207054 260854
rect 206434 243174 207054 260618
rect 206434 242938 206466 243174
rect 206702 242938 206786 243174
rect 207022 242938 207054 243174
rect 206434 242854 207054 242938
rect 206434 242618 206466 242854
rect 206702 242618 206786 242854
rect 207022 242618 207054 242854
rect 206434 225174 207054 242618
rect 206434 224938 206466 225174
rect 206702 224938 206786 225174
rect 207022 224938 207054 225174
rect 206434 224854 207054 224938
rect 206434 224618 206466 224854
rect 206702 224618 206786 224854
rect 207022 224618 207054 224854
rect 206434 207174 207054 224618
rect 206434 206938 206466 207174
rect 206702 206938 206786 207174
rect 207022 206938 207054 207174
rect 206434 206854 207054 206938
rect 206434 206618 206466 206854
rect 206702 206618 206786 206854
rect 207022 206618 207054 206854
rect 206434 189174 207054 206618
rect 206434 188938 206466 189174
rect 206702 188938 206786 189174
rect 207022 188938 207054 189174
rect 206434 188854 207054 188938
rect 206434 188618 206466 188854
rect 206702 188618 206786 188854
rect 207022 188618 207054 188854
rect 206434 171174 207054 188618
rect 206434 170938 206466 171174
rect 206702 170938 206786 171174
rect 207022 170938 207054 171174
rect 206434 170854 207054 170938
rect 206434 170618 206466 170854
rect 206702 170618 206786 170854
rect 207022 170618 207054 170854
rect 206434 153174 207054 170618
rect 206434 152938 206466 153174
rect 206702 152938 206786 153174
rect 207022 152938 207054 153174
rect 206434 152854 207054 152938
rect 206434 152618 206466 152854
rect 206702 152618 206786 152854
rect 207022 152618 207054 152854
rect 206434 135174 207054 152618
rect 206434 134938 206466 135174
rect 206702 134938 206786 135174
rect 207022 134938 207054 135174
rect 206434 134854 207054 134938
rect 206434 134618 206466 134854
rect 206702 134618 206786 134854
rect 207022 134618 207054 134854
rect 206434 117174 207054 134618
rect 206434 116938 206466 117174
rect 206702 116938 206786 117174
rect 207022 116938 207054 117174
rect 206434 116854 207054 116938
rect 206434 116618 206466 116854
rect 206702 116618 206786 116854
rect 207022 116618 207054 116854
rect 206434 99174 207054 116618
rect 206434 98938 206466 99174
rect 206702 98938 206786 99174
rect 207022 98938 207054 99174
rect 206434 98854 207054 98938
rect 206434 98618 206466 98854
rect 206702 98618 206786 98854
rect 207022 98618 207054 98854
rect 206434 81174 207054 98618
rect 206434 80938 206466 81174
rect 206702 80938 206786 81174
rect 207022 80938 207054 81174
rect 206434 80854 207054 80938
rect 206434 80618 206466 80854
rect 206702 80618 206786 80854
rect 207022 80618 207054 80854
rect 206434 63174 207054 80618
rect 206434 62938 206466 63174
rect 206702 62938 206786 63174
rect 207022 62938 207054 63174
rect 206434 62854 207054 62938
rect 206434 62618 206466 62854
rect 206702 62618 206786 62854
rect 207022 62618 207054 62854
rect 206434 45174 207054 62618
rect 206434 44938 206466 45174
rect 206702 44938 206786 45174
rect 207022 44938 207054 45174
rect 206434 44854 207054 44938
rect 206434 44618 206466 44854
rect 206702 44618 206786 44854
rect 207022 44618 207054 44854
rect 206434 27174 207054 44618
rect 206434 26938 206466 27174
rect 206702 26938 206786 27174
rect 207022 26938 207054 27174
rect 206434 26854 207054 26938
rect 206434 26618 206466 26854
rect 206702 26618 206786 26854
rect 207022 26618 207054 26854
rect 206434 9174 207054 26618
rect 206434 8938 206466 9174
rect 206702 8938 206786 9174
rect 207022 8938 207054 9174
rect 206434 8854 207054 8938
rect 206434 8618 206466 8854
rect 206702 8618 206786 8854
rect 207022 8618 207054 8854
rect 206434 -1816 207054 8618
rect 206434 -2052 206466 -1816
rect 206702 -2052 206786 -1816
rect 207022 -2052 207054 -1816
rect 206434 -2136 207054 -2052
rect 206434 -2372 206466 -2136
rect 206702 -2372 206786 -2136
rect 207022 -2372 207054 -2136
rect 206434 -4324 207054 -2372
rect 210154 463012 210774 464004
rect 210154 462776 210186 463012
rect 210422 462776 210506 463012
rect 210742 462776 210774 463012
rect 210154 462692 210774 462776
rect 210154 462456 210186 462692
rect 210422 462456 210506 462692
rect 210742 462456 210774 462692
rect 210154 444894 210774 462456
rect 210154 444658 210186 444894
rect 210422 444658 210506 444894
rect 210742 444658 210774 444894
rect 210154 444574 210774 444658
rect 210154 444338 210186 444574
rect 210422 444338 210506 444574
rect 210742 444338 210774 444574
rect 210154 426894 210774 444338
rect 210154 426658 210186 426894
rect 210422 426658 210506 426894
rect 210742 426658 210774 426894
rect 210154 426574 210774 426658
rect 210154 426338 210186 426574
rect 210422 426338 210506 426574
rect 210742 426338 210774 426574
rect 210154 408894 210774 426338
rect 210154 408658 210186 408894
rect 210422 408658 210506 408894
rect 210742 408658 210774 408894
rect 210154 408574 210774 408658
rect 210154 408338 210186 408574
rect 210422 408338 210506 408574
rect 210742 408338 210774 408574
rect 210154 390894 210774 408338
rect 210154 390658 210186 390894
rect 210422 390658 210506 390894
rect 210742 390658 210774 390894
rect 210154 390574 210774 390658
rect 210154 390338 210186 390574
rect 210422 390338 210506 390574
rect 210742 390338 210774 390574
rect 210154 372894 210774 390338
rect 210154 372658 210186 372894
rect 210422 372658 210506 372894
rect 210742 372658 210774 372894
rect 210154 372574 210774 372658
rect 210154 372338 210186 372574
rect 210422 372338 210506 372574
rect 210742 372338 210774 372574
rect 210154 354894 210774 372338
rect 210154 354658 210186 354894
rect 210422 354658 210506 354894
rect 210742 354658 210774 354894
rect 210154 354574 210774 354658
rect 210154 354338 210186 354574
rect 210422 354338 210506 354574
rect 210742 354338 210774 354574
rect 210154 336894 210774 354338
rect 210154 336658 210186 336894
rect 210422 336658 210506 336894
rect 210742 336658 210774 336894
rect 210154 336574 210774 336658
rect 210154 336338 210186 336574
rect 210422 336338 210506 336574
rect 210742 336338 210774 336574
rect 210154 318894 210774 336338
rect 210154 318658 210186 318894
rect 210422 318658 210506 318894
rect 210742 318658 210774 318894
rect 210154 318574 210774 318658
rect 210154 318338 210186 318574
rect 210422 318338 210506 318574
rect 210742 318338 210774 318574
rect 210154 300894 210774 318338
rect 210154 300658 210186 300894
rect 210422 300658 210506 300894
rect 210742 300658 210774 300894
rect 210154 300574 210774 300658
rect 210154 300338 210186 300574
rect 210422 300338 210506 300574
rect 210742 300338 210774 300574
rect 210154 282894 210774 300338
rect 210154 282658 210186 282894
rect 210422 282658 210506 282894
rect 210742 282658 210774 282894
rect 210154 282574 210774 282658
rect 210154 282338 210186 282574
rect 210422 282338 210506 282574
rect 210742 282338 210774 282574
rect 210154 264894 210774 282338
rect 210154 264658 210186 264894
rect 210422 264658 210506 264894
rect 210742 264658 210774 264894
rect 210154 264574 210774 264658
rect 210154 264338 210186 264574
rect 210422 264338 210506 264574
rect 210742 264338 210774 264574
rect 210154 246894 210774 264338
rect 210154 246658 210186 246894
rect 210422 246658 210506 246894
rect 210742 246658 210774 246894
rect 210154 246574 210774 246658
rect 210154 246338 210186 246574
rect 210422 246338 210506 246574
rect 210742 246338 210774 246574
rect 210154 228894 210774 246338
rect 210154 228658 210186 228894
rect 210422 228658 210506 228894
rect 210742 228658 210774 228894
rect 210154 228574 210774 228658
rect 210154 228338 210186 228574
rect 210422 228338 210506 228574
rect 210742 228338 210774 228574
rect 210154 210894 210774 228338
rect 210154 210658 210186 210894
rect 210422 210658 210506 210894
rect 210742 210658 210774 210894
rect 210154 210574 210774 210658
rect 210154 210338 210186 210574
rect 210422 210338 210506 210574
rect 210742 210338 210774 210574
rect 210154 192894 210774 210338
rect 210154 192658 210186 192894
rect 210422 192658 210506 192894
rect 210742 192658 210774 192894
rect 210154 192574 210774 192658
rect 210154 192338 210186 192574
rect 210422 192338 210506 192574
rect 210742 192338 210774 192574
rect 210154 174894 210774 192338
rect 210154 174658 210186 174894
rect 210422 174658 210506 174894
rect 210742 174658 210774 174894
rect 210154 174574 210774 174658
rect 210154 174338 210186 174574
rect 210422 174338 210506 174574
rect 210742 174338 210774 174574
rect 210154 156894 210774 174338
rect 210154 156658 210186 156894
rect 210422 156658 210506 156894
rect 210742 156658 210774 156894
rect 210154 156574 210774 156658
rect 210154 156338 210186 156574
rect 210422 156338 210506 156574
rect 210742 156338 210774 156574
rect 210154 138894 210774 156338
rect 210154 138658 210186 138894
rect 210422 138658 210506 138894
rect 210742 138658 210774 138894
rect 210154 138574 210774 138658
rect 210154 138338 210186 138574
rect 210422 138338 210506 138574
rect 210742 138338 210774 138574
rect 210154 120894 210774 138338
rect 210154 120658 210186 120894
rect 210422 120658 210506 120894
rect 210742 120658 210774 120894
rect 210154 120574 210774 120658
rect 210154 120338 210186 120574
rect 210422 120338 210506 120574
rect 210742 120338 210774 120574
rect 210154 102894 210774 120338
rect 210154 102658 210186 102894
rect 210422 102658 210506 102894
rect 210742 102658 210774 102894
rect 210154 102574 210774 102658
rect 210154 102338 210186 102574
rect 210422 102338 210506 102574
rect 210742 102338 210774 102574
rect 210154 84894 210774 102338
rect 210154 84658 210186 84894
rect 210422 84658 210506 84894
rect 210742 84658 210774 84894
rect 210154 84574 210774 84658
rect 210154 84338 210186 84574
rect 210422 84338 210506 84574
rect 210742 84338 210774 84574
rect 210154 66894 210774 84338
rect 210154 66658 210186 66894
rect 210422 66658 210506 66894
rect 210742 66658 210774 66894
rect 210154 66574 210774 66658
rect 210154 66338 210186 66574
rect 210422 66338 210506 66574
rect 210742 66338 210774 66574
rect 210154 48894 210774 66338
rect 210154 48658 210186 48894
rect 210422 48658 210506 48894
rect 210742 48658 210774 48894
rect 210154 48574 210774 48658
rect 210154 48338 210186 48574
rect 210422 48338 210506 48574
rect 210742 48338 210774 48574
rect 210154 30894 210774 48338
rect 210154 30658 210186 30894
rect 210422 30658 210506 30894
rect 210742 30658 210774 30894
rect 210154 30574 210774 30658
rect 210154 30338 210186 30574
rect 210422 30338 210506 30574
rect 210742 30338 210774 30574
rect 210154 12894 210774 30338
rect 210154 12658 210186 12894
rect 210422 12658 210506 12894
rect 210742 12658 210774 12894
rect 210154 12574 210774 12658
rect 210154 12338 210186 12574
rect 210422 12338 210506 12574
rect 210742 12338 210774 12574
rect 210154 -2776 210774 12338
rect 210154 -3012 210186 -2776
rect 210422 -3012 210506 -2776
rect 210742 -3012 210774 -2776
rect 210154 -3096 210774 -3012
rect 210154 -3332 210186 -3096
rect 210422 -3332 210506 -3096
rect 210742 -3332 210774 -3096
rect 210154 -4324 210774 -3332
rect 213874 463972 214494 464004
rect 213874 463736 213906 463972
rect 214142 463736 214226 463972
rect 214462 463736 214494 463972
rect 213874 463652 214494 463736
rect 213874 463416 213906 463652
rect 214142 463416 214226 463652
rect 214462 463416 214494 463652
rect 213874 448614 214494 463416
rect 213874 448378 213906 448614
rect 214142 448378 214226 448614
rect 214462 448378 214494 448614
rect 213874 448294 214494 448378
rect 213874 448058 213906 448294
rect 214142 448058 214226 448294
rect 214462 448058 214494 448294
rect 213874 430614 214494 448058
rect 213874 430378 213906 430614
rect 214142 430378 214226 430614
rect 214462 430378 214494 430614
rect 213874 430294 214494 430378
rect 213874 430058 213906 430294
rect 214142 430058 214226 430294
rect 214462 430058 214494 430294
rect 213874 412614 214494 430058
rect 213874 412378 213906 412614
rect 214142 412378 214226 412614
rect 214462 412378 214494 412614
rect 213874 412294 214494 412378
rect 213874 412058 213906 412294
rect 214142 412058 214226 412294
rect 214462 412058 214494 412294
rect 213874 394614 214494 412058
rect 213874 394378 213906 394614
rect 214142 394378 214226 394614
rect 214462 394378 214494 394614
rect 213874 394294 214494 394378
rect 213874 394058 213906 394294
rect 214142 394058 214226 394294
rect 214462 394058 214494 394294
rect 213874 376614 214494 394058
rect 213874 376378 213906 376614
rect 214142 376378 214226 376614
rect 214462 376378 214494 376614
rect 213874 376294 214494 376378
rect 213874 376058 213906 376294
rect 214142 376058 214226 376294
rect 214462 376058 214494 376294
rect 213874 358614 214494 376058
rect 213874 358378 213906 358614
rect 214142 358378 214226 358614
rect 214462 358378 214494 358614
rect 213874 358294 214494 358378
rect 213874 358058 213906 358294
rect 214142 358058 214226 358294
rect 214462 358058 214494 358294
rect 213874 340614 214494 358058
rect 213874 340378 213906 340614
rect 214142 340378 214226 340614
rect 214462 340378 214494 340614
rect 213874 340294 214494 340378
rect 213874 340058 213906 340294
rect 214142 340058 214226 340294
rect 214462 340058 214494 340294
rect 213874 322614 214494 340058
rect 213874 322378 213906 322614
rect 214142 322378 214226 322614
rect 214462 322378 214494 322614
rect 213874 322294 214494 322378
rect 213874 322058 213906 322294
rect 214142 322058 214226 322294
rect 214462 322058 214494 322294
rect 213874 304614 214494 322058
rect 213874 304378 213906 304614
rect 214142 304378 214226 304614
rect 214462 304378 214494 304614
rect 213874 304294 214494 304378
rect 213874 304058 213906 304294
rect 214142 304058 214226 304294
rect 214462 304058 214494 304294
rect 213874 286614 214494 304058
rect 213874 286378 213906 286614
rect 214142 286378 214226 286614
rect 214462 286378 214494 286614
rect 213874 286294 214494 286378
rect 213874 286058 213906 286294
rect 214142 286058 214226 286294
rect 214462 286058 214494 286294
rect 213874 268614 214494 286058
rect 213874 268378 213906 268614
rect 214142 268378 214226 268614
rect 214462 268378 214494 268614
rect 213874 268294 214494 268378
rect 213874 268058 213906 268294
rect 214142 268058 214226 268294
rect 214462 268058 214494 268294
rect 213874 250614 214494 268058
rect 213874 250378 213906 250614
rect 214142 250378 214226 250614
rect 214462 250378 214494 250614
rect 213874 250294 214494 250378
rect 213874 250058 213906 250294
rect 214142 250058 214226 250294
rect 214462 250058 214494 250294
rect 213874 232614 214494 250058
rect 213874 232378 213906 232614
rect 214142 232378 214226 232614
rect 214462 232378 214494 232614
rect 213874 232294 214494 232378
rect 213874 232058 213906 232294
rect 214142 232058 214226 232294
rect 214462 232058 214494 232294
rect 213874 214614 214494 232058
rect 213874 214378 213906 214614
rect 214142 214378 214226 214614
rect 214462 214378 214494 214614
rect 213874 214294 214494 214378
rect 213874 214058 213906 214294
rect 214142 214058 214226 214294
rect 214462 214058 214494 214294
rect 213874 196614 214494 214058
rect 213874 196378 213906 196614
rect 214142 196378 214226 196614
rect 214462 196378 214494 196614
rect 213874 196294 214494 196378
rect 213874 196058 213906 196294
rect 214142 196058 214226 196294
rect 214462 196058 214494 196294
rect 213874 178614 214494 196058
rect 213874 178378 213906 178614
rect 214142 178378 214226 178614
rect 214462 178378 214494 178614
rect 213874 178294 214494 178378
rect 213874 178058 213906 178294
rect 214142 178058 214226 178294
rect 214462 178058 214494 178294
rect 213874 160614 214494 178058
rect 213874 160378 213906 160614
rect 214142 160378 214226 160614
rect 214462 160378 214494 160614
rect 213874 160294 214494 160378
rect 213874 160058 213906 160294
rect 214142 160058 214226 160294
rect 214462 160058 214494 160294
rect 213874 142614 214494 160058
rect 213874 142378 213906 142614
rect 214142 142378 214226 142614
rect 214462 142378 214494 142614
rect 213874 142294 214494 142378
rect 213874 142058 213906 142294
rect 214142 142058 214226 142294
rect 214462 142058 214494 142294
rect 213874 124614 214494 142058
rect 213874 124378 213906 124614
rect 214142 124378 214226 124614
rect 214462 124378 214494 124614
rect 213874 124294 214494 124378
rect 213874 124058 213906 124294
rect 214142 124058 214226 124294
rect 214462 124058 214494 124294
rect 213874 106614 214494 124058
rect 213874 106378 213906 106614
rect 214142 106378 214226 106614
rect 214462 106378 214494 106614
rect 213874 106294 214494 106378
rect 213874 106058 213906 106294
rect 214142 106058 214226 106294
rect 214462 106058 214494 106294
rect 213874 88614 214494 106058
rect 213874 88378 213906 88614
rect 214142 88378 214226 88614
rect 214462 88378 214494 88614
rect 213874 88294 214494 88378
rect 213874 88058 213906 88294
rect 214142 88058 214226 88294
rect 214462 88058 214494 88294
rect 213874 70614 214494 88058
rect 213874 70378 213906 70614
rect 214142 70378 214226 70614
rect 214462 70378 214494 70614
rect 213874 70294 214494 70378
rect 213874 70058 213906 70294
rect 214142 70058 214226 70294
rect 214462 70058 214494 70294
rect 213874 52614 214494 70058
rect 213874 52378 213906 52614
rect 214142 52378 214226 52614
rect 214462 52378 214494 52614
rect 213874 52294 214494 52378
rect 213874 52058 213906 52294
rect 214142 52058 214226 52294
rect 214462 52058 214494 52294
rect 213874 34614 214494 52058
rect 213874 34378 213906 34614
rect 214142 34378 214226 34614
rect 214462 34378 214494 34614
rect 213874 34294 214494 34378
rect 213874 34058 213906 34294
rect 214142 34058 214226 34294
rect 214462 34058 214494 34294
rect 213874 16614 214494 34058
rect 213874 16378 213906 16614
rect 214142 16378 214226 16614
rect 214462 16378 214494 16614
rect 213874 16294 214494 16378
rect 213874 16058 213906 16294
rect 214142 16058 214226 16294
rect 214462 16058 214494 16294
rect 213874 -3736 214494 16058
rect 213874 -3972 213906 -3736
rect 214142 -3972 214226 -3736
rect 214462 -3972 214494 -3736
rect 213874 -4056 214494 -3972
rect 213874 -4292 213906 -4056
rect 214142 -4292 214226 -4056
rect 214462 -4292 214494 -4056
rect 213874 -4324 214494 -4292
rect 220714 461092 221334 464004
rect 220714 460856 220746 461092
rect 220982 460856 221066 461092
rect 221302 460856 221334 461092
rect 220714 460772 221334 460856
rect 220714 460536 220746 460772
rect 220982 460536 221066 460772
rect 221302 460536 221334 460772
rect 220714 455454 221334 460536
rect 220714 455218 220746 455454
rect 220982 455218 221066 455454
rect 221302 455218 221334 455454
rect 220714 455134 221334 455218
rect 220714 454898 220746 455134
rect 220982 454898 221066 455134
rect 221302 454898 221334 455134
rect 220714 437454 221334 454898
rect 220714 437218 220746 437454
rect 220982 437218 221066 437454
rect 221302 437218 221334 437454
rect 220714 437134 221334 437218
rect 220714 436898 220746 437134
rect 220982 436898 221066 437134
rect 221302 436898 221334 437134
rect 220714 419454 221334 436898
rect 220714 419218 220746 419454
rect 220982 419218 221066 419454
rect 221302 419218 221334 419454
rect 220714 419134 221334 419218
rect 220714 418898 220746 419134
rect 220982 418898 221066 419134
rect 221302 418898 221334 419134
rect 220714 401454 221334 418898
rect 220714 401218 220746 401454
rect 220982 401218 221066 401454
rect 221302 401218 221334 401454
rect 220714 401134 221334 401218
rect 220714 400898 220746 401134
rect 220982 400898 221066 401134
rect 221302 400898 221334 401134
rect 220714 383454 221334 400898
rect 220714 383218 220746 383454
rect 220982 383218 221066 383454
rect 221302 383218 221334 383454
rect 220714 383134 221334 383218
rect 220714 382898 220746 383134
rect 220982 382898 221066 383134
rect 221302 382898 221334 383134
rect 220714 365454 221334 382898
rect 220714 365218 220746 365454
rect 220982 365218 221066 365454
rect 221302 365218 221334 365454
rect 220714 365134 221334 365218
rect 220714 364898 220746 365134
rect 220982 364898 221066 365134
rect 221302 364898 221334 365134
rect 220714 347454 221334 364898
rect 220714 347218 220746 347454
rect 220982 347218 221066 347454
rect 221302 347218 221334 347454
rect 220714 347134 221334 347218
rect 220714 346898 220746 347134
rect 220982 346898 221066 347134
rect 221302 346898 221334 347134
rect 220714 329454 221334 346898
rect 220714 329218 220746 329454
rect 220982 329218 221066 329454
rect 221302 329218 221334 329454
rect 220714 329134 221334 329218
rect 220714 328898 220746 329134
rect 220982 328898 221066 329134
rect 221302 328898 221334 329134
rect 220714 311454 221334 328898
rect 220714 311218 220746 311454
rect 220982 311218 221066 311454
rect 221302 311218 221334 311454
rect 220714 311134 221334 311218
rect 220714 310898 220746 311134
rect 220982 310898 221066 311134
rect 221302 310898 221334 311134
rect 220714 293454 221334 310898
rect 220714 293218 220746 293454
rect 220982 293218 221066 293454
rect 221302 293218 221334 293454
rect 220714 293134 221334 293218
rect 220714 292898 220746 293134
rect 220982 292898 221066 293134
rect 221302 292898 221334 293134
rect 220714 275454 221334 292898
rect 220714 275218 220746 275454
rect 220982 275218 221066 275454
rect 221302 275218 221334 275454
rect 220714 275134 221334 275218
rect 220714 274898 220746 275134
rect 220982 274898 221066 275134
rect 221302 274898 221334 275134
rect 220714 257454 221334 274898
rect 220714 257218 220746 257454
rect 220982 257218 221066 257454
rect 221302 257218 221334 257454
rect 220714 257134 221334 257218
rect 220714 256898 220746 257134
rect 220982 256898 221066 257134
rect 221302 256898 221334 257134
rect 220714 239454 221334 256898
rect 220714 239218 220746 239454
rect 220982 239218 221066 239454
rect 221302 239218 221334 239454
rect 220714 239134 221334 239218
rect 220714 238898 220746 239134
rect 220982 238898 221066 239134
rect 221302 238898 221334 239134
rect 220714 221454 221334 238898
rect 220714 221218 220746 221454
rect 220982 221218 221066 221454
rect 221302 221218 221334 221454
rect 220714 221134 221334 221218
rect 220714 220898 220746 221134
rect 220982 220898 221066 221134
rect 221302 220898 221334 221134
rect 220714 203454 221334 220898
rect 220714 203218 220746 203454
rect 220982 203218 221066 203454
rect 221302 203218 221334 203454
rect 220714 203134 221334 203218
rect 220714 202898 220746 203134
rect 220982 202898 221066 203134
rect 221302 202898 221334 203134
rect 220714 185454 221334 202898
rect 220714 185218 220746 185454
rect 220982 185218 221066 185454
rect 221302 185218 221334 185454
rect 220714 185134 221334 185218
rect 220714 184898 220746 185134
rect 220982 184898 221066 185134
rect 221302 184898 221334 185134
rect 220714 167454 221334 184898
rect 220714 167218 220746 167454
rect 220982 167218 221066 167454
rect 221302 167218 221334 167454
rect 220714 167134 221334 167218
rect 220714 166898 220746 167134
rect 220982 166898 221066 167134
rect 221302 166898 221334 167134
rect 220714 149454 221334 166898
rect 220714 149218 220746 149454
rect 220982 149218 221066 149454
rect 221302 149218 221334 149454
rect 220714 149134 221334 149218
rect 220714 148898 220746 149134
rect 220982 148898 221066 149134
rect 221302 148898 221334 149134
rect 220714 131454 221334 148898
rect 220714 131218 220746 131454
rect 220982 131218 221066 131454
rect 221302 131218 221334 131454
rect 220714 131134 221334 131218
rect 220714 130898 220746 131134
rect 220982 130898 221066 131134
rect 221302 130898 221334 131134
rect 220714 113454 221334 130898
rect 220714 113218 220746 113454
rect 220982 113218 221066 113454
rect 221302 113218 221334 113454
rect 220714 113134 221334 113218
rect 220714 112898 220746 113134
rect 220982 112898 221066 113134
rect 221302 112898 221334 113134
rect 220714 95454 221334 112898
rect 220714 95218 220746 95454
rect 220982 95218 221066 95454
rect 221302 95218 221334 95454
rect 220714 95134 221334 95218
rect 220714 94898 220746 95134
rect 220982 94898 221066 95134
rect 221302 94898 221334 95134
rect 220714 77454 221334 94898
rect 220714 77218 220746 77454
rect 220982 77218 221066 77454
rect 221302 77218 221334 77454
rect 220714 77134 221334 77218
rect 220714 76898 220746 77134
rect 220982 76898 221066 77134
rect 221302 76898 221334 77134
rect 220714 59454 221334 76898
rect 220714 59218 220746 59454
rect 220982 59218 221066 59454
rect 221302 59218 221334 59454
rect 220714 59134 221334 59218
rect 220714 58898 220746 59134
rect 220982 58898 221066 59134
rect 221302 58898 221334 59134
rect 220714 41454 221334 58898
rect 220714 41218 220746 41454
rect 220982 41218 221066 41454
rect 221302 41218 221334 41454
rect 220714 41134 221334 41218
rect 220714 40898 220746 41134
rect 220982 40898 221066 41134
rect 221302 40898 221334 41134
rect 220714 23454 221334 40898
rect 220714 23218 220746 23454
rect 220982 23218 221066 23454
rect 221302 23218 221334 23454
rect 220714 23134 221334 23218
rect 220714 22898 220746 23134
rect 220982 22898 221066 23134
rect 221302 22898 221334 23134
rect 220714 5454 221334 22898
rect 220714 5218 220746 5454
rect 220982 5218 221066 5454
rect 221302 5218 221334 5454
rect 220714 5134 221334 5218
rect 220714 4898 220746 5134
rect 220982 4898 221066 5134
rect 221302 4898 221334 5134
rect 220714 -856 221334 4898
rect 220714 -1092 220746 -856
rect 220982 -1092 221066 -856
rect 221302 -1092 221334 -856
rect 220714 -1176 221334 -1092
rect 220714 -1412 220746 -1176
rect 220982 -1412 221066 -1176
rect 221302 -1412 221334 -1176
rect 220714 -4324 221334 -1412
rect 224434 462052 225054 464004
rect 224434 461816 224466 462052
rect 224702 461816 224786 462052
rect 225022 461816 225054 462052
rect 224434 461732 225054 461816
rect 224434 461496 224466 461732
rect 224702 461496 224786 461732
rect 225022 461496 225054 461732
rect 224434 441174 225054 461496
rect 224434 440938 224466 441174
rect 224702 440938 224786 441174
rect 225022 440938 225054 441174
rect 224434 440854 225054 440938
rect 224434 440618 224466 440854
rect 224702 440618 224786 440854
rect 225022 440618 225054 440854
rect 224434 423174 225054 440618
rect 224434 422938 224466 423174
rect 224702 422938 224786 423174
rect 225022 422938 225054 423174
rect 224434 422854 225054 422938
rect 224434 422618 224466 422854
rect 224702 422618 224786 422854
rect 225022 422618 225054 422854
rect 224434 405174 225054 422618
rect 224434 404938 224466 405174
rect 224702 404938 224786 405174
rect 225022 404938 225054 405174
rect 224434 404854 225054 404938
rect 224434 404618 224466 404854
rect 224702 404618 224786 404854
rect 225022 404618 225054 404854
rect 224434 387174 225054 404618
rect 224434 386938 224466 387174
rect 224702 386938 224786 387174
rect 225022 386938 225054 387174
rect 224434 386854 225054 386938
rect 224434 386618 224466 386854
rect 224702 386618 224786 386854
rect 225022 386618 225054 386854
rect 224434 369174 225054 386618
rect 224434 368938 224466 369174
rect 224702 368938 224786 369174
rect 225022 368938 225054 369174
rect 224434 368854 225054 368938
rect 224434 368618 224466 368854
rect 224702 368618 224786 368854
rect 225022 368618 225054 368854
rect 224434 351174 225054 368618
rect 224434 350938 224466 351174
rect 224702 350938 224786 351174
rect 225022 350938 225054 351174
rect 224434 350854 225054 350938
rect 224434 350618 224466 350854
rect 224702 350618 224786 350854
rect 225022 350618 225054 350854
rect 224434 333174 225054 350618
rect 224434 332938 224466 333174
rect 224702 332938 224786 333174
rect 225022 332938 225054 333174
rect 224434 332854 225054 332938
rect 224434 332618 224466 332854
rect 224702 332618 224786 332854
rect 225022 332618 225054 332854
rect 224434 315174 225054 332618
rect 224434 314938 224466 315174
rect 224702 314938 224786 315174
rect 225022 314938 225054 315174
rect 224434 314854 225054 314938
rect 224434 314618 224466 314854
rect 224702 314618 224786 314854
rect 225022 314618 225054 314854
rect 224434 297174 225054 314618
rect 224434 296938 224466 297174
rect 224702 296938 224786 297174
rect 225022 296938 225054 297174
rect 224434 296854 225054 296938
rect 224434 296618 224466 296854
rect 224702 296618 224786 296854
rect 225022 296618 225054 296854
rect 224434 279174 225054 296618
rect 224434 278938 224466 279174
rect 224702 278938 224786 279174
rect 225022 278938 225054 279174
rect 224434 278854 225054 278938
rect 224434 278618 224466 278854
rect 224702 278618 224786 278854
rect 225022 278618 225054 278854
rect 224434 261174 225054 278618
rect 224434 260938 224466 261174
rect 224702 260938 224786 261174
rect 225022 260938 225054 261174
rect 224434 260854 225054 260938
rect 224434 260618 224466 260854
rect 224702 260618 224786 260854
rect 225022 260618 225054 260854
rect 224434 243174 225054 260618
rect 224434 242938 224466 243174
rect 224702 242938 224786 243174
rect 225022 242938 225054 243174
rect 224434 242854 225054 242938
rect 224434 242618 224466 242854
rect 224702 242618 224786 242854
rect 225022 242618 225054 242854
rect 224434 225174 225054 242618
rect 224434 224938 224466 225174
rect 224702 224938 224786 225174
rect 225022 224938 225054 225174
rect 224434 224854 225054 224938
rect 224434 224618 224466 224854
rect 224702 224618 224786 224854
rect 225022 224618 225054 224854
rect 224434 207174 225054 224618
rect 224434 206938 224466 207174
rect 224702 206938 224786 207174
rect 225022 206938 225054 207174
rect 224434 206854 225054 206938
rect 224434 206618 224466 206854
rect 224702 206618 224786 206854
rect 225022 206618 225054 206854
rect 224434 189174 225054 206618
rect 224434 188938 224466 189174
rect 224702 188938 224786 189174
rect 225022 188938 225054 189174
rect 224434 188854 225054 188938
rect 224434 188618 224466 188854
rect 224702 188618 224786 188854
rect 225022 188618 225054 188854
rect 224434 171174 225054 188618
rect 224434 170938 224466 171174
rect 224702 170938 224786 171174
rect 225022 170938 225054 171174
rect 224434 170854 225054 170938
rect 224434 170618 224466 170854
rect 224702 170618 224786 170854
rect 225022 170618 225054 170854
rect 224434 153174 225054 170618
rect 224434 152938 224466 153174
rect 224702 152938 224786 153174
rect 225022 152938 225054 153174
rect 224434 152854 225054 152938
rect 224434 152618 224466 152854
rect 224702 152618 224786 152854
rect 225022 152618 225054 152854
rect 224434 135174 225054 152618
rect 224434 134938 224466 135174
rect 224702 134938 224786 135174
rect 225022 134938 225054 135174
rect 224434 134854 225054 134938
rect 224434 134618 224466 134854
rect 224702 134618 224786 134854
rect 225022 134618 225054 134854
rect 224434 117174 225054 134618
rect 224434 116938 224466 117174
rect 224702 116938 224786 117174
rect 225022 116938 225054 117174
rect 224434 116854 225054 116938
rect 224434 116618 224466 116854
rect 224702 116618 224786 116854
rect 225022 116618 225054 116854
rect 224434 99174 225054 116618
rect 224434 98938 224466 99174
rect 224702 98938 224786 99174
rect 225022 98938 225054 99174
rect 224434 98854 225054 98938
rect 224434 98618 224466 98854
rect 224702 98618 224786 98854
rect 225022 98618 225054 98854
rect 224434 81174 225054 98618
rect 224434 80938 224466 81174
rect 224702 80938 224786 81174
rect 225022 80938 225054 81174
rect 224434 80854 225054 80938
rect 224434 80618 224466 80854
rect 224702 80618 224786 80854
rect 225022 80618 225054 80854
rect 224434 63174 225054 80618
rect 224434 62938 224466 63174
rect 224702 62938 224786 63174
rect 225022 62938 225054 63174
rect 224434 62854 225054 62938
rect 224434 62618 224466 62854
rect 224702 62618 224786 62854
rect 225022 62618 225054 62854
rect 224434 45174 225054 62618
rect 224434 44938 224466 45174
rect 224702 44938 224786 45174
rect 225022 44938 225054 45174
rect 224434 44854 225054 44938
rect 224434 44618 224466 44854
rect 224702 44618 224786 44854
rect 225022 44618 225054 44854
rect 224434 27174 225054 44618
rect 224434 26938 224466 27174
rect 224702 26938 224786 27174
rect 225022 26938 225054 27174
rect 224434 26854 225054 26938
rect 224434 26618 224466 26854
rect 224702 26618 224786 26854
rect 225022 26618 225054 26854
rect 224434 9174 225054 26618
rect 224434 8938 224466 9174
rect 224702 8938 224786 9174
rect 225022 8938 225054 9174
rect 224434 8854 225054 8938
rect 224434 8618 224466 8854
rect 224702 8618 224786 8854
rect 225022 8618 225054 8854
rect 224434 -1816 225054 8618
rect 224434 -2052 224466 -1816
rect 224702 -2052 224786 -1816
rect 225022 -2052 225054 -1816
rect 224434 -2136 225054 -2052
rect 224434 -2372 224466 -2136
rect 224702 -2372 224786 -2136
rect 225022 -2372 225054 -2136
rect 224434 -4324 225054 -2372
rect 228154 463012 228774 464004
rect 228154 462776 228186 463012
rect 228422 462776 228506 463012
rect 228742 462776 228774 463012
rect 228154 462692 228774 462776
rect 228154 462456 228186 462692
rect 228422 462456 228506 462692
rect 228742 462456 228774 462692
rect 228154 444894 228774 462456
rect 228154 444658 228186 444894
rect 228422 444658 228506 444894
rect 228742 444658 228774 444894
rect 228154 444574 228774 444658
rect 228154 444338 228186 444574
rect 228422 444338 228506 444574
rect 228742 444338 228774 444574
rect 228154 426894 228774 444338
rect 228154 426658 228186 426894
rect 228422 426658 228506 426894
rect 228742 426658 228774 426894
rect 228154 426574 228774 426658
rect 228154 426338 228186 426574
rect 228422 426338 228506 426574
rect 228742 426338 228774 426574
rect 228154 408894 228774 426338
rect 228154 408658 228186 408894
rect 228422 408658 228506 408894
rect 228742 408658 228774 408894
rect 228154 408574 228774 408658
rect 228154 408338 228186 408574
rect 228422 408338 228506 408574
rect 228742 408338 228774 408574
rect 228154 390894 228774 408338
rect 228154 390658 228186 390894
rect 228422 390658 228506 390894
rect 228742 390658 228774 390894
rect 228154 390574 228774 390658
rect 228154 390338 228186 390574
rect 228422 390338 228506 390574
rect 228742 390338 228774 390574
rect 228154 372894 228774 390338
rect 228154 372658 228186 372894
rect 228422 372658 228506 372894
rect 228742 372658 228774 372894
rect 228154 372574 228774 372658
rect 228154 372338 228186 372574
rect 228422 372338 228506 372574
rect 228742 372338 228774 372574
rect 228154 354894 228774 372338
rect 228154 354658 228186 354894
rect 228422 354658 228506 354894
rect 228742 354658 228774 354894
rect 228154 354574 228774 354658
rect 228154 354338 228186 354574
rect 228422 354338 228506 354574
rect 228742 354338 228774 354574
rect 228154 336894 228774 354338
rect 228154 336658 228186 336894
rect 228422 336658 228506 336894
rect 228742 336658 228774 336894
rect 228154 336574 228774 336658
rect 228154 336338 228186 336574
rect 228422 336338 228506 336574
rect 228742 336338 228774 336574
rect 228154 318894 228774 336338
rect 228154 318658 228186 318894
rect 228422 318658 228506 318894
rect 228742 318658 228774 318894
rect 228154 318574 228774 318658
rect 228154 318338 228186 318574
rect 228422 318338 228506 318574
rect 228742 318338 228774 318574
rect 228154 300894 228774 318338
rect 228154 300658 228186 300894
rect 228422 300658 228506 300894
rect 228742 300658 228774 300894
rect 228154 300574 228774 300658
rect 228154 300338 228186 300574
rect 228422 300338 228506 300574
rect 228742 300338 228774 300574
rect 228154 282894 228774 300338
rect 228154 282658 228186 282894
rect 228422 282658 228506 282894
rect 228742 282658 228774 282894
rect 228154 282574 228774 282658
rect 228154 282338 228186 282574
rect 228422 282338 228506 282574
rect 228742 282338 228774 282574
rect 228154 264894 228774 282338
rect 228154 264658 228186 264894
rect 228422 264658 228506 264894
rect 228742 264658 228774 264894
rect 228154 264574 228774 264658
rect 228154 264338 228186 264574
rect 228422 264338 228506 264574
rect 228742 264338 228774 264574
rect 228154 246894 228774 264338
rect 228154 246658 228186 246894
rect 228422 246658 228506 246894
rect 228742 246658 228774 246894
rect 228154 246574 228774 246658
rect 228154 246338 228186 246574
rect 228422 246338 228506 246574
rect 228742 246338 228774 246574
rect 228154 228894 228774 246338
rect 228154 228658 228186 228894
rect 228422 228658 228506 228894
rect 228742 228658 228774 228894
rect 228154 228574 228774 228658
rect 228154 228338 228186 228574
rect 228422 228338 228506 228574
rect 228742 228338 228774 228574
rect 228154 210894 228774 228338
rect 228154 210658 228186 210894
rect 228422 210658 228506 210894
rect 228742 210658 228774 210894
rect 228154 210574 228774 210658
rect 228154 210338 228186 210574
rect 228422 210338 228506 210574
rect 228742 210338 228774 210574
rect 228154 192894 228774 210338
rect 228154 192658 228186 192894
rect 228422 192658 228506 192894
rect 228742 192658 228774 192894
rect 228154 192574 228774 192658
rect 228154 192338 228186 192574
rect 228422 192338 228506 192574
rect 228742 192338 228774 192574
rect 228154 174894 228774 192338
rect 228154 174658 228186 174894
rect 228422 174658 228506 174894
rect 228742 174658 228774 174894
rect 228154 174574 228774 174658
rect 228154 174338 228186 174574
rect 228422 174338 228506 174574
rect 228742 174338 228774 174574
rect 228154 156894 228774 174338
rect 228154 156658 228186 156894
rect 228422 156658 228506 156894
rect 228742 156658 228774 156894
rect 228154 156574 228774 156658
rect 228154 156338 228186 156574
rect 228422 156338 228506 156574
rect 228742 156338 228774 156574
rect 228154 138894 228774 156338
rect 228154 138658 228186 138894
rect 228422 138658 228506 138894
rect 228742 138658 228774 138894
rect 228154 138574 228774 138658
rect 228154 138338 228186 138574
rect 228422 138338 228506 138574
rect 228742 138338 228774 138574
rect 228154 120894 228774 138338
rect 228154 120658 228186 120894
rect 228422 120658 228506 120894
rect 228742 120658 228774 120894
rect 228154 120574 228774 120658
rect 228154 120338 228186 120574
rect 228422 120338 228506 120574
rect 228742 120338 228774 120574
rect 228154 102894 228774 120338
rect 228154 102658 228186 102894
rect 228422 102658 228506 102894
rect 228742 102658 228774 102894
rect 228154 102574 228774 102658
rect 228154 102338 228186 102574
rect 228422 102338 228506 102574
rect 228742 102338 228774 102574
rect 228154 84894 228774 102338
rect 228154 84658 228186 84894
rect 228422 84658 228506 84894
rect 228742 84658 228774 84894
rect 228154 84574 228774 84658
rect 228154 84338 228186 84574
rect 228422 84338 228506 84574
rect 228742 84338 228774 84574
rect 228154 66894 228774 84338
rect 228154 66658 228186 66894
rect 228422 66658 228506 66894
rect 228742 66658 228774 66894
rect 228154 66574 228774 66658
rect 228154 66338 228186 66574
rect 228422 66338 228506 66574
rect 228742 66338 228774 66574
rect 228154 48894 228774 66338
rect 228154 48658 228186 48894
rect 228422 48658 228506 48894
rect 228742 48658 228774 48894
rect 228154 48574 228774 48658
rect 228154 48338 228186 48574
rect 228422 48338 228506 48574
rect 228742 48338 228774 48574
rect 228154 30894 228774 48338
rect 228154 30658 228186 30894
rect 228422 30658 228506 30894
rect 228742 30658 228774 30894
rect 228154 30574 228774 30658
rect 228154 30338 228186 30574
rect 228422 30338 228506 30574
rect 228742 30338 228774 30574
rect 228154 12894 228774 30338
rect 228154 12658 228186 12894
rect 228422 12658 228506 12894
rect 228742 12658 228774 12894
rect 228154 12574 228774 12658
rect 228154 12338 228186 12574
rect 228422 12338 228506 12574
rect 228742 12338 228774 12574
rect 228154 -2776 228774 12338
rect 228154 -3012 228186 -2776
rect 228422 -3012 228506 -2776
rect 228742 -3012 228774 -2776
rect 228154 -3096 228774 -3012
rect 228154 -3332 228186 -3096
rect 228422 -3332 228506 -3096
rect 228742 -3332 228774 -3096
rect 228154 -4324 228774 -3332
rect 231874 463972 232494 464004
rect 231874 463736 231906 463972
rect 232142 463736 232226 463972
rect 232462 463736 232494 463972
rect 231874 463652 232494 463736
rect 231874 463416 231906 463652
rect 232142 463416 232226 463652
rect 232462 463416 232494 463652
rect 231874 448614 232494 463416
rect 231874 448378 231906 448614
rect 232142 448378 232226 448614
rect 232462 448378 232494 448614
rect 231874 448294 232494 448378
rect 231874 448058 231906 448294
rect 232142 448058 232226 448294
rect 232462 448058 232494 448294
rect 231874 430614 232494 448058
rect 231874 430378 231906 430614
rect 232142 430378 232226 430614
rect 232462 430378 232494 430614
rect 231874 430294 232494 430378
rect 231874 430058 231906 430294
rect 232142 430058 232226 430294
rect 232462 430058 232494 430294
rect 231874 412614 232494 430058
rect 231874 412378 231906 412614
rect 232142 412378 232226 412614
rect 232462 412378 232494 412614
rect 231874 412294 232494 412378
rect 231874 412058 231906 412294
rect 232142 412058 232226 412294
rect 232462 412058 232494 412294
rect 231874 394614 232494 412058
rect 231874 394378 231906 394614
rect 232142 394378 232226 394614
rect 232462 394378 232494 394614
rect 231874 394294 232494 394378
rect 231874 394058 231906 394294
rect 232142 394058 232226 394294
rect 232462 394058 232494 394294
rect 231874 376614 232494 394058
rect 231874 376378 231906 376614
rect 232142 376378 232226 376614
rect 232462 376378 232494 376614
rect 231874 376294 232494 376378
rect 231874 376058 231906 376294
rect 232142 376058 232226 376294
rect 232462 376058 232494 376294
rect 231874 358614 232494 376058
rect 231874 358378 231906 358614
rect 232142 358378 232226 358614
rect 232462 358378 232494 358614
rect 231874 358294 232494 358378
rect 231874 358058 231906 358294
rect 232142 358058 232226 358294
rect 232462 358058 232494 358294
rect 231874 340614 232494 358058
rect 231874 340378 231906 340614
rect 232142 340378 232226 340614
rect 232462 340378 232494 340614
rect 231874 340294 232494 340378
rect 231874 340058 231906 340294
rect 232142 340058 232226 340294
rect 232462 340058 232494 340294
rect 231874 322614 232494 340058
rect 231874 322378 231906 322614
rect 232142 322378 232226 322614
rect 232462 322378 232494 322614
rect 231874 322294 232494 322378
rect 231874 322058 231906 322294
rect 232142 322058 232226 322294
rect 232462 322058 232494 322294
rect 231874 304614 232494 322058
rect 231874 304378 231906 304614
rect 232142 304378 232226 304614
rect 232462 304378 232494 304614
rect 231874 304294 232494 304378
rect 231874 304058 231906 304294
rect 232142 304058 232226 304294
rect 232462 304058 232494 304294
rect 231874 286614 232494 304058
rect 231874 286378 231906 286614
rect 232142 286378 232226 286614
rect 232462 286378 232494 286614
rect 231874 286294 232494 286378
rect 231874 286058 231906 286294
rect 232142 286058 232226 286294
rect 232462 286058 232494 286294
rect 231874 268614 232494 286058
rect 231874 268378 231906 268614
rect 232142 268378 232226 268614
rect 232462 268378 232494 268614
rect 231874 268294 232494 268378
rect 231874 268058 231906 268294
rect 232142 268058 232226 268294
rect 232462 268058 232494 268294
rect 231874 250614 232494 268058
rect 231874 250378 231906 250614
rect 232142 250378 232226 250614
rect 232462 250378 232494 250614
rect 231874 250294 232494 250378
rect 231874 250058 231906 250294
rect 232142 250058 232226 250294
rect 232462 250058 232494 250294
rect 231874 232614 232494 250058
rect 231874 232378 231906 232614
rect 232142 232378 232226 232614
rect 232462 232378 232494 232614
rect 231874 232294 232494 232378
rect 231874 232058 231906 232294
rect 232142 232058 232226 232294
rect 232462 232058 232494 232294
rect 231874 214614 232494 232058
rect 231874 214378 231906 214614
rect 232142 214378 232226 214614
rect 232462 214378 232494 214614
rect 231874 214294 232494 214378
rect 231874 214058 231906 214294
rect 232142 214058 232226 214294
rect 232462 214058 232494 214294
rect 231874 196614 232494 214058
rect 231874 196378 231906 196614
rect 232142 196378 232226 196614
rect 232462 196378 232494 196614
rect 231874 196294 232494 196378
rect 231874 196058 231906 196294
rect 232142 196058 232226 196294
rect 232462 196058 232494 196294
rect 231874 178614 232494 196058
rect 231874 178378 231906 178614
rect 232142 178378 232226 178614
rect 232462 178378 232494 178614
rect 231874 178294 232494 178378
rect 231874 178058 231906 178294
rect 232142 178058 232226 178294
rect 232462 178058 232494 178294
rect 231874 160614 232494 178058
rect 231874 160378 231906 160614
rect 232142 160378 232226 160614
rect 232462 160378 232494 160614
rect 231874 160294 232494 160378
rect 231874 160058 231906 160294
rect 232142 160058 232226 160294
rect 232462 160058 232494 160294
rect 231874 142614 232494 160058
rect 231874 142378 231906 142614
rect 232142 142378 232226 142614
rect 232462 142378 232494 142614
rect 231874 142294 232494 142378
rect 231874 142058 231906 142294
rect 232142 142058 232226 142294
rect 232462 142058 232494 142294
rect 231874 124614 232494 142058
rect 231874 124378 231906 124614
rect 232142 124378 232226 124614
rect 232462 124378 232494 124614
rect 231874 124294 232494 124378
rect 231874 124058 231906 124294
rect 232142 124058 232226 124294
rect 232462 124058 232494 124294
rect 231874 106614 232494 124058
rect 231874 106378 231906 106614
rect 232142 106378 232226 106614
rect 232462 106378 232494 106614
rect 231874 106294 232494 106378
rect 231874 106058 231906 106294
rect 232142 106058 232226 106294
rect 232462 106058 232494 106294
rect 231874 88614 232494 106058
rect 231874 88378 231906 88614
rect 232142 88378 232226 88614
rect 232462 88378 232494 88614
rect 231874 88294 232494 88378
rect 231874 88058 231906 88294
rect 232142 88058 232226 88294
rect 232462 88058 232494 88294
rect 231874 70614 232494 88058
rect 231874 70378 231906 70614
rect 232142 70378 232226 70614
rect 232462 70378 232494 70614
rect 231874 70294 232494 70378
rect 231874 70058 231906 70294
rect 232142 70058 232226 70294
rect 232462 70058 232494 70294
rect 231874 52614 232494 70058
rect 231874 52378 231906 52614
rect 232142 52378 232226 52614
rect 232462 52378 232494 52614
rect 231874 52294 232494 52378
rect 231874 52058 231906 52294
rect 232142 52058 232226 52294
rect 232462 52058 232494 52294
rect 231874 34614 232494 52058
rect 231874 34378 231906 34614
rect 232142 34378 232226 34614
rect 232462 34378 232494 34614
rect 231874 34294 232494 34378
rect 231874 34058 231906 34294
rect 232142 34058 232226 34294
rect 232462 34058 232494 34294
rect 231874 16614 232494 34058
rect 231874 16378 231906 16614
rect 232142 16378 232226 16614
rect 232462 16378 232494 16614
rect 231874 16294 232494 16378
rect 231874 16058 231906 16294
rect 232142 16058 232226 16294
rect 232462 16058 232494 16294
rect 231874 -3736 232494 16058
rect 231874 -3972 231906 -3736
rect 232142 -3972 232226 -3736
rect 232462 -3972 232494 -3736
rect 231874 -4056 232494 -3972
rect 231874 -4292 231906 -4056
rect 232142 -4292 232226 -4056
rect 232462 -4292 232494 -4056
rect 231874 -4324 232494 -4292
rect 238714 461092 239334 464004
rect 238714 460856 238746 461092
rect 238982 460856 239066 461092
rect 239302 460856 239334 461092
rect 238714 460772 239334 460856
rect 238714 460536 238746 460772
rect 238982 460536 239066 460772
rect 239302 460536 239334 460772
rect 238714 455454 239334 460536
rect 238714 455218 238746 455454
rect 238982 455218 239066 455454
rect 239302 455218 239334 455454
rect 238714 455134 239334 455218
rect 238714 454898 238746 455134
rect 238982 454898 239066 455134
rect 239302 454898 239334 455134
rect 238714 437454 239334 454898
rect 238714 437218 238746 437454
rect 238982 437218 239066 437454
rect 239302 437218 239334 437454
rect 238714 437134 239334 437218
rect 238714 436898 238746 437134
rect 238982 436898 239066 437134
rect 239302 436898 239334 437134
rect 238714 419454 239334 436898
rect 238714 419218 238746 419454
rect 238982 419218 239066 419454
rect 239302 419218 239334 419454
rect 238714 419134 239334 419218
rect 238714 418898 238746 419134
rect 238982 418898 239066 419134
rect 239302 418898 239334 419134
rect 238714 401454 239334 418898
rect 238714 401218 238746 401454
rect 238982 401218 239066 401454
rect 239302 401218 239334 401454
rect 238714 401134 239334 401218
rect 238714 400898 238746 401134
rect 238982 400898 239066 401134
rect 239302 400898 239334 401134
rect 238714 383454 239334 400898
rect 238714 383218 238746 383454
rect 238982 383218 239066 383454
rect 239302 383218 239334 383454
rect 238714 383134 239334 383218
rect 238714 382898 238746 383134
rect 238982 382898 239066 383134
rect 239302 382898 239334 383134
rect 238714 365454 239334 382898
rect 238714 365218 238746 365454
rect 238982 365218 239066 365454
rect 239302 365218 239334 365454
rect 238714 365134 239334 365218
rect 238714 364898 238746 365134
rect 238982 364898 239066 365134
rect 239302 364898 239334 365134
rect 238714 347454 239334 364898
rect 238714 347218 238746 347454
rect 238982 347218 239066 347454
rect 239302 347218 239334 347454
rect 238714 347134 239334 347218
rect 238714 346898 238746 347134
rect 238982 346898 239066 347134
rect 239302 346898 239334 347134
rect 238714 329454 239334 346898
rect 238714 329218 238746 329454
rect 238982 329218 239066 329454
rect 239302 329218 239334 329454
rect 238714 329134 239334 329218
rect 238714 328898 238746 329134
rect 238982 328898 239066 329134
rect 239302 328898 239334 329134
rect 238714 311454 239334 328898
rect 238714 311218 238746 311454
rect 238982 311218 239066 311454
rect 239302 311218 239334 311454
rect 238714 311134 239334 311218
rect 238714 310898 238746 311134
rect 238982 310898 239066 311134
rect 239302 310898 239334 311134
rect 238714 293454 239334 310898
rect 238714 293218 238746 293454
rect 238982 293218 239066 293454
rect 239302 293218 239334 293454
rect 238714 293134 239334 293218
rect 238714 292898 238746 293134
rect 238982 292898 239066 293134
rect 239302 292898 239334 293134
rect 238714 275454 239334 292898
rect 238714 275218 238746 275454
rect 238982 275218 239066 275454
rect 239302 275218 239334 275454
rect 238714 275134 239334 275218
rect 238714 274898 238746 275134
rect 238982 274898 239066 275134
rect 239302 274898 239334 275134
rect 238714 257454 239334 274898
rect 238714 257218 238746 257454
rect 238982 257218 239066 257454
rect 239302 257218 239334 257454
rect 238714 257134 239334 257218
rect 238714 256898 238746 257134
rect 238982 256898 239066 257134
rect 239302 256898 239334 257134
rect 238714 239454 239334 256898
rect 238714 239218 238746 239454
rect 238982 239218 239066 239454
rect 239302 239218 239334 239454
rect 238714 239134 239334 239218
rect 238714 238898 238746 239134
rect 238982 238898 239066 239134
rect 239302 238898 239334 239134
rect 238714 221454 239334 238898
rect 238714 221218 238746 221454
rect 238982 221218 239066 221454
rect 239302 221218 239334 221454
rect 238714 221134 239334 221218
rect 238714 220898 238746 221134
rect 238982 220898 239066 221134
rect 239302 220898 239334 221134
rect 238714 203454 239334 220898
rect 238714 203218 238746 203454
rect 238982 203218 239066 203454
rect 239302 203218 239334 203454
rect 238714 203134 239334 203218
rect 238714 202898 238746 203134
rect 238982 202898 239066 203134
rect 239302 202898 239334 203134
rect 238714 185454 239334 202898
rect 238714 185218 238746 185454
rect 238982 185218 239066 185454
rect 239302 185218 239334 185454
rect 238714 185134 239334 185218
rect 238714 184898 238746 185134
rect 238982 184898 239066 185134
rect 239302 184898 239334 185134
rect 238714 167454 239334 184898
rect 238714 167218 238746 167454
rect 238982 167218 239066 167454
rect 239302 167218 239334 167454
rect 238714 167134 239334 167218
rect 238714 166898 238746 167134
rect 238982 166898 239066 167134
rect 239302 166898 239334 167134
rect 238714 149454 239334 166898
rect 238714 149218 238746 149454
rect 238982 149218 239066 149454
rect 239302 149218 239334 149454
rect 238714 149134 239334 149218
rect 238714 148898 238746 149134
rect 238982 148898 239066 149134
rect 239302 148898 239334 149134
rect 238714 131454 239334 148898
rect 238714 131218 238746 131454
rect 238982 131218 239066 131454
rect 239302 131218 239334 131454
rect 238714 131134 239334 131218
rect 238714 130898 238746 131134
rect 238982 130898 239066 131134
rect 239302 130898 239334 131134
rect 238714 113454 239334 130898
rect 238714 113218 238746 113454
rect 238982 113218 239066 113454
rect 239302 113218 239334 113454
rect 238714 113134 239334 113218
rect 238714 112898 238746 113134
rect 238982 112898 239066 113134
rect 239302 112898 239334 113134
rect 238714 95454 239334 112898
rect 238714 95218 238746 95454
rect 238982 95218 239066 95454
rect 239302 95218 239334 95454
rect 238714 95134 239334 95218
rect 238714 94898 238746 95134
rect 238982 94898 239066 95134
rect 239302 94898 239334 95134
rect 238714 77454 239334 94898
rect 238714 77218 238746 77454
rect 238982 77218 239066 77454
rect 239302 77218 239334 77454
rect 238714 77134 239334 77218
rect 238714 76898 238746 77134
rect 238982 76898 239066 77134
rect 239302 76898 239334 77134
rect 238714 59454 239334 76898
rect 238714 59218 238746 59454
rect 238982 59218 239066 59454
rect 239302 59218 239334 59454
rect 238714 59134 239334 59218
rect 238714 58898 238746 59134
rect 238982 58898 239066 59134
rect 239302 58898 239334 59134
rect 238714 41454 239334 58898
rect 238714 41218 238746 41454
rect 238982 41218 239066 41454
rect 239302 41218 239334 41454
rect 238714 41134 239334 41218
rect 238714 40898 238746 41134
rect 238982 40898 239066 41134
rect 239302 40898 239334 41134
rect 238714 23454 239334 40898
rect 238714 23218 238746 23454
rect 238982 23218 239066 23454
rect 239302 23218 239334 23454
rect 238714 23134 239334 23218
rect 238714 22898 238746 23134
rect 238982 22898 239066 23134
rect 239302 22898 239334 23134
rect 238714 5454 239334 22898
rect 238714 5218 238746 5454
rect 238982 5218 239066 5454
rect 239302 5218 239334 5454
rect 238714 5134 239334 5218
rect 238714 4898 238746 5134
rect 238982 4898 239066 5134
rect 239302 4898 239334 5134
rect 238714 -856 239334 4898
rect 238714 -1092 238746 -856
rect 238982 -1092 239066 -856
rect 239302 -1092 239334 -856
rect 238714 -1176 239334 -1092
rect 238714 -1412 238746 -1176
rect 238982 -1412 239066 -1176
rect 239302 -1412 239334 -1176
rect 238714 -4324 239334 -1412
rect 242434 462052 243054 464004
rect 242434 461816 242466 462052
rect 242702 461816 242786 462052
rect 243022 461816 243054 462052
rect 242434 461732 243054 461816
rect 242434 461496 242466 461732
rect 242702 461496 242786 461732
rect 243022 461496 243054 461732
rect 242434 441174 243054 461496
rect 242434 440938 242466 441174
rect 242702 440938 242786 441174
rect 243022 440938 243054 441174
rect 242434 440854 243054 440938
rect 242434 440618 242466 440854
rect 242702 440618 242786 440854
rect 243022 440618 243054 440854
rect 242434 423174 243054 440618
rect 242434 422938 242466 423174
rect 242702 422938 242786 423174
rect 243022 422938 243054 423174
rect 242434 422854 243054 422938
rect 242434 422618 242466 422854
rect 242702 422618 242786 422854
rect 243022 422618 243054 422854
rect 242434 405174 243054 422618
rect 242434 404938 242466 405174
rect 242702 404938 242786 405174
rect 243022 404938 243054 405174
rect 242434 404854 243054 404938
rect 242434 404618 242466 404854
rect 242702 404618 242786 404854
rect 243022 404618 243054 404854
rect 242434 387174 243054 404618
rect 242434 386938 242466 387174
rect 242702 386938 242786 387174
rect 243022 386938 243054 387174
rect 242434 386854 243054 386938
rect 242434 386618 242466 386854
rect 242702 386618 242786 386854
rect 243022 386618 243054 386854
rect 242434 369174 243054 386618
rect 242434 368938 242466 369174
rect 242702 368938 242786 369174
rect 243022 368938 243054 369174
rect 242434 368854 243054 368938
rect 242434 368618 242466 368854
rect 242702 368618 242786 368854
rect 243022 368618 243054 368854
rect 242434 351174 243054 368618
rect 242434 350938 242466 351174
rect 242702 350938 242786 351174
rect 243022 350938 243054 351174
rect 242434 350854 243054 350938
rect 242434 350618 242466 350854
rect 242702 350618 242786 350854
rect 243022 350618 243054 350854
rect 242434 333174 243054 350618
rect 242434 332938 242466 333174
rect 242702 332938 242786 333174
rect 243022 332938 243054 333174
rect 242434 332854 243054 332938
rect 242434 332618 242466 332854
rect 242702 332618 242786 332854
rect 243022 332618 243054 332854
rect 242434 315174 243054 332618
rect 242434 314938 242466 315174
rect 242702 314938 242786 315174
rect 243022 314938 243054 315174
rect 242434 314854 243054 314938
rect 242434 314618 242466 314854
rect 242702 314618 242786 314854
rect 243022 314618 243054 314854
rect 242434 297174 243054 314618
rect 242434 296938 242466 297174
rect 242702 296938 242786 297174
rect 243022 296938 243054 297174
rect 242434 296854 243054 296938
rect 242434 296618 242466 296854
rect 242702 296618 242786 296854
rect 243022 296618 243054 296854
rect 242434 279174 243054 296618
rect 242434 278938 242466 279174
rect 242702 278938 242786 279174
rect 243022 278938 243054 279174
rect 242434 278854 243054 278938
rect 242434 278618 242466 278854
rect 242702 278618 242786 278854
rect 243022 278618 243054 278854
rect 242434 261174 243054 278618
rect 242434 260938 242466 261174
rect 242702 260938 242786 261174
rect 243022 260938 243054 261174
rect 242434 260854 243054 260938
rect 242434 260618 242466 260854
rect 242702 260618 242786 260854
rect 243022 260618 243054 260854
rect 242434 243174 243054 260618
rect 242434 242938 242466 243174
rect 242702 242938 242786 243174
rect 243022 242938 243054 243174
rect 242434 242854 243054 242938
rect 242434 242618 242466 242854
rect 242702 242618 242786 242854
rect 243022 242618 243054 242854
rect 242434 225174 243054 242618
rect 242434 224938 242466 225174
rect 242702 224938 242786 225174
rect 243022 224938 243054 225174
rect 242434 224854 243054 224938
rect 242434 224618 242466 224854
rect 242702 224618 242786 224854
rect 243022 224618 243054 224854
rect 242434 207174 243054 224618
rect 242434 206938 242466 207174
rect 242702 206938 242786 207174
rect 243022 206938 243054 207174
rect 242434 206854 243054 206938
rect 242434 206618 242466 206854
rect 242702 206618 242786 206854
rect 243022 206618 243054 206854
rect 242434 189174 243054 206618
rect 242434 188938 242466 189174
rect 242702 188938 242786 189174
rect 243022 188938 243054 189174
rect 242434 188854 243054 188938
rect 242434 188618 242466 188854
rect 242702 188618 242786 188854
rect 243022 188618 243054 188854
rect 242434 171174 243054 188618
rect 242434 170938 242466 171174
rect 242702 170938 242786 171174
rect 243022 170938 243054 171174
rect 242434 170854 243054 170938
rect 242434 170618 242466 170854
rect 242702 170618 242786 170854
rect 243022 170618 243054 170854
rect 242434 153174 243054 170618
rect 242434 152938 242466 153174
rect 242702 152938 242786 153174
rect 243022 152938 243054 153174
rect 242434 152854 243054 152938
rect 242434 152618 242466 152854
rect 242702 152618 242786 152854
rect 243022 152618 243054 152854
rect 242434 135174 243054 152618
rect 242434 134938 242466 135174
rect 242702 134938 242786 135174
rect 243022 134938 243054 135174
rect 242434 134854 243054 134938
rect 242434 134618 242466 134854
rect 242702 134618 242786 134854
rect 243022 134618 243054 134854
rect 242434 117174 243054 134618
rect 242434 116938 242466 117174
rect 242702 116938 242786 117174
rect 243022 116938 243054 117174
rect 242434 116854 243054 116938
rect 242434 116618 242466 116854
rect 242702 116618 242786 116854
rect 243022 116618 243054 116854
rect 242434 99174 243054 116618
rect 242434 98938 242466 99174
rect 242702 98938 242786 99174
rect 243022 98938 243054 99174
rect 242434 98854 243054 98938
rect 242434 98618 242466 98854
rect 242702 98618 242786 98854
rect 243022 98618 243054 98854
rect 242434 81174 243054 98618
rect 242434 80938 242466 81174
rect 242702 80938 242786 81174
rect 243022 80938 243054 81174
rect 242434 80854 243054 80938
rect 242434 80618 242466 80854
rect 242702 80618 242786 80854
rect 243022 80618 243054 80854
rect 242434 63174 243054 80618
rect 242434 62938 242466 63174
rect 242702 62938 242786 63174
rect 243022 62938 243054 63174
rect 242434 62854 243054 62938
rect 242434 62618 242466 62854
rect 242702 62618 242786 62854
rect 243022 62618 243054 62854
rect 242434 45174 243054 62618
rect 242434 44938 242466 45174
rect 242702 44938 242786 45174
rect 243022 44938 243054 45174
rect 242434 44854 243054 44938
rect 242434 44618 242466 44854
rect 242702 44618 242786 44854
rect 243022 44618 243054 44854
rect 242434 27174 243054 44618
rect 242434 26938 242466 27174
rect 242702 26938 242786 27174
rect 243022 26938 243054 27174
rect 242434 26854 243054 26938
rect 242434 26618 242466 26854
rect 242702 26618 242786 26854
rect 243022 26618 243054 26854
rect 242434 9174 243054 26618
rect 242434 8938 242466 9174
rect 242702 8938 242786 9174
rect 243022 8938 243054 9174
rect 242434 8854 243054 8938
rect 242434 8618 242466 8854
rect 242702 8618 242786 8854
rect 243022 8618 243054 8854
rect 242434 -1816 243054 8618
rect 242434 -2052 242466 -1816
rect 242702 -2052 242786 -1816
rect 243022 -2052 243054 -1816
rect 242434 -2136 243054 -2052
rect 242434 -2372 242466 -2136
rect 242702 -2372 242786 -2136
rect 243022 -2372 243054 -2136
rect 242434 -4324 243054 -2372
rect 246154 463012 246774 464004
rect 246154 462776 246186 463012
rect 246422 462776 246506 463012
rect 246742 462776 246774 463012
rect 246154 462692 246774 462776
rect 246154 462456 246186 462692
rect 246422 462456 246506 462692
rect 246742 462456 246774 462692
rect 246154 444894 246774 462456
rect 246154 444658 246186 444894
rect 246422 444658 246506 444894
rect 246742 444658 246774 444894
rect 246154 444574 246774 444658
rect 246154 444338 246186 444574
rect 246422 444338 246506 444574
rect 246742 444338 246774 444574
rect 246154 426894 246774 444338
rect 246154 426658 246186 426894
rect 246422 426658 246506 426894
rect 246742 426658 246774 426894
rect 246154 426574 246774 426658
rect 246154 426338 246186 426574
rect 246422 426338 246506 426574
rect 246742 426338 246774 426574
rect 246154 408894 246774 426338
rect 246154 408658 246186 408894
rect 246422 408658 246506 408894
rect 246742 408658 246774 408894
rect 246154 408574 246774 408658
rect 246154 408338 246186 408574
rect 246422 408338 246506 408574
rect 246742 408338 246774 408574
rect 246154 390894 246774 408338
rect 246154 390658 246186 390894
rect 246422 390658 246506 390894
rect 246742 390658 246774 390894
rect 246154 390574 246774 390658
rect 246154 390338 246186 390574
rect 246422 390338 246506 390574
rect 246742 390338 246774 390574
rect 246154 372894 246774 390338
rect 246154 372658 246186 372894
rect 246422 372658 246506 372894
rect 246742 372658 246774 372894
rect 246154 372574 246774 372658
rect 246154 372338 246186 372574
rect 246422 372338 246506 372574
rect 246742 372338 246774 372574
rect 246154 354894 246774 372338
rect 246154 354658 246186 354894
rect 246422 354658 246506 354894
rect 246742 354658 246774 354894
rect 246154 354574 246774 354658
rect 246154 354338 246186 354574
rect 246422 354338 246506 354574
rect 246742 354338 246774 354574
rect 246154 336894 246774 354338
rect 246154 336658 246186 336894
rect 246422 336658 246506 336894
rect 246742 336658 246774 336894
rect 246154 336574 246774 336658
rect 246154 336338 246186 336574
rect 246422 336338 246506 336574
rect 246742 336338 246774 336574
rect 246154 318894 246774 336338
rect 246154 318658 246186 318894
rect 246422 318658 246506 318894
rect 246742 318658 246774 318894
rect 246154 318574 246774 318658
rect 246154 318338 246186 318574
rect 246422 318338 246506 318574
rect 246742 318338 246774 318574
rect 246154 300894 246774 318338
rect 246154 300658 246186 300894
rect 246422 300658 246506 300894
rect 246742 300658 246774 300894
rect 246154 300574 246774 300658
rect 246154 300338 246186 300574
rect 246422 300338 246506 300574
rect 246742 300338 246774 300574
rect 246154 282894 246774 300338
rect 246154 282658 246186 282894
rect 246422 282658 246506 282894
rect 246742 282658 246774 282894
rect 246154 282574 246774 282658
rect 246154 282338 246186 282574
rect 246422 282338 246506 282574
rect 246742 282338 246774 282574
rect 246154 264894 246774 282338
rect 246154 264658 246186 264894
rect 246422 264658 246506 264894
rect 246742 264658 246774 264894
rect 246154 264574 246774 264658
rect 246154 264338 246186 264574
rect 246422 264338 246506 264574
rect 246742 264338 246774 264574
rect 246154 246894 246774 264338
rect 246154 246658 246186 246894
rect 246422 246658 246506 246894
rect 246742 246658 246774 246894
rect 246154 246574 246774 246658
rect 246154 246338 246186 246574
rect 246422 246338 246506 246574
rect 246742 246338 246774 246574
rect 246154 228894 246774 246338
rect 246154 228658 246186 228894
rect 246422 228658 246506 228894
rect 246742 228658 246774 228894
rect 246154 228574 246774 228658
rect 246154 228338 246186 228574
rect 246422 228338 246506 228574
rect 246742 228338 246774 228574
rect 246154 210894 246774 228338
rect 246154 210658 246186 210894
rect 246422 210658 246506 210894
rect 246742 210658 246774 210894
rect 246154 210574 246774 210658
rect 246154 210338 246186 210574
rect 246422 210338 246506 210574
rect 246742 210338 246774 210574
rect 246154 192894 246774 210338
rect 246154 192658 246186 192894
rect 246422 192658 246506 192894
rect 246742 192658 246774 192894
rect 246154 192574 246774 192658
rect 246154 192338 246186 192574
rect 246422 192338 246506 192574
rect 246742 192338 246774 192574
rect 246154 174894 246774 192338
rect 246154 174658 246186 174894
rect 246422 174658 246506 174894
rect 246742 174658 246774 174894
rect 246154 174574 246774 174658
rect 246154 174338 246186 174574
rect 246422 174338 246506 174574
rect 246742 174338 246774 174574
rect 246154 156894 246774 174338
rect 246154 156658 246186 156894
rect 246422 156658 246506 156894
rect 246742 156658 246774 156894
rect 246154 156574 246774 156658
rect 246154 156338 246186 156574
rect 246422 156338 246506 156574
rect 246742 156338 246774 156574
rect 246154 138894 246774 156338
rect 246154 138658 246186 138894
rect 246422 138658 246506 138894
rect 246742 138658 246774 138894
rect 246154 138574 246774 138658
rect 246154 138338 246186 138574
rect 246422 138338 246506 138574
rect 246742 138338 246774 138574
rect 246154 120894 246774 138338
rect 246154 120658 246186 120894
rect 246422 120658 246506 120894
rect 246742 120658 246774 120894
rect 246154 120574 246774 120658
rect 246154 120338 246186 120574
rect 246422 120338 246506 120574
rect 246742 120338 246774 120574
rect 246154 102894 246774 120338
rect 246154 102658 246186 102894
rect 246422 102658 246506 102894
rect 246742 102658 246774 102894
rect 246154 102574 246774 102658
rect 246154 102338 246186 102574
rect 246422 102338 246506 102574
rect 246742 102338 246774 102574
rect 246154 84894 246774 102338
rect 246154 84658 246186 84894
rect 246422 84658 246506 84894
rect 246742 84658 246774 84894
rect 246154 84574 246774 84658
rect 246154 84338 246186 84574
rect 246422 84338 246506 84574
rect 246742 84338 246774 84574
rect 246154 66894 246774 84338
rect 246154 66658 246186 66894
rect 246422 66658 246506 66894
rect 246742 66658 246774 66894
rect 246154 66574 246774 66658
rect 246154 66338 246186 66574
rect 246422 66338 246506 66574
rect 246742 66338 246774 66574
rect 246154 48894 246774 66338
rect 246154 48658 246186 48894
rect 246422 48658 246506 48894
rect 246742 48658 246774 48894
rect 246154 48574 246774 48658
rect 246154 48338 246186 48574
rect 246422 48338 246506 48574
rect 246742 48338 246774 48574
rect 246154 30894 246774 48338
rect 246154 30658 246186 30894
rect 246422 30658 246506 30894
rect 246742 30658 246774 30894
rect 246154 30574 246774 30658
rect 246154 30338 246186 30574
rect 246422 30338 246506 30574
rect 246742 30338 246774 30574
rect 246154 12894 246774 30338
rect 246154 12658 246186 12894
rect 246422 12658 246506 12894
rect 246742 12658 246774 12894
rect 246154 12574 246774 12658
rect 246154 12338 246186 12574
rect 246422 12338 246506 12574
rect 246742 12338 246774 12574
rect 246154 -2776 246774 12338
rect 246154 -3012 246186 -2776
rect 246422 -3012 246506 -2776
rect 246742 -3012 246774 -2776
rect 246154 -3096 246774 -3012
rect 246154 -3332 246186 -3096
rect 246422 -3332 246506 -3096
rect 246742 -3332 246774 -3096
rect 246154 -4324 246774 -3332
rect 249874 463972 250494 464004
rect 249874 463736 249906 463972
rect 250142 463736 250226 463972
rect 250462 463736 250494 463972
rect 249874 463652 250494 463736
rect 249874 463416 249906 463652
rect 250142 463416 250226 463652
rect 250462 463416 250494 463652
rect 249874 448614 250494 463416
rect 249874 448378 249906 448614
rect 250142 448378 250226 448614
rect 250462 448378 250494 448614
rect 249874 448294 250494 448378
rect 249874 448058 249906 448294
rect 250142 448058 250226 448294
rect 250462 448058 250494 448294
rect 249874 430614 250494 448058
rect 249874 430378 249906 430614
rect 250142 430378 250226 430614
rect 250462 430378 250494 430614
rect 249874 430294 250494 430378
rect 249874 430058 249906 430294
rect 250142 430058 250226 430294
rect 250462 430058 250494 430294
rect 249874 412614 250494 430058
rect 249874 412378 249906 412614
rect 250142 412378 250226 412614
rect 250462 412378 250494 412614
rect 249874 412294 250494 412378
rect 249874 412058 249906 412294
rect 250142 412058 250226 412294
rect 250462 412058 250494 412294
rect 249874 394614 250494 412058
rect 249874 394378 249906 394614
rect 250142 394378 250226 394614
rect 250462 394378 250494 394614
rect 249874 394294 250494 394378
rect 249874 394058 249906 394294
rect 250142 394058 250226 394294
rect 250462 394058 250494 394294
rect 249874 376614 250494 394058
rect 249874 376378 249906 376614
rect 250142 376378 250226 376614
rect 250462 376378 250494 376614
rect 249874 376294 250494 376378
rect 249874 376058 249906 376294
rect 250142 376058 250226 376294
rect 250462 376058 250494 376294
rect 249874 358614 250494 376058
rect 249874 358378 249906 358614
rect 250142 358378 250226 358614
rect 250462 358378 250494 358614
rect 249874 358294 250494 358378
rect 249874 358058 249906 358294
rect 250142 358058 250226 358294
rect 250462 358058 250494 358294
rect 249874 340614 250494 358058
rect 249874 340378 249906 340614
rect 250142 340378 250226 340614
rect 250462 340378 250494 340614
rect 249874 340294 250494 340378
rect 249874 340058 249906 340294
rect 250142 340058 250226 340294
rect 250462 340058 250494 340294
rect 249874 322614 250494 340058
rect 249874 322378 249906 322614
rect 250142 322378 250226 322614
rect 250462 322378 250494 322614
rect 249874 322294 250494 322378
rect 249874 322058 249906 322294
rect 250142 322058 250226 322294
rect 250462 322058 250494 322294
rect 249874 304614 250494 322058
rect 249874 304378 249906 304614
rect 250142 304378 250226 304614
rect 250462 304378 250494 304614
rect 249874 304294 250494 304378
rect 249874 304058 249906 304294
rect 250142 304058 250226 304294
rect 250462 304058 250494 304294
rect 249874 286614 250494 304058
rect 249874 286378 249906 286614
rect 250142 286378 250226 286614
rect 250462 286378 250494 286614
rect 249874 286294 250494 286378
rect 249874 286058 249906 286294
rect 250142 286058 250226 286294
rect 250462 286058 250494 286294
rect 249874 268614 250494 286058
rect 249874 268378 249906 268614
rect 250142 268378 250226 268614
rect 250462 268378 250494 268614
rect 249874 268294 250494 268378
rect 249874 268058 249906 268294
rect 250142 268058 250226 268294
rect 250462 268058 250494 268294
rect 249874 250614 250494 268058
rect 249874 250378 249906 250614
rect 250142 250378 250226 250614
rect 250462 250378 250494 250614
rect 249874 250294 250494 250378
rect 249874 250058 249906 250294
rect 250142 250058 250226 250294
rect 250462 250058 250494 250294
rect 249874 232614 250494 250058
rect 249874 232378 249906 232614
rect 250142 232378 250226 232614
rect 250462 232378 250494 232614
rect 249874 232294 250494 232378
rect 249874 232058 249906 232294
rect 250142 232058 250226 232294
rect 250462 232058 250494 232294
rect 249874 214614 250494 232058
rect 249874 214378 249906 214614
rect 250142 214378 250226 214614
rect 250462 214378 250494 214614
rect 249874 214294 250494 214378
rect 249874 214058 249906 214294
rect 250142 214058 250226 214294
rect 250462 214058 250494 214294
rect 249874 196614 250494 214058
rect 249874 196378 249906 196614
rect 250142 196378 250226 196614
rect 250462 196378 250494 196614
rect 249874 196294 250494 196378
rect 249874 196058 249906 196294
rect 250142 196058 250226 196294
rect 250462 196058 250494 196294
rect 249874 178614 250494 196058
rect 249874 178378 249906 178614
rect 250142 178378 250226 178614
rect 250462 178378 250494 178614
rect 249874 178294 250494 178378
rect 249874 178058 249906 178294
rect 250142 178058 250226 178294
rect 250462 178058 250494 178294
rect 249874 160614 250494 178058
rect 249874 160378 249906 160614
rect 250142 160378 250226 160614
rect 250462 160378 250494 160614
rect 249874 160294 250494 160378
rect 249874 160058 249906 160294
rect 250142 160058 250226 160294
rect 250462 160058 250494 160294
rect 249874 142614 250494 160058
rect 249874 142378 249906 142614
rect 250142 142378 250226 142614
rect 250462 142378 250494 142614
rect 249874 142294 250494 142378
rect 249874 142058 249906 142294
rect 250142 142058 250226 142294
rect 250462 142058 250494 142294
rect 249874 124614 250494 142058
rect 249874 124378 249906 124614
rect 250142 124378 250226 124614
rect 250462 124378 250494 124614
rect 249874 124294 250494 124378
rect 249874 124058 249906 124294
rect 250142 124058 250226 124294
rect 250462 124058 250494 124294
rect 249874 106614 250494 124058
rect 249874 106378 249906 106614
rect 250142 106378 250226 106614
rect 250462 106378 250494 106614
rect 249874 106294 250494 106378
rect 249874 106058 249906 106294
rect 250142 106058 250226 106294
rect 250462 106058 250494 106294
rect 249874 88614 250494 106058
rect 249874 88378 249906 88614
rect 250142 88378 250226 88614
rect 250462 88378 250494 88614
rect 249874 88294 250494 88378
rect 249874 88058 249906 88294
rect 250142 88058 250226 88294
rect 250462 88058 250494 88294
rect 249874 70614 250494 88058
rect 249874 70378 249906 70614
rect 250142 70378 250226 70614
rect 250462 70378 250494 70614
rect 249874 70294 250494 70378
rect 249874 70058 249906 70294
rect 250142 70058 250226 70294
rect 250462 70058 250494 70294
rect 249874 52614 250494 70058
rect 249874 52378 249906 52614
rect 250142 52378 250226 52614
rect 250462 52378 250494 52614
rect 249874 52294 250494 52378
rect 249874 52058 249906 52294
rect 250142 52058 250226 52294
rect 250462 52058 250494 52294
rect 249874 34614 250494 52058
rect 249874 34378 249906 34614
rect 250142 34378 250226 34614
rect 250462 34378 250494 34614
rect 249874 34294 250494 34378
rect 249874 34058 249906 34294
rect 250142 34058 250226 34294
rect 250462 34058 250494 34294
rect 249874 16614 250494 34058
rect 249874 16378 249906 16614
rect 250142 16378 250226 16614
rect 250462 16378 250494 16614
rect 249874 16294 250494 16378
rect 249874 16058 249906 16294
rect 250142 16058 250226 16294
rect 250462 16058 250494 16294
rect 249874 -3736 250494 16058
rect 249874 -3972 249906 -3736
rect 250142 -3972 250226 -3736
rect 250462 -3972 250494 -3736
rect 249874 -4056 250494 -3972
rect 249874 -4292 249906 -4056
rect 250142 -4292 250226 -4056
rect 250462 -4292 250494 -4056
rect 249874 -4324 250494 -4292
rect 256714 461092 257334 464004
rect 256714 460856 256746 461092
rect 256982 460856 257066 461092
rect 257302 460856 257334 461092
rect 256714 460772 257334 460856
rect 256714 460536 256746 460772
rect 256982 460536 257066 460772
rect 257302 460536 257334 460772
rect 256714 455454 257334 460536
rect 256714 455218 256746 455454
rect 256982 455218 257066 455454
rect 257302 455218 257334 455454
rect 256714 455134 257334 455218
rect 256714 454898 256746 455134
rect 256982 454898 257066 455134
rect 257302 454898 257334 455134
rect 256714 437454 257334 454898
rect 256714 437218 256746 437454
rect 256982 437218 257066 437454
rect 257302 437218 257334 437454
rect 256714 437134 257334 437218
rect 256714 436898 256746 437134
rect 256982 436898 257066 437134
rect 257302 436898 257334 437134
rect 256714 419454 257334 436898
rect 256714 419218 256746 419454
rect 256982 419218 257066 419454
rect 257302 419218 257334 419454
rect 256714 419134 257334 419218
rect 256714 418898 256746 419134
rect 256982 418898 257066 419134
rect 257302 418898 257334 419134
rect 256714 401454 257334 418898
rect 256714 401218 256746 401454
rect 256982 401218 257066 401454
rect 257302 401218 257334 401454
rect 256714 401134 257334 401218
rect 256714 400898 256746 401134
rect 256982 400898 257066 401134
rect 257302 400898 257334 401134
rect 256714 383454 257334 400898
rect 256714 383218 256746 383454
rect 256982 383218 257066 383454
rect 257302 383218 257334 383454
rect 256714 383134 257334 383218
rect 256714 382898 256746 383134
rect 256982 382898 257066 383134
rect 257302 382898 257334 383134
rect 256714 365454 257334 382898
rect 256714 365218 256746 365454
rect 256982 365218 257066 365454
rect 257302 365218 257334 365454
rect 256714 365134 257334 365218
rect 256714 364898 256746 365134
rect 256982 364898 257066 365134
rect 257302 364898 257334 365134
rect 256714 347454 257334 364898
rect 256714 347218 256746 347454
rect 256982 347218 257066 347454
rect 257302 347218 257334 347454
rect 256714 347134 257334 347218
rect 256714 346898 256746 347134
rect 256982 346898 257066 347134
rect 257302 346898 257334 347134
rect 256714 329454 257334 346898
rect 256714 329218 256746 329454
rect 256982 329218 257066 329454
rect 257302 329218 257334 329454
rect 256714 329134 257334 329218
rect 256714 328898 256746 329134
rect 256982 328898 257066 329134
rect 257302 328898 257334 329134
rect 256714 311454 257334 328898
rect 256714 311218 256746 311454
rect 256982 311218 257066 311454
rect 257302 311218 257334 311454
rect 256714 311134 257334 311218
rect 256714 310898 256746 311134
rect 256982 310898 257066 311134
rect 257302 310898 257334 311134
rect 256714 293454 257334 310898
rect 256714 293218 256746 293454
rect 256982 293218 257066 293454
rect 257302 293218 257334 293454
rect 256714 293134 257334 293218
rect 256714 292898 256746 293134
rect 256982 292898 257066 293134
rect 257302 292898 257334 293134
rect 256714 275454 257334 292898
rect 256714 275218 256746 275454
rect 256982 275218 257066 275454
rect 257302 275218 257334 275454
rect 256714 275134 257334 275218
rect 256714 274898 256746 275134
rect 256982 274898 257066 275134
rect 257302 274898 257334 275134
rect 256714 257454 257334 274898
rect 256714 257218 256746 257454
rect 256982 257218 257066 257454
rect 257302 257218 257334 257454
rect 256714 257134 257334 257218
rect 256714 256898 256746 257134
rect 256982 256898 257066 257134
rect 257302 256898 257334 257134
rect 256714 239454 257334 256898
rect 256714 239218 256746 239454
rect 256982 239218 257066 239454
rect 257302 239218 257334 239454
rect 256714 239134 257334 239218
rect 256714 238898 256746 239134
rect 256982 238898 257066 239134
rect 257302 238898 257334 239134
rect 256714 221454 257334 238898
rect 256714 221218 256746 221454
rect 256982 221218 257066 221454
rect 257302 221218 257334 221454
rect 256714 221134 257334 221218
rect 256714 220898 256746 221134
rect 256982 220898 257066 221134
rect 257302 220898 257334 221134
rect 256714 203454 257334 220898
rect 256714 203218 256746 203454
rect 256982 203218 257066 203454
rect 257302 203218 257334 203454
rect 256714 203134 257334 203218
rect 256714 202898 256746 203134
rect 256982 202898 257066 203134
rect 257302 202898 257334 203134
rect 256714 185454 257334 202898
rect 256714 185218 256746 185454
rect 256982 185218 257066 185454
rect 257302 185218 257334 185454
rect 256714 185134 257334 185218
rect 256714 184898 256746 185134
rect 256982 184898 257066 185134
rect 257302 184898 257334 185134
rect 256714 167454 257334 184898
rect 256714 167218 256746 167454
rect 256982 167218 257066 167454
rect 257302 167218 257334 167454
rect 256714 167134 257334 167218
rect 256714 166898 256746 167134
rect 256982 166898 257066 167134
rect 257302 166898 257334 167134
rect 256714 149454 257334 166898
rect 256714 149218 256746 149454
rect 256982 149218 257066 149454
rect 257302 149218 257334 149454
rect 256714 149134 257334 149218
rect 256714 148898 256746 149134
rect 256982 148898 257066 149134
rect 257302 148898 257334 149134
rect 256714 131454 257334 148898
rect 256714 131218 256746 131454
rect 256982 131218 257066 131454
rect 257302 131218 257334 131454
rect 256714 131134 257334 131218
rect 256714 130898 256746 131134
rect 256982 130898 257066 131134
rect 257302 130898 257334 131134
rect 256714 113454 257334 130898
rect 256714 113218 256746 113454
rect 256982 113218 257066 113454
rect 257302 113218 257334 113454
rect 256714 113134 257334 113218
rect 256714 112898 256746 113134
rect 256982 112898 257066 113134
rect 257302 112898 257334 113134
rect 256714 95454 257334 112898
rect 256714 95218 256746 95454
rect 256982 95218 257066 95454
rect 257302 95218 257334 95454
rect 256714 95134 257334 95218
rect 256714 94898 256746 95134
rect 256982 94898 257066 95134
rect 257302 94898 257334 95134
rect 256714 77454 257334 94898
rect 256714 77218 256746 77454
rect 256982 77218 257066 77454
rect 257302 77218 257334 77454
rect 256714 77134 257334 77218
rect 256714 76898 256746 77134
rect 256982 76898 257066 77134
rect 257302 76898 257334 77134
rect 256714 59454 257334 76898
rect 256714 59218 256746 59454
rect 256982 59218 257066 59454
rect 257302 59218 257334 59454
rect 256714 59134 257334 59218
rect 256714 58898 256746 59134
rect 256982 58898 257066 59134
rect 257302 58898 257334 59134
rect 256714 41454 257334 58898
rect 256714 41218 256746 41454
rect 256982 41218 257066 41454
rect 257302 41218 257334 41454
rect 256714 41134 257334 41218
rect 256714 40898 256746 41134
rect 256982 40898 257066 41134
rect 257302 40898 257334 41134
rect 256714 23454 257334 40898
rect 256714 23218 256746 23454
rect 256982 23218 257066 23454
rect 257302 23218 257334 23454
rect 256714 23134 257334 23218
rect 256714 22898 256746 23134
rect 256982 22898 257066 23134
rect 257302 22898 257334 23134
rect 256714 5454 257334 22898
rect 256714 5218 256746 5454
rect 256982 5218 257066 5454
rect 257302 5218 257334 5454
rect 256714 5134 257334 5218
rect 256714 4898 256746 5134
rect 256982 4898 257066 5134
rect 257302 4898 257334 5134
rect 256714 -856 257334 4898
rect 256714 -1092 256746 -856
rect 256982 -1092 257066 -856
rect 257302 -1092 257334 -856
rect 256714 -1176 257334 -1092
rect 256714 -1412 256746 -1176
rect 256982 -1412 257066 -1176
rect 257302 -1412 257334 -1176
rect 256714 -4324 257334 -1412
rect 260434 462052 261054 464004
rect 260434 461816 260466 462052
rect 260702 461816 260786 462052
rect 261022 461816 261054 462052
rect 260434 461732 261054 461816
rect 260434 461496 260466 461732
rect 260702 461496 260786 461732
rect 261022 461496 261054 461732
rect 260434 441174 261054 461496
rect 260434 440938 260466 441174
rect 260702 440938 260786 441174
rect 261022 440938 261054 441174
rect 260434 440854 261054 440938
rect 260434 440618 260466 440854
rect 260702 440618 260786 440854
rect 261022 440618 261054 440854
rect 260434 423174 261054 440618
rect 260434 422938 260466 423174
rect 260702 422938 260786 423174
rect 261022 422938 261054 423174
rect 260434 422854 261054 422938
rect 260434 422618 260466 422854
rect 260702 422618 260786 422854
rect 261022 422618 261054 422854
rect 260434 405174 261054 422618
rect 260434 404938 260466 405174
rect 260702 404938 260786 405174
rect 261022 404938 261054 405174
rect 260434 404854 261054 404938
rect 260434 404618 260466 404854
rect 260702 404618 260786 404854
rect 261022 404618 261054 404854
rect 260434 387174 261054 404618
rect 260434 386938 260466 387174
rect 260702 386938 260786 387174
rect 261022 386938 261054 387174
rect 260434 386854 261054 386938
rect 260434 386618 260466 386854
rect 260702 386618 260786 386854
rect 261022 386618 261054 386854
rect 260434 369174 261054 386618
rect 260434 368938 260466 369174
rect 260702 368938 260786 369174
rect 261022 368938 261054 369174
rect 260434 368854 261054 368938
rect 260434 368618 260466 368854
rect 260702 368618 260786 368854
rect 261022 368618 261054 368854
rect 260434 351174 261054 368618
rect 260434 350938 260466 351174
rect 260702 350938 260786 351174
rect 261022 350938 261054 351174
rect 260434 350854 261054 350938
rect 260434 350618 260466 350854
rect 260702 350618 260786 350854
rect 261022 350618 261054 350854
rect 260434 333174 261054 350618
rect 260434 332938 260466 333174
rect 260702 332938 260786 333174
rect 261022 332938 261054 333174
rect 260434 332854 261054 332938
rect 260434 332618 260466 332854
rect 260702 332618 260786 332854
rect 261022 332618 261054 332854
rect 260434 315174 261054 332618
rect 260434 314938 260466 315174
rect 260702 314938 260786 315174
rect 261022 314938 261054 315174
rect 260434 314854 261054 314938
rect 260434 314618 260466 314854
rect 260702 314618 260786 314854
rect 261022 314618 261054 314854
rect 260434 297174 261054 314618
rect 260434 296938 260466 297174
rect 260702 296938 260786 297174
rect 261022 296938 261054 297174
rect 260434 296854 261054 296938
rect 260434 296618 260466 296854
rect 260702 296618 260786 296854
rect 261022 296618 261054 296854
rect 260434 279174 261054 296618
rect 260434 278938 260466 279174
rect 260702 278938 260786 279174
rect 261022 278938 261054 279174
rect 260434 278854 261054 278938
rect 260434 278618 260466 278854
rect 260702 278618 260786 278854
rect 261022 278618 261054 278854
rect 260434 261174 261054 278618
rect 260434 260938 260466 261174
rect 260702 260938 260786 261174
rect 261022 260938 261054 261174
rect 260434 260854 261054 260938
rect 260434 260618 260466 260854
rect 260702 260618 260786 260854
rect 261022 260618 261054 260854
rect 260434 243174 261054 260618
rect 260434 242938 260466 243174
rect 260702 242938 260786 243174
rect 261022 242938 261054 243174
rect 260434 242854 261054 242938
rect 260434 242618 260466 242854
rect 260702 242618 260786 242854
rect 261022 242618 261054 242854
rect 260434 225174 261054 242618
rect 260434 224938 260466 225174
rect 260702 224938 260786 225174
rect 261022 224938 261054 225174
rect 260434 224854 261054 224938
rect 260434 224618 260466 224854
rect 260702 224618 260786 224854
rect 261022 224618 261054 224854
rect 260434 207174 261054 224618
rect 260434 206938 260466 207174
rect 260702 206938 260786 207174
rect 261022 206938 261054 207174
rect 260434 206854 261054 206938
rect 260434 206618 260466 206854
rect 260702 206618 260786 206854
rect 261022 206618 261054 206854
rect 260434 189174 261054 206618
rect 260434 188938 260466 189174
rect 260702 188938 260786 189174
rect 261022 188938 261054 189174
rect 260434 188854 261054 188938
rect 260434 188618 260466 188854
rect 260702 188618 260786 188854
rect 261022 188618 261054 188854
rect 260434 171174 261054 188618
rect 260434 170938 260466 171174
rect 260702 170938 260786 171174
rect 261022 170938 261054 171174
rect 260434 170854 261054 170938
rect 260434 170618 260466 170854
rect 260702 170618 260786 170854
rect 261022 170618 261054 170854
rect 260434 153174 261054 170618
rect 260434 152938 260466 153174
rect 260702 152938 260786 153174
rect 261022 152938 261054 153174
rect 260434 152854 261054 152938
rect 260434 152618 260466 152854
rect 260702 152618 260786 152854
rect 261022 152618 261054 152854
rect 260434 135174 261054 152618
rect 260434 134938 260466 135174
rect 260702 134938 260786 135174
rect 261022 134938 261054 135174
rect 260434 134854 261054 134938
rect 260434 134618 260466 134854
rect 260702 134618 260786 134854
rect 261022 134618 261054 134854
rect 260434 117174 261054 134618
rect 260434 116938 260466 117174
rect 260702 116938 260786 117174
rect 261022 116938 261054 117174
rect 260434 116854 261054 116938
rect 260434 116618 260466 116854
rect 260702 116618 260786 116854
rect 261022 116618 261054 116854
rect 260434 99174 261054 116618
rect 260434 98938 260466 99174
rect 260702 98938 260786 99174
rect 261022 98938 261054 99174
rect 260434 98854 261054 98938
rect 260434 98618 260466 98854
rect 260702 98618 260786 98854
rect 261022 98618 261054 98854
rect 260434 81174 261054 98618
rect 260434 80938 260466 81174
rect 260702 80938 260786 81174
rect 261022 80938 261054 81174
rect 260434 80854 261054 80938
rect 260434 80618 260466 80854
rect 260702 80618 260786 80854
rect 261022 80618 261054 80854
rect 260434 63174 261054 80618
rect 260434 62938 260466 63174
rect 260702 62938 260786 63174
rect 261022 62938 261054 63174
rect 260434 62854 261054 62938
rect 260434 62618 260466 62854
rect 260702 62618 260786 62854
rect 261022 62618 261054 62854
rect 260434 45174 261054 62618
rect 260434 44938 260466 45174
rect 260702 44938 260786 45174
rect 261022 44938 261054 45174
rect 260434 44854 261054 44938
rect 260434 44618 260466 44854
rect 260702 44618 260786 44854
rect 261022 44618 261054 44854
rect 260434 27174 261054 44618
rect 260434 26938 260466 27174
rect 260702 26938 260786 27174
rect 261022 26938 261054 27174
rect 260434 26854 261054 26938
rect 260434 26618 260466 26854
rect 260702 26618 260786 26854
rect 261022 26618 261054 26854
rect 260434 9174 261054 26618
rect 260434 8938 260466 9174
rect 260702 8938 260786 9174
rect 261022 8938 261054 9174
rect 260434 8854 261054 8938
rect 260434 8618 260466 8854
rect 260702 8618 260786 8854
rect 261022 8618 261054 8854
rect 260434 -1816 261054 8618
rect 260434 -2052 260466 -1816
rect 260702 -2052 260786 -1816
rect 261022 -2052 261054 -1816
rect 260434 -2136 261054 -2052
rect 260434 -2372 260466 -2136
rect 260702 -2372 260786 -2136
rect 261022 -2372 261054 -2136
rect 260434 -4324 261054 -2372
rect 264154 463012 264774 464004
rect 264154 462776 264186 463012
rect 264422 462776 264506 463012
rect 264742 462776 264774 463012
rect 264154 462692 264774 462776
rect 264154 462456 264186 462692
rect 264422 462456 264506 462692
rect 264742 462456 264774 462692
rect 264154 444894 264774 462456
rect 264154 444658 264186 444894
rect 264422 444658 264506 444894
rect 264742 444658 264774 444894
rect 264154 444574 264774 444658
rect 264154 444338 264186 444574
rect 264422 444338 264506 444574
rect 264742 444338 264774 444574
rect 264154 426894 264774 444338
rect 264154 426658 264186 426894
rect 264422 426658 264506 426894
rect 264742 426658 264774 426894
rect 264154 426574 264774 426658
rect 264154 426338 264186 426574
rect 264422 426338 264506 426574
rect 264742 426338 264774 426574
rect 264154 408894 264774 426338
rect 264154 408658 264186 408894
rect 264422 408658 264506 408894
rect 264742 408658 264774 408894
rect 264154 408574 264774 408658
rect 264154 408338 264186 408574
rect 264422 408338 264506 408574
rect 264742 408338 264774 408574
rect 264154 390894 264774 408338
rect 264154 390658 264186 390894
rect 264422 390658 264506 390894
rect 264742 390658 264774 390894
rect 264154 390574 264774 390658
rect 264154 390338 264186 390574
rect 264422 390338 264506 390574
rect 264742 390338 264774 390574
rect 264154 372894 264774 390338
rect 264154 372658 264186 372894
rect 264422 372658 264506 372894
rect 264742 372658 264774 372894
rect 264154 372574 264774 372658
rect 264154 372338 264186 372574
rect 264422 372338 264506 372574
rect 264742 372338 264774 372574
rect 264154 354894 264774 372338
rect 264154 354658 264186 354894
rect 264422 354658 264506 354894
rect 264742 354658 264774 354894
rect 264154 354574 264774 354658
rect 264154 354338 264186 354574
rect 264422 354338 264506 354574
rect 264742 354338 264774 354574
rect 264154 336894 264774 354338
rect 264154 336658 264186 336894
rect 264422 336658 264506 336894
rect 264742 336658 264774 336894
rect 264154 336574 264774 336658
rect 264154 336338 264186 336574
rect 264422 336338 264506 336574
rect 264742 336338 264774 336574
rect 264154 318894 264774 336338
rect 264154 318658 264186 318894
rect 264422 318658 264506 318894
rect 264742 318658 264774 318894
rect 264154 318574 264774 318658
rect 264154 318338 264186 318574
rect 264422 318338 264506 318574
rect 264742 318338 264774 318574
rect 264154 300894 264774 318338
rect 264154 300658 264186 300894
rect 264422 300658 264506 300894
rect 264742 300658 264774 300894
rect 264154 300574 264774 300658
rect 264154 300338 264186 300574
rect 264422 300338 264506 300574
rect 264742 300338 264774 300574
rect 264154 282894 264774 300338
rect 264154 282658 264186 282894
rect 264422 282658 264506 282894
rect 264742 282658 264774 282894
rect 264154 282574 264774 282658
rect 264154 282338 264186 282574
rect 264422 282338 264506 282574
rect 264742 282338 264774 282574
rect 264154 264894 264774 282338
rect 264154 264658 264186 264894
rect 264422 264658 264506 264894
rect 264742 264658 264774 264894
rect 264154 264574 264774 264658
rect 264154 264338 264186 264574
rect 264422 264338 264506 264574
rect 264742 264338 264774 264574
rect 264154 246894 264774 264338
rect 264154 246658 264186 246894
rect 264422 246658 264506 246894
rect 264742 246658 264774 246894
rect 264154 246574 264774 246658
rect 264154 246338 264186 246574
rect 264422 246338 264506 246574
rect 264742 246338 264774 246574
rect 264154 228894 264774 246338
rect 264154 228658 264186 228894
rect 264422 228658 264506 228894
rect 264742 228658 264774 228894
rect 264154 228574 264774 228658
rect 264154 228338 264186 228574
rect 264422 228338 264506 228574
rect 264742 228338 264774 228574
rect 264154 210894 264774 228338
rect 264154 210658 264186 210894
rect 264422 210658 264506 210894
rect 264742 210658 264774 210894
rect 264154 210574 264774 210658
rect 264154 210338 264186 210574
rect 264422 210338 264506 210574
rect 264742 210338 264774 210574
rect 264154 192894 264774 210338
rect 264154 192658 264186 192894
rect 264422 192658 264506 192894
rect 264742 192658 264774 192894
rect 264154 192574 264774 192658
rect 264154 192338 264186 192574
rect 264422 192338 264506 192574
rect 264742 192338 264774 192574
rect 264154 174894 264774 192338
rect 264154 174658 264186 174894
rect 264422 174658 264506 174894
rect 264742 174658 264774 174894
rect 264154 174574 264774 174658
rect 264154 174338 264186 174574
rect 264422 174338 264506 174574
rect 264742 174338 264774 174574
rect 264154 156894 264774 174338
rect 264154 156658 264186 156894
rect 264422 156658 264506 156894
rect 264742 156658 264774 156894
rect 264154 156574 264774 156658
rect 264154 156338 264186 156574
rect 264422 156338 264506 156574
rect 264742 156338 264774 156574
rect 264154 138894 264774 156338
rect 264154 138658 264186 138894
rect 264422 138658 264506 138894
rect 264742 138658 264774 138894
rect 264154 138574 264774 138658
rect 264154 138338 264186 138574
rect 264422 138338 264506 138574
rect 264742 138338 264774 138574
rect 264154 120894 264774 138338
rect 264154 120658 264186 120894
rect 264422 120658 264506 120894
rect 264742 120658 264774 120894
rect 264154 120574 264774 120658
rect 264154 120338 264186 120574
rect 264422 120338 264506 120574
rect 264742 120338 264774 120574
rect 264154 102894 264774 120338
rect 264154 102658 264186 102894
rect 264422 102658 264506 102894
rect 264742 102658 264774 102894
rect 264154 102574 264774 102658
rect 264154 102338 264186 102574
rect 264422 102338 264506 102574
rect 264742 102338 264774 102574
rect 264154 84894 264774 102338
rect 264154 84658 264186 84894
rect 264422 84658 264506 84894
rect 264742 84658 264774 84894
rect 264154 84574 264774 84658
rect 264154 84338 264186 84574
rect 264422 84338 264506 84574
rect 264742 84338 264774 84574
rect 264154 66894 264774 84338
rect 264154 66658 264186 66894
rect 264422 66658 264506 66894
rect 264742 66658 264774 66894
rect 264154 66574 264774 66658
rect 264154 66338 264186 66574
rect 264422 66338 264506 66574
rect 264742 66338 264774 66574
rect 264154 48894 264774 66338
rect 264154 48658 264186 48894
rect 264422 48658 264506 48894
rect 264742 48658 264774 48894
rect 264154 48574 264774 48658
rect 264154 48338 264186 48574
rect 264422 48338 264506 48574
rect 264742 48338 264774 48574
rect 264154 30894 264774 48338
rect 264154 30658 264186 30894
rect 264422 30658 264506 30894
rect 264742 30658 264774 30894
rect 264154 30574 264774 30658
rect 264154 30338 264186 30574
rect 264422 30338 264506 30574
rect 264742 30338 264774 30574
rect 264154 12894 264774 30338
rect 264154 12658 264186 12894
rect 264422 12658 264506 12894
rect 264742 12658 264774 12894
rect 264154 12574 264774 12658
rect 264154 12338 264186 12574
rect 264422 12338 264506 12574
rect 264742 12338 264774 12574
rect 264154 -2776 264774 12338
rect 264154 -3012 264186 -2776
rect 264422 -3012 264506 -2776
rect 264742 -3012 264774 -2776
rect 264154 -3096 264774 -3012
rect 264154 -3332 264186 -3096
rect 264422 -3332 264506 -3096
rect 264742 -3332 264774 -3096
rect 264154 -4324 264774 -3332
rect 267874 463972 268494 464004
rect 267874 463736 267906 463972
rect 268142 463736 268226 463972
rect 268462 463736 268494 463972
rect 267874 463652 268494 463736
rect 267874 463416 267906 463652
rect 268142 463416 268226 463652
rect 268462 463416 268494 463652
rect 267874 448614 268494 463416
rect 267874 448378 267906 448614
rect 268142 448378 268226 448614
rect 268462 448378 268494 448614
rect 267874 448294 268494 448378
rect 267874 448058 267906 448294
rect 268142 448058 268226 448294
rect 268462 448058 268494 448294
rect 267874 430614 268494 448058
rect 267874 430378 267906 430614
rect 268142 430378 268226 430614
rect 268462 430378 268494 430614
rect 267874 430294 268494 430378
rect 267874 430058 267906 430294
rect 268142 430058 268226 430294
rect 268462 430058 268494 430294
rect 267874 412614 268494 430058
rect 267874 412378 267906 412614
rect 268142 412378 268226 412614
rect 268462 412378 268494 412614
rect 267874 412294 268494 412378
rect 267874 412058 267906 412294
rect 268142 412058 268226 412294
rect 268462 412058 268494 412294
rect 267874 394614 268494 412058
rect 267874 394378 267906 394614
rect 268142 394378 268226 394614
rect 268462 394378 268494 394614
rect 267874 394294 268494 394378
rect 267874 394058 267906 394294
rect 268142 394058 268226 394294
rect 268462 394058 268494 394294
rect 267874 376614 268494 394058
rect 267874 376378 267906 376614
rect 268142 376378 268226 376614
rect 268462 376378 268494 376614
rect 267874 376294 268494 376378
rect 267874 376058 267906 376294
rect 268142 376058 268226 376294
rect 268462 376058 268494 376294
rect 267874 358614 268494 376058
rect 267874 358378 267906 358614
rect 268142 358378 268226 358614
rect 268462 358378 268494 358614
rect 267874 358294 268494 358378
rect 267874 358058 267906 358294
rect 268142 358058 268226 358294
rect 268462 358058 268494 358294
rect 267874 340614 268494 358058
rect 267874 340378 267906 340614
rect 268142 340378 268226 340614
rect 268462 340378 268494 340614
rect 267874 340294 268494 340378
rect 267874 340058 267906 340294
rect 268142 340058 268226 340294
rect 268462 340058 268494 340294
rect 267874 322614 268494 340058
rect 267874 322378 267906 322614
rect 268142 322378 268226 322614
rect 268462 322378 268494 322614
rect 267874 322294 268494 322378
rect 267874 322058 267906 322294
rect 268142 322058 268226 322294
rect 268462 322058 268494 322294
rect 267874 304614 268494 322058
rect 267874 304378 267906 304614
rect 268142 304378 268226 304614
rect 268462 304378 268494 304614
rect 267874 304294 268494 304378
rect 267874 304058 267906 304294
rect 268142 304058 268226 304294
rect 268462 304058 268494 304294
rect 267874 286614 268494 304058
rect 267874 286378 267906 286614
rect 268142 286378 268226 286614
rect 268462 286378 268494 286614
rect 267874 286294 268494 286378
rect 267874 286058 267906 286294
rect 268142 286058 268226 286294
rect 268462 286058 268494 286294
rect 267874 268614 268494 286058
rect 267874 268378 267906 268614
rect 268142 268378 268226 268614
rect 268462 268378 268494 268614
rect 267874 268294 268494 268378
rect 267874 268058 267906 268294
rect 268142 268058 268226 268294
rect 268462 268058 268494 268294
rect 267874 250614 268494 268058
rect 267874 250378 267906 250614
rect 268142 250378 268226 250614
rect 268462 250378 268494 250614
rect 267874 250294 268494 250378
rect 267874 250058 267906 250294
rect 268142 250058 268226 250294
rect 268462 250058 268494 250294
rect 267874 232614 268494 250058
rect 267874 232378 267906 232614
rect 268142 232378 268226 232614
rect 268462 232378 268494 232614
rect 267874 232294 268494 232378
rect 267874 232058 267906 232294
rect 268142 232058 268226 232294
rect 268462 232058 268494 232294
rect 267874 214614 268494 232058
rect 267874 214378 267906 214614
rect 268142 214378 268226 214614
rect 268462 214378 268494 214614
rect 267874 214294 268494 214378
rect 267874 214058 267906 214294
rect 268142 214058 268226 214294
rect 268462 214058 268494 214294
rect 267874 196614 268494 214058
rect 267874 196378 267906 196614
rect 268142 196378 268226 196614
rect 268462 196378 268494 196614
rect 267874 196294 268494 196378
rect 267874 196058 267906 196294
rect 268142 196058 268226 196294
rect 268462 196058 268494 196294
rect 267874 178614 268494 196058
rect 267874 178378 267906 178614
rect 268142 178378 268226 178614
rect 268462 178378 268494 178614
rect 267874 178294 268494 178378
rect 267874 178058 267906 178294
rect 268142 178058 268226 178294
rect 268462 178058 268494 178294
rect 267874 160614 268494 178058
rect 267874 160378 267906 160614
rect 268142 160378 268226 160614
rect 268462 160378 268494 160614
rect 267874 160294 268494 160378
rect 267874 160058 267906 160294
rect 268142 160058 268226 160294
rect 268462 160058 268494 160294
rect 267874 142614 268494 160058
rect 267874 142378 267906 142614
rect 268142 142378 268226 142614
rect 268462 142378 268494 142614
rect 267874 142294 268494 142378
rect 267874 142058 267906 142294
rect 268142 142058 268226 142294
rect 268462 142058 268494 142294
rect 267874 124614 268494 142058
rect 267874 124378 267906 124614
rect 268142 124378 268226 124614
rect 268462 124378 268494 124614
rect 267874 124294 268494 124378
rect 267874 124058 267906 124294
rect 268142 124058 268226 124294
rect 268462 124058 268494 124294
rect 267874 106614 268494 124058
rect 267874 106378 267906 106614
rect 268142 106378 268226 106614
rect 268462 106378 268494 106614
rect 267874 106294 268494 106378
rect 267874 106058 267906 106294
rect 268142 106058 268226 106294
rect 268462 106058 268494 106294
rect 267874 88614 268494 106058
rect 267874 88378 267906 88614
rect 268142 88378 268226 88614
rect 268462 88378 268494 88614
rect 267874 88294 268494 88378
rect 267874 88058 267906 88294
rect 268142 88058 268226 88294
rect 268462 88058 268494 88294
rect 267874 70614 268494 88058
rect 267874 70378 267906 70614
rect 268142 70378 268226 70614
rect 268462 70378 268494 70614
rect 267874 70294 268494 70378
rect 267874 70058 267906 70294
rect 268142 70058 268226 70294
rect 268462 70058 268494 70294
rect 267874 52614 268494 70058
rect 267874 52378 267906 52614
rect 268142 52378 268226 52614
rect 268462 52378 268494 52614
rect 267874 52294 268494 52378
rect 267874 52058 267906 52294
rect 268142 52058 268226 52294
rect 268462 52058 268494 52294
rect 267874 34614 268494 52058
rect 267874 34378 267906 34614
rect 268142 34378 268226 34614
rect 268462 34378 268494 34614
rect 267874 34294 268494 34378
rect 267874 34058 267906 34294
rect 268142 34058 268226 34294
rect 268462 34058 268494 34294
rect 267874 16614 268494 34058
rect 267874 16378 267906 16614
rect 268142 16378 268226 16614
rect 268462 16378 268494 16614
rect 267874 16294 268494 16378
rect 267874 16058 267906 16294
rect 268142 16058 268226 16294
rect 268462 16058 268494 16294
rect 267874 -3736 268494 16058
rect 267874 -3972 267906 -3736
rect 268142 -3972 268226 -3736
rect 268462 -3972 268494 -3736
rect 267874 -4056 268494 -3972
rect 267874 -4292 267906 -4056
rect 268142 -4292 268226 -4056
rect 268462 -4292 268494 -4056
rect 267874 -4324 268494 -4292
rect 274714 461092 275334 464004
rect 274714 460856 274746 461092
rect 274982 460856 275066 461092
rect 275302 460856 275334 461092
rect 274714 460772 275334 460856
rect 274714 460536 274746 460772
rect 274982 460536 275066 460772
rect 275302 460536 275334 460772
rect 274714 455454 275334 460536
rect 274714 455218 274746 455454
rect 274982 455218 275066 455454
rect 275302 455218 275334 455454
rect 274714 455134 275334 455218
rect 274714 454898 274746 455134
rect 274982 454898 275066 455134
rect 275302 454898 275334 455134
rect 274714 437454 275334 454898
rect 274714 437218 274746 437454
rect 274982 437218 275066 437454
rect 275302 437218 275334 437454
rect 274714 437134 275334 437218
rect 274714 436898 274746 437134
rect 274982 436898 275066 437134
rect 275302 436898 275334 437134
rect 274714 419454 275334 436898
rect 274714 419218 274746 419454
rect 274982 419218 275066 419454
rect 275302 419218 275334 419454
rect 274714 419134 275334 419218
rect 274714 418898 274746 419134
rect 274982 418898 275066 419134
rect 275302 418898 275334 419134
rect 274714 401454 275334 418898
rect 274714 401218 274746 401454
rect 274982 401218 275066 401454
rect 275302 401218 275334 401454
rect 274714 401134 275334 401218
rect 274714 400898 274746 401134
rect 274982 400898 275066 401134
rect 275302 400898 275334 401134
rect 274714 383454 275334 400898
rect 274714 383218 274746 383454
rect 274982 383218 275066 383454
rect 275302 383218 275334 383454
rect 274714 383134 275334 383218
rect 274714 382898 274746 383134
rect 274982 382898 275066 383134
rect 275302 382898 275334 383134
rect 274714 365454 275334 382898
rect 274714 365218 274746 365454
rect 274982 365218 275066 365454
rect 275302 365218 275334 365454
rect 274714 365134 275334 365218
rect 274714 364898 274746 365134
rect 274982 364898 275066 365134
rect 275302 364898 275334 365134
rect 274714 347454 275334 364898
rect 274714 347218 274746 347454
rect 274982 347218 275066 347454
rect 275302 347218 275334 347454
rect 274714 347134 275334 347218
rect 274714 346898 274746 347134
rect 274982 346898 275066 347134
rect 275302 346898 275334 347134
rect 274714 329454 275334 346898
rect 274714 329218 274746 329454
rect 274982 329218 275066 329454
rect 275302 329218 275334 329454
rect 274714 329134 275334 329218
rect 274714 328898 274746 329134
rect 274982 328898 275066 329134
rect 275302 328898 275334 329134
rect 274714 311454 275334 328898
rect 274714 311218 274746 311454
rect 274982 311218 275066 311454
rect 275302 311218 275334 311454
rect 274714 311134 275334 311218
rect 274714 310898 274746 311134
rect 274982 310898 275066 311134
rect 275302 310898 275334 311134
rect 274714 293454 275334 310898
rect 274714 293218 274746 293454
rect 274982 293218 275066 293454
rect 275302 293218 275334 293454
rect 274714 293134 275334 293218
rect 274714 292898 274746 293134
rect 274982 292898 275066 293134
rect 275302 292898 275334 293134
rect 274714 275454 275334 292898
rect 274714 275218 274746 275454
rect 274982 275218 275066 275454
rect 275302 275218 275334 275454
rect 274714 275134 275334 275218
rect 274714 274898 274746 275134
rect 274982 274898 275066 275134
rect 275302 274898 275334 275134
rect 274714 257454 275334 274898
rect 274714 257218 274746 257454
rect 274982 257218 275066 257454
rect 275302 257218 275334 257454
rect 274714 257134 275334 257218
rect 274714 256898 274746 257134
rect 274982 256898 275066 257134
rect 275302 256898 275334 257134
rect 274714 239454 275334 256898
rect 274714 239218 274746 239454
rect 274982 239218 275066 239454
rect 275302 239218 275334 239454
rect 274714 239134 275334 239218
rect 274714 238898 274746 239134
rect 274982 238898 275066 239134
rect 275302 238898 275334 239134
rect 274714 221454 275334 238898
rect 274714 221218 274746 221454
rect 274982 221218 275066 221454
rect 275302 221218 275334 221454
rect 274714 221134 275334 221218
rect 274714 220898 274746 221134
rect 274982 220898 275066 221134
rect 275302 220898 275334 221134
rect 274714 203454 275334 220898
rect 274714 203218 274746 203454
rect 274982 203218 275066 203454
rect 275302 203218 275334 203454
rect 274714 203134 275334 203218
rect 274714 202898 274746 203134
rect 274982 202898 275066 203134
rect 275302 202898 275334 203134
rect 274714 185454 275334 202898
rect 274714 185218 274746 185454
rect 274982 185218 275066 185454
rect 275302 185218 275334 185454
rect 274714 185134 275334 185218
rect 274714 184898 274746 185134
rect 274982 184898 275066 185134
rect 275302 184898 275334 185134
rect 274714 167454 275334 184898
rect 274714 167218 274746 167454
rect 274982 167218 275066 167454
rect 275302 167218 275334 167454
rect 274714 167134 275334 167218
rect 274714 166898 274746 167134
rect 274982 166898 275066 167134
rect 275302 166898 275334 167134
rect 274714 149454 275334 166898
rect 274714 149218 274746 149454
rect 274982 149218 275066 149454
rect 275302 149218 275334 149454
rect 274714 149134 275334 149218
rect 274714 148898 274746 149134
rect 274982 148898 275066 149134
rect 275302 148898 275334 149134
rect 274714 131454 275334 148898
rect 274714 131218 274746 131454
rect 274982 131218 275066 131454
rect 275302 131218 275334 131454
rect 274714 131134 275334 131218
rect 274714 130898 274746 131134
rect 274982 130898 275066 131134
rect 275302 130898 275334 131134
rect 274714 113454 275334 130898
rect 274714 113218 274746 113454
rect 274982 113218 275066 113454
rect 275302 113218 275334 113454
rect 274714 113134 275334 113218
rect 274714 112898 274746 113134
rect 274982 112898 275066 113134
rect 275302 112898 275334 113134
rect 274714 95454 275334 112898
rect 274714 95218 274746 95454
rect 274982 95218 275066 95454
rect 275302 95218 275334 95454
rect 274714 95134 275334 95218
rect 274714 94898 274746 95134
rect 274982 94898 275066 95134
rect 275302 94898 275334 95134
rect 274714 77454 275334 94898
rect 274714 77218 274746 77454
rect 274982 77218 275066 77454
rect 275302 77218 275334 77454
rect 274714 77134 275334 77218
rect 274714 76898 274746 77134
rect 274982 76898 275066 77134
rect 275302 76898 275334 77134
rect 274714 59454 275334 76898
rect 274714 59218 274746 59454
rect 274982 59218 275066 59454
rect 275302 59218 275334 59454
rect 274714 59134 275334 59218
rect 274714 58898 274746 59134
rect 274982 58898 275066 59134
rect 275302 58898 275334 59134
rect 274714 41454 275334 58898
rect 274714 41218 274746 41454
rect 274982 41218 275066 41454
rect 275302 41218 275334 41454
rect 274714 41134 275334 41218
rect 274714 40898 274746 41134
rect 274982 40898 275066 41134
rect 275302 40898 275334 41134
rect 274714 23454 275334 40898
rect 274714 23218 274746 23454
rect 274982 23218 275066 23454
rect 275302 23218 275334 23454
rect 274714 23134 275334 23218
rect 274714 22898 274746 23134
rect 274982 22898 275066 23134
rect 275302 22898 275334 23134
rect 274714 5454 275334 22898
rect 274714 5218 274746 5454
rect 274982 5218 275066 5454
rect 275302 5218 275334 5454
rect 274714 5134 275334 5218
rect 274714 4898 274746 5134
rect 274982 4898 275066 5134
rect 275302 4898 275334 5134
rect 274714 -856 275334 4898
rect 274714 -1092 274746 -856
rect 274982 -1092 275066 -856
rect 275302 -1092 275334 -856
rect 274714 -1176 275334 -1092
rect 274714 -1412 274746 -1176
rect 274982 -1412 275066 -1176
rect 275302 -1412 275334 -1176
rect 274714 -4324 275334 -1412
rect 278434 462052 279054 464004
rect 278434 461816 278466 462052
rect 278702 461816 278786 462052
rect 279022 461816 279054 462052
rect 278434 461732 279054 461816
rect 278434 461496 278466 461732
rect 278702 461496 278786 461732
rect 279022 461496 279054 461732
rect 278434 441174 279054 461496
rect 278434 440938 278466 441174
rect 278702 440938 278786 441174
rect 279022 440938 279054 441174
rect 278434 440854 279054 440938
rect 278434 440618 278466 440854
rect 278702 440618 278786 440854
rect 279022 440618 279054 440854
rect 278434 423174 279054 440618
rect 278434 422938 278466 423174
rect 278702 422938 278786 423174
rect 279022 422938 279054 423174
rect 278434 422854 279054 422938
rect 278434 422618 278466 422854
rect 278702 422618 278786 422854
rect 279022 422618 279054 422854
rect 278434 405174 279054 422618
rect 278434 404938 278466 405174
rect 278702 404938 278786 405174
rect 279022 404938 279054 405174
rect 278434 404854 279054 404938
rect 278434 404618 278466 404854
rect 278702 404618 278786 404854
rect 279022 404618 279054 404854
rect 278434 387174 279054 404618
rect 278434 386938 278466 387174
rect 278702 386938 278786 387174
rect 279022 386938 279054 387174
rect 278434 386854 279054 386938
rect 278434 386618 278466 386854
rect 278702 386618 278786 386854
rect 279022 386618 279054 386854
rect 278434 369174 279054 386618
rect 278434 368938 278466 369174
rect 278702 368938 278786 369174
rect 279022 368938 279054 369174
rect 278434 368854 279054 368938
rect 278434 368618 278466 368854
rect 278702 368618 278786 368854
rect 279022 368618 279054 368854
rect 278434 351174 279054 368618
rect 278434 350938 278466 351174
rect 278702 350938 278786 351174
rect 279022 350938 279054 351174
rect 278434 350854 279054 350938
rect 278434 350618 278466 350854
rect 278702 350618 278786 350854
rect 279022 350618 279054 350854
rect 278434 333174 279054 350618
rect 278434 332938 278466 333174
rect 278702 332938 278786 333174
rect 279022 332938 279054 333174
rect 278434 332854 279054 332938
rect 278434 332618 278466 332854
rect 278702 332618 278786 332854
rect 279022 332618 279054 332854
rect 278434 315174 279054 332618
rect 278434 314938 278466 315174
rect 278702 314938 278786 315174
rect 279022 314938 279054 315174
rect 278434 314854 279054 314938
rect 278434 314618 278466 314854
rect 278702 314618 278786 314854
rect 279022 314618 279054 314854
rect 278434 297174 279054 314618
rect 278434 296938 278466 297174
rect 278702 296938 278786 297174
rect 279022 296938 279054 297174
rect 278434 296854 279054 296938
rect 278434 296618 278466 296854
rect 278702 296618 278786 296854
rect 279022 296618 279054 296854
rect 278434 279174 279054 296618
rect 278434 278938 278466 279174
rect 278702 278938 278786 279174
rect 279022 278938 279054 279174
rect 278434 278854 279054 278938
rect 278434 278618 278466 278854
rect 278702 278618 278786 278854
rect 279022 278618 279054 278854
rect 278434 261174 279054 278618
rect 278434 260938 278466 261174
rect 278702 260938 278786 261174
rect 279022 260938 279054 261174
rect 278434 260854 279054 260938
rect 278434 260618 278466 260854
rect 278702 260618 278786 260854
rect 279022 260618 279054 260854
rect 278434 243174 279054 260618
rect 278434 242938 278466 243174
rect 278702 242938 278786 243174
rect 279022 242938 279054 243174
rect 278434 242854 279054 242938
rect 278434 242618 278466 242854
rect 278702 242618 278786 242854
rect 279022 242618 279054 242854
rect 278434 225174 279054 242618
rect 278434 224938 278466 225174
rect 278702 224938 278786 225174
rect 279022 224938 279054 225174
rect 278434 224854 279054 224938
rect 278434 224618 278466 224854
rect 278702 224618 278786 224854
rect 279022 224618 279054 224854
rect 278434 207174 279054 224618
rect 278434 206938 278466 207174
rect 278702 206938 278786 207174
rect 279022 206938 279054 207174
rect 278434 206854 279054 206938
rect 278434 206618 278466 206854
rect 278702 206618 278786 206854
rect 279022 206618 279054 206854
rect 278434 189174 279054 206618
rect 278434 188938 278466 189174
rect 278702 188938 278786 189174
rect 279022 188938 279054 189174
rect 278434 188854 279054 188938
rect 278434 188618 278466 188854
rect 278702 188618 278786 188854
rect 279022 188618 279054 188854
rect 278434 171174 279054 188618
rect 278434 170938 278466 171174
rect 278702 170938 278786 171174
rect 279022 170938 279054 171174
rect 278434 170854 279054 170938
rect 278434 170618 278466 170854
rect 278702 170618 278786 170854
rect 279022 170618 279054 170854
rect 278434 153174 279054 170618
rect 278434 152938 278466 153174
rect 278702 152938 278786 153174
rect 279022 152938 279054 153174
rect 278434 152854 279054 152938
rect 278434 152618 278466 152854
rect 278702 152618 278786 152854
rect 279022 152618 279054 152854
rect 278434 135174 279054 152618
rect 278434 134938 278466 135174
rect 278702 134938 278786 135174
rect 279022 134938 279054 135174
rect 278434 134854 279054 134938
rect 278434 134618 278466 134854
rect 278702 134618 278786 134854
rect 279022 134618 279054 134854
rect 278434 117174 279054 134618
rect 278434 116938 278466 117174
rect 278702 116938 278786 117174
rect 279022 116938 279054 117174
rect 278434 116854 279054 116938
rect 278434 116618 278466 116854
rect 278702 116618 278786 116854
rect 279022 116618 279054 116854
rect 278434 99174 279054 116618
rect 278434 98938 278466 99174
rect 278702 98938 278786 99174
rect 279022 98938 279054 99174
rect 278434 98854 279054 98938
rect 278434 98618 278466 98854
rect 278702 98618 278786 98854
rect 279022 98618 279054 98854
rect 278434 81174 279054 98618
rect 278434 80938 278466 81174
rect 278702 80938 278786 81174
rect 279022 80938 279054 81174
rect 278434 80854 279054 80938
rect 278434 80618 278466 80854
rect 278702 80618 278786 80854
rect 279022 80618 279054 80854
rect 278434 63174 279054 80618
rect 278434 62938 278466 63174
rect 278702 62938 278786 63174
rect 279022 62938 279054 63174
rect 278434 62854 279054 62938
rect 278434 62618 278466 62854
rect 278702 62618 278786 62854
rect 279022 62618 279054 62854
rect 278434 45174 279054 62618
rect 278434 44938 278466 45174
rect 278702 44938 278786 45174
rect 279022 44938 279054 45174
rect 278434 44854 279054 44938
rect 278434 44618 278466 44854
rect 278702 44618 278786 44854
rect 279022 44618 279054 44854
rect 278434 27174 279054 44618
rect 278434 26938 278466 27174
rect 278702 26938 278786 27174
rect 279022 26938 279054 27174
rect 278434 26854 279054 26938
rect 278434 26618 278466 26854
rect 278702 26618 278786 26854
rect 279022 26618 279054 26854
rect 278434 9174 279054 26618
rect 278434 8938 278466 9174
rect 278702 8938 278786 9174
rect 279022 8938 279054 9174
rect 278434 8854 279054 8938
rect 278434 8618 278466 8854
rect 278702 8618 278786 8854
rect 279022 8618 279054 8854
rect 278434 -1816 279054 8618
rect 278434 -2052 278466 -1816
rect 278702 -2052 278786 -1816
rect 279022 -2052 279054 -1816
rect 278434 -2136 279054 -2052
rect 278434 -2372 278466 -2136
rect 278702 -2372 278786 -2136
rect 279022 -2372 279054 -2136
rect 278434 -4324 279054 -2372
rect 282154 463012 282774 464004
rect 282154 462776 282186 463012
rect 282422 462776 282506 463012
rect 282742 462776 282774 463012
rect 282154 462692 282774 462776
rect 282154 462456 282186 462692
rect 282422 462456 282506 462692
rect 282742 462456 282774 462692
rect 282154 444894 282774 462456
rect 282154 444658 282186 444894
rect 282422 444658 282506 444894
rect 282742 444658 282774 444894
rect 282154 444574 282774 444658
rect 282154 444338 282186 444574
rect 282422 444338 282506 444574
rect 282742 444338 282774 444574
rect 282154 426894 282774 444338
rect 282154 426658 282186 426894
rect 282422 426658 282506 426894
rect 282742 426658 282774 426894
rect 282154 426574 282774 426658
rect 282154 426338 282186 426574
rect 282422 426338 282506 426574
rect 282742 426338 282774 426574
rect 282154 408894 282774 426338
rect 282154 408658 282186 408894
rect 282422 408658 282506 408894
rect 282742 408658 282774 408894
rect 282154 408574 282774 408658
rect 282154 408338 282186 408574
rect 282422 408338 282506 408574
rect 282742 408338 282774 408574
rect 282154 390894 282774 408338
rect 282154 390658 282186 390894
rect 282422 390658 282506 390894
rect 282742 390658 282774 390894
rect 282154 390574 282774 390658
rect 282154 390338 282186 390574
rect 282422 390338 282506 390574
rect 282742 390338 282774 390574
rect 282154 372894 282774 390338
rect 282154 372658 282186 372894
rect 282422 372658 282506 372894
rect 282742 372658 282774 372894
rect 282154 372574 282774 372658
rect 282154 372338 282186 372574
rect 282422 372338 282506 372574
rect 282742 372338 282774 372574
rect 282154 354894 282774 372338
rect 282154 354658 282186 354894
rect 282422 354658 282506 354894
rect 282742 354658 282774 354894
rect 282154 354574 282774 354658
rect 282154 354338 282186 354574
rect 282422 354338 282506 354574
rect 282742 354338 282774 354574
rect 282154 336894 282774 354338
rect 282154 336658 282186 336894
rect 282422 336658 282506 336894
rect 282742 336658 282774 336894
rect 282154 336574 282774 336658
rect 282154 336338 282186 336574
rect 282422 336338 282506 336574
rect 282742 336338 282774 336574
rect 282154 318894 282774 336338
rect 282154 318658 282186 318894
rect 282422 318658 282506 318894
rect 282742 318658 282774 318894
rect 282154 318574 282774 318658
rect 282154 318338 282186 318574
rect 282422 318338 282506 318574
rect 282742 318338 282774 318574
rect 282154 300894 282774 318338
rect 282154 300658 282186 300894
rect 282422 300658 282506 300894
rect 282742 300658 282774 300894
rect 282154 300574 282774 300658
rect 282154 300338 282186 300574
rect 282422 300338 282506 300574
rect 282742 300338 282774 300574
rect 282154 282894 282774 300338
rect 282154 282658 282186 282894
rect 282422 282658 282506 282894
rect 282742 282658 282774 282894
rect 282154 282574 282774 282658
rect 282154 282338 282186 282574
rect 282422 282338 282506 282574
rect 282742 282338 282774 282574
rect 282154 264894 282774 282338
rect 282154 264658 282186 264894
rect 282422 264658 282506 264894
rect 282742 264658 282774 264894
rect 282154 264574 282774 264658
rect 282154 264338 282186 264574
rect 282422 264338 282506 264574
rect 282742 264338 282774 264574
rect 282154 246894 282774 264338
rect 282154 246658 282186 246894
rect 282422 246658 282506 246894
rect 282742 246658 282774 246894
rect 282154 246574 282774 246658
rect 282154 246338 282186 246574
rect 282422 246338 282506 246574
rect 282742 246338 282774 246574
rect 282154 228894 282774 246338
rect 282154 228658 282186 228894
rect 282422 228658 282506 228894
rect 282742 228658 282774 228894
rect 282154 228574 282774 228658
rect 282154 228338 282186 228574
rect 282422 228338 282506 228574
rect 282742 228338 282774 228574
rect 282154 210894 282774 228338
rect 282154 210658 282186 210894
rect 282422 210658 282506 210894
rect 282742 210658 282774 210894
rect 282154 210574 282774 210658
rect 282154 210338 282186 210574
rect 282422 210338 282506 210574
rect 282742 210338 282774 210574
rect 282154 192894 282774 210338
rect 282154 192658 282186 192894
rect 282422 192658 282506 192894
rect 282742 192658 282774 192894
rect 282154 192574 282774 192658
rect 282154 192338 282186 192574
rect 282422 192338 282506 192574
rect 282742 192338 282774 192574
rect 282154 174894 282774 192338
rect 282154 174658 282186 174894
rect 282422 174658 282506 174894
rect 282742 174658 282774 174894
rect 282154 174574 282774 174658
rect 282154 174338 282186 174574
rect 282422 174338 282506 174574
rect 282742 174338 282774 174574
rect 282154 156894 282774 174338
rect 282154 156658 282186 156894
rect 282422 156658 282506 156894
rect 282742 156658 282774 156894
rect 282154 156574 282774 156658
rect 282154 156338 282186 156574
rect 282422 156338 282506 156574
rect 282742 156338 282774 156574
rect 282154 138894 282774 156338
rect 282154 138658 282186 138894
rect 282422 138658 282506 138894
rect 282742 138658 282774 138894
rect 282154 138574 282774 138658
rect 282154 138338 282186 138574
rect 282422 138338 282506 138574
rect 282742 138338 282774 138574
rect 282154 120894 282774 138338
rect 282154 120658 282186 120894
rect 282422 120658 282506 120894
rect 282742 120658 282774 120894
rect 282154 120574 282774 120658
rect 282154 120338 282186 120574
rect 282422 120338 282506 120574
rect 282742 120338 282774 120574
rect 282154 102894 282774 120338
rect 282154 102658 282186 102894
rect 282422 102658 282506 102894
rect 282742 102658 282774 102894
rect 282154 102574 282774 102658
rect 282154 102338 282186 102574
rect 282422 102338 282506 102574
rect 282742 102338 282774 102574
rect 282154 84894 282774 102338
rect 282154 84658 282186 84894
rect 282422 84658 282506 84894
rect 282742 84658 282774 84894
rect 282154 84574 282774 84658
rect 282154 84338 282186 84574
rect 282422 84338 282506 84574
rect 282742 84338 282774 84574
rect 282154 66894 282774 84338
rect 282154 66658 282186 66894
rect 282422 66658 282506 66894
rect 282742 66658 282774 66894
rect 282154 66574 282774 66658
rect 282154 66338 282186 66574
rect 282422 66338 282506 66574
rect 282742 66338 282774 66574
rect 282154 48894 282774 66338
rect 282154 48658 282186 48894
rect 282422 48658 282506 48894
rect 282742 48658 282774 48894
rect 282154 48574 282774 48658
rect 282154 48338 282186 48574
rect 282422 48338 282506 48574
rect 282742 48338 282774 48574
rect 282154 30894 282774 48338
rect 282154 30658 282186 30894
rect 282422 30658 282506 30894
rect 282742 30658 282774 30894
rect 282154 30574 282774 30658
rect 282154 30338 282186 30574
rect 282422 30338 282506 30574
rect 282742 30338 282774 30574
rect 282154 12894 282774 30338
rect 282154 12658 282186 12894
rect 282422 12658 282506 12894
rect 282742 12658 282774 12894
rect 282154 12574 282774 12658
rect 282154 12338 282186 12574
rect 282422 12338 282506 12574
rect 282742 12338 282774 12574
rect 282154 -2776 282774 12338
rect 282154 -3012 282186 -2776
rect 282422 -3012 282506 -2776
rect 282742 -3012 282774 -2776
rect 282154 -3096 282774 -3012
rect 282154 -3332 282186 -3096
rect 282422 -3332 282506 -3096
rect 282742 -3332 282774 -3096
rect 282154 -4324 282774 -3332
rect 285874 463972 286494 464004
rect 285874 463736 285906 463972
rect 286142 463736 286226 463972
rect 286462 463736 286494 463972
rect 285874 463652 286494 463736
rect 285874 463416 285906 463652
rect 286142 463416 286226 463652
rect 286462 463416 286494 463652
rect 285874 448614 286494 463416
rect 285874 448378 285906 448614
rect 286142 448378 286226 448614
rect 286462 448378 286494 448614
rect 285874 448294 286494 448378
rect 285874 448058 285906 448294
rect 286142 448058 286226 448294
rect 286462 448058 286494 448294
rect 285874 430614 286494 448058
rect 285874 430378 285906 430614
rect 286142 430378 286226 430614
rect 286462 430378 286494 430614
rect 285874 430294 286494 430378
rect 285874 430058 285906 430294
rect 286142 430058 286226 430294
rect 286462 430058 286494 430294
rect 285874 412614 286494 430058
rect 285874 412378 285906 412614
rect 286142 412378 286226 412614
rect 286462 412378 286494 412614
rect 285874 412294 286494 412378
rect 285874 412058 285906 412294
rect 286142 412058 286226 412294
rect 286462 412058 286494 412294
rect 285874 394614 286494 412058
rect 285874 394378 285906 394614
rect 286142 394378 286226 394614
rect 286462 394378 286494 394614
rect 285874 394294 286494 394378
rect 285874 394058 285906 394294
rect 286142 394058 286226 394294
rect 286462 394058 286494 394294
rect 285874 376614 286494 394058
rect 285874 376378 285906 376614
rect 286142 376378 286226 376614
rect 286462 376378 286494 376614
rect 285874 376294 286494 376378
rect 285874 376058 285906 376294
rect 286142 376058 286226 376294
rect 286462 376058 286494 376294
rect 285874 358614 286494 376058
rect 285874 358378 285906 358614
rect 286142 358378 286226 358614
rect 286462 358378 286494 358614
rect 285874 358294 286494 358378
rect 285874 358058 285906 358294
rect 286142 358058 286226 358294
rect 286462 358058 286494 358294
rect 285874 340614 286494 358058
rect 285874 340378 285906 340614
rect 286142 340378 286226 340614
rect 286462 340378 286494 340614
rect 285874 340294 286494 340378
rect 285874 340058 285906 340294
rect 286142 340058 286226 340294
rect 286462 340058 286494 340294
rect 285874 322614 286494 340058
rect 285874 322378 285906 322614
rect 286142 322378 286226 322614
rect 286462 322378 286494 322614
rect 285874 322294 286494 322378
rect 285874 322058 285906 322294
rect 286142 322058 286226 322294
rect 286462 322058 286494 322294
rect 285874 304614 286494 322058
rect 285874 304378 285906 304614
rect 286142 304378 286226 304614
rect 286462 304378 286494 304614
rect 285874 304294 286494 304378
rect 285874 304058 285906 304294
rect 286142 304058 286226 304294
rect 286462 304058 286494 304294
rect 285874 286614 286494 304058
rect 285874 286378 285906 286614
rect 286142 286378 286226 286614
rect 286462 286378 286494 286614
rect 285874 286294 286494 286378
rect 285874 286058 285906 286294
rect 286142 286058 286226 286294
rect 286462 286058 286494 286294
rect 285874 268614 286494 286058
rect 285874 268378 285906 268614
rect 286142 268378 286226 268614
rect 286462 268378 286494 268614
rect 285874 268294 286494 268378
rect 285874 268058 285906 268294
rect 286142 268058 286226 268294
rect 286462 268058 286494 268294
rect 285874 250614 286494 268058
rect 285874 250378 285906 250614
rect 286142 250378 286226 250614
rect 286462 250378 286494 250614
rect 285874 250294 286494 250378
rect 285874 250058 285906 250294
rect 286142 250058 286226 250294
rect 286462 250058 286494 250294
rect 285874 232614 286494 250058
rect 285874 232378 285906 232614
rect 286142 232378 286226 232614
rect 286462 232378 286494 232614
rect 285874 232294 286494 232378
rect 285874 232058 285906 232294
rect 286142 232058 286226 232294
rect 286462 232058 286494 232294
rect 285874 214614 286494 232058
rect 285874 214378 285906 214614
rect 286142 214378 286226 214614
rect 286462 214378 286494 214614
rect 285874 214294 286494 214378
rect 285874 214058 285906 214294
rect 286142 214058 286226 214294
rect 286462 214058 286494 214294
rect 285874 196614 286494 214058
rect 285874 196378 285906 196614
rect 286142 196378 286226 196614
rect 286462 196378 286494 196614
rect 285874 196294 286494 196378
rect 285874 196058 285906 196294
rect 286142 196058 286226 196294
rect 286462 196058 286494 196294
rect 285874 178614 286494 196058
rect 285874 178378 285906 178614
rect 286142 178378 286226 178614
rect 286462 178378 286494 178614
rect 285874 178294 286494 178378
rect 285874 178058 285906 178294
rect 286142 178058 286226 178294
rect 286462 178058 286494 178294
rect 285874 160614 286494 178058
rect 285874 160378 285906 160614
rect 286142 160378 286226 160614
rect 286462 160378 286494 160614
rect 285874 160294 286494 160378
rect 285874 160058 285906 160294
rect 286142 160058 286226 160294
rect 286462 160058 286494 160294
rect 285874 142614 286494 160058
rect 285874 142378 285906 142614
rect 286142 142378 286226 142614
rect 286462 142378 286494 142614
rect 285874 142294 286494 142378
rect 285874 142058 285906 142294
rect 286142 142058 286226 142294
rect 286462 142058 286494 142294
rect 285874 124614 286494 142058
rect 285874 124378 285906 124614
rect 286142 124378 286226 124614
rect 286462 124378 286494 124614
rect 285874 124294 286494 124378
rect 285874 124058 285906 124294
rect 286142 124058 286226 124294
rect 286462 124058 286494 124294
rect 285874 106614 286494 124058
rect 285874 106378 285906 106614
rect 286142 106378 286226 106614
rect 286462 106378 286494 106614
rect 285874 106294 286494 106378
rect 285874 106058 285906 106294
rect 286142 106058 286226 106294
rect 286462 106058 286494 106294
rect 285874 88614 286494 106058
rect 285874 88378 285906 88614
rect 286142 88378 286226 88614
rect 286462 88378 286494 88614
rect 285874 88294 286494 88378
rect 285874 88058 285906 88294
rect 286142 88058 286226 88294
rect 286462 88058 286494 88294
rect 285874 70614 286494 88058
rect 285874 70378 285906 70614
rect 286142 70378 286226 70614
rect 286462 70378 286494 70614
rect 285874 70294 286494 70378
rect 285874 70058 285906 70294
rect 286142 70058 286226 70294
rect 286462 70058 286494 70294
rect 285874 52614 286494 70058
rect 285874 52378 285906 52614
rect 286142 52378 286226 52614
rect 286462 52378 286494 52614
rect 285874 52294 286494 52378
rect 285874 52058 285906 52294
rect 286142 52058 286226 52294
rect 286462 52058 286494 52294
rect 285874 34614 286494 52058
rect 285874 34378 285906 34614
rect 286142 34378 286226 34614
rect 286462 34378 286494 34614
rect 285874 34294 286494 34378
rect 285874 34058 285906 34294
rect 286142 34058 286226 34294
rect 286462 34058 286494 34294
rect 285874 16614 286494 34058
rect 285874 16378 285906 16614
rect 286142 16378 286226 16614
rect 286462 16378 286494 16614
rect 285874 16294 286494 16378
rect 285874 16058 285906 16294
rect 286142 16058 286226 16294
rect 286462 16058 286494 16294
rect 285874 -3736 286494 16058
rect 285874 -3972 285906 -3736
rect 286142 -3972 286226 -3736
rect 286462 -3972 286494 -3736
rect 285874 -4056 286494 -3972
rect 285874 -4292 285906 -4056
rect 286142 -4292 286226 -4056
rect 286462 -4292 286494 -4056
rect 285874 -4324 286494 -4292
rect 292714 461092 293334 464004
rect 292714 460856 292746 461092
rect 292982 460856 293066 461092
rect 293302 460856 293334 461092
rect 292714 460772 293334 460856
rect 292714 460536 292746 460772
rect 292982 460536 293066 460772
rect 293302 460536 293334 460772
rect 292714 455454 293334 460536
rect 292714 455218 292746 455454
rect 292982 455218 293066 455454
rect 293302 455218 293334 455454
rect 292714 455134 293334 455218
rect 292714 454898 292746 455134
rect 292982 454898 293066 455134
rect 293302 454898 293334 455134
rect 292714 437454 293334 454898
rect 292714 437218 292746 437454
rect 292982 437218 293066 437454
rect 293302 437218 293334 437454
rect 292714 437134 293334 437218
rect 292714 436898 292746 437134
rect 292982 436898 293066 437134
rect 293302 436898 293334 437134
rect 292714 419454 293334 436898
rect 292714 419218 292746 419454
rect 292982 419218 293066 419454
rect 293302 419218 293334 419454
rect 292714 419134 293334 419218
rect 292714 418898 292746 419134
rect 292982 418898 293066 419134
rect 293302 418898 293334 419134
rect 292714 401454 293334 418898
rect 292714 401218 292746 401454
rect 292982 401218 293066 401454
rect 293302 401218 293334 401454
rect 292714 401134 293334 401218
rect 292714 400898 292746 401134
rect 292982 400898 293066 401134
rect 293302 400898 293334 401134
rect 292714 383454 293334 400898
rect 292714 383218 292746 383454
rect 292982 383218 293066 383454
rect 293302 383218 293334 383454
rect 292714 383134 293334 383218
rect 292714 382898 292746 383134
rect 292982 382898 293066 383134
rect 293302 382898 293334 383134
rect 292714 365454 293334 382898
rect 292714 365218 292746 365454
rect 292982 365218 293066 365454
rect 293302 365218 293334 365454
rect 292714 365134 293334 365218
rect 292714 364898 292746 365134
rect 292982 364898 293066 365134
rect 293302 364898 293334 365134
rect 292714 347454 293334 364898
rect 292714 347218 292746 347454
rect 292982 347218 293066 347454
rect 293302 347218 293334 347454
rect 292714 347134 293334 347218
rect 292714 346898 292746 347134
rect 292982 346898 293066 347134
rect 293302 346898 293334 347134
rect 292714 329454 293334 346898
rect 292714 329218 292746 329454
rect 292982 329218 293066 329454
rect 293302 329218 293334 329454
rect 292714 329134 293334 329218
rect 292714 328898 292746 329134
rect 292982 328898 293066 329134
rect 293302 328898 293334 329134
rect 292714 311454 293334 328898
rect 292714 311218 292746 311454
rect 292982 311218 293066 311454
rect 293302 311218 293334 311454
rect 292714 311134 293334 311218
rect 292714 310898 292746 311134
rect 292982 310898 293066 311134
rect 293302 310898 293334 311134
rect 292714 293454 293334 310898
rect 292714 293218 292746 293454
rect 292982 293218 293066 293454
rect 293302 293218 293334 293454
rect 292714 293134 293334 293218
rect 292714 292898 292746 293134
rect 292982 292898 293066 293134
rect 293302 292898 293334 293134
rect 292714 275454 293334 292898
rect 292714 275218 292746 275454
rect 292982 275218 293066 275454
rect 293302 275218 293334 275454
rect 292714 275134 293334 275218
rect 292714 274898 292746 275134
rect 292982 274898 293066 275134
rect 293302 274898 293334 275134
rect 292714 257454 293334 274898
rect 292714 257218 292746 257454
rect 292982 257218 293066 257454
rect 293302 257218 293334 257454
rect 292714 257134 293334 257218
rect 292714 256898 292746 257134
rect 292982 256898 293066 257134
rect 293302 256898 293334 257134
rect 292714 239454 293334 256898
rect 292714 239218 292746 239454
rect 292982 239218 293066 239454
rect 293302 239218 293334 239454
rect 292714 239134 293334 239218
rect 292714 238898 292746 239134
rect 292982 238898 293066 239134
rect 293302 238898 293334 239134
rect 292714 221454 293334 238898
rect 292714 221218 292746 221454
rect 292982 221218 293066 221454
rect 293302 221218 293334 221454
rect 292714 221134 293334 221218
rect 292714 220898 292746 221134
rect 292982 220898 293066 221134
rect 293302 220898 293334 221134
rect 292714 203454 293334 220898
rect 292714 203218 292746 203454
rect 292982 203218 293066 203454
rect 293302 203218 293334 203454
rect 292714 203134 293334 203218
rect 292714 202898 292746 203134
rect 292982 202898 293066 203134
rect 293302 202898 293334 203134
rect 292714 185454 293334 202898
rect 292714 185218 292746 185454
rect 292982 185218 293066 185454
rect 293302 185218 293334 185454
rect 292714 185134 293334 185218
rect 292714 184898 292746 185134
rect 292982 184898 293066 185134
rect 293302 184898 293334 185134
rect 292714 167454 293334 184898
rect 292714 167218 292746 167454
rect 292982 167218 293066 167454
rect 293302 167218 293334 167454
rect 292714 167134 293334 167218
rect 292714 166898 292746 167134
rect 292982 166898 293066 167134
rect 293302 166898 293334 167134
rect 292714 149454 293334 166898
rect 292714 149218 292746 149454
rect 292982 149218 293066 149454
rect 293302 149218 293334 149454
rect 292714 149134 293334 149218
rect 292714 148898 292746 149134
rect 292982 148898 293066 149134
rect 293302 148898 293334 149134
rect 292714 131454 293334 148898
rect 292714 131218 292746 131454
rect 292982 131218 293066 131454
rect 293302 131218 293334 131454
rect 292714 131134 293334 131218
rect 292714 130898 292746 131134
rect 292982 130898 293066 131134
rect 293302 130898 293334 131134
rect 292714 113454 293334 130898
rect 292714 113218 292746 113454
rect 292982 113218 293066 113454
rect 293302 113218 293334 113454
rect 292714 113134 293334 113218
rect 292714 112898 292746 113134
rect 292982 112898 293066 113134
rect 293302 112898 293334 113134
rect 292714 95454 293334 112898
rect 292714 95218 292746 95454
rect 292982 95218 293066 95454
rect 293302 95218 293334 95454
rect 292714 95134 293334 95218
rect 292714 94898 292746 95134
rect 292982 94898 293066 95134
rect 293302 94898 293334 95134
rect 292714 77454 293334 94898
rect 292714 77218 292746 77454
rect 292982 77218 293066 77454
rect 293302 77218 293334 77454
rect 292714 77134 293334 77218
rect 292714 76898 292746 77134
rect 292982 76898 293066 77134
rect 293302 76898 293334 77134
rect 292714 59454 293334 76898
rect 292714 59218 292746 59454
rect 292982 59218 293066 59454
rect 293302 59218 293334 59454
rect 292714 59134 293334 59218
rect 292714 58898 292746 59134
rect 292982 58898 293066 59134
rect 293302 58898 293334 59134
rect 292714 41454 293334 58898
rect 292714 41218 292746 41454
rect 292982 41218 293066 41454
rect 293302 41218 293334 41454
rect 292714 41134 293334 41218
rect 292714 40898 292746 41134
rect 292982 40898 293066 41134
rect 293302 40898 293334 41134
rect 292714 23454 293334 40898
rect 292714 23218 292746 23454
rect 292982 23218 293066 23454
rect 293302 23218 293334 23454
rect 292714 23134 293334 23218
rect 292714 22898 292746 23134
rect 292982 22898 293066 23134
rect 293302 22898 293334 23134
rect 292714 5454 293334 22898
rect 292714 5218 292746 5454
rect 292982 5218 293066 5454
rect 293302 5218 293334 5454
rect 292714 5134 293334 5218
rect 292714 4898 292746 5134
rect 292982 4898 293066 5134
rect 293302 4898 293334 5134
rect 292714 -856 293334 4898
rect 292714 -1092 292746 -856
rect 292982 -1092 293066 -856
rect 293302 -1092 293334 -856
rect 292714 -1176 293334 -1092
rect 292714 -1412 292746 -1176
rect 292982 -1412 293066 -1176
rect 293302 -1412 293334 -1176
rect 292714 -4324 293334 -1412
rect 296434 462052 297054 464004
rect 296434 461816 296466 462052
rect 296702 461816 296786 462052
rect 297022 461816 297054 462052
rect 296434 461732 297054 461816
rect 296434 461496 296466 461732
rect 296702 461496 296786 461732
rect 297022 461496 297054 461732
rect 296434 441174 297054 461496
rect 296434 440938 296466 441174
rect 296702 440938 296786 441174
rect 297022 440938 297054 441174
rect 296434 440854 297054 440938
rect 296434 440618 296466 440854
rect 296702 440618 296786 440854
rect 297022 440618 297054 440854
rect 296434 423174 297054 440618
rect 296434 422938 296466 423174
rect 296702 422938 296786 423174
rect 297022 422938 297054 423174
rect 296434 422854 297054 422938
rect 296434 422618 296466 422854
rect 296702 422618 296786 422854
rect 297022 422618 297054 422854
rect 296434 405174 297054 422618
rect 296434 404938 296466 405174
rect 296702 404938 296786 405174
rect 297022 404938 297054 405174
rect 296434 404854 297054 404938
rect 296434 404618 296466 404854
rect 296702 404618 296786 404854
rect 297022 404618 297054 404854
rect 296434 387174 297054 404618
rect 296434 386938 296466 387174
rect 296702 386938 296786 387174
rect 297022 386938 297054 387174
rect 296434 386854 297054 386938
rect 296434 386618 296466 386854
rect 296702 386618 296786 386854
rect 297022 386618 297054 386854
rect 296434 369174 297054 386618
rect 296434 368938 296466 369174
rect 296702 368938 296786 369174
rect 297022 368938 297054 369174
rect 296434 368854 297054 368938
rect 296434 368618 296466 368854
rect 296702 368618 296786 368854
rect 297022 368618 297054 368854
rect 296434 351174 297054 368618
rect 296434 350938 296466 351174
rect 296702 350938 296786 351174
rect 297022 350938 297054 351174
rect 296434 350854 297054 350938
rect 296434 350618 296466 350854
rect 296702 350618 296786 350854
rect 297022 350618 297054 350854
rect 296434 333174 297054 350618
rect 296434 332938 296466 333174
rect 296702 332938 296786 333174
rect 297022 332938 297054 333174
rect 296434 332854 297054 332938
rect 296434 332618 296466 332854
rect 296702 332618 296786 332854
rect 297022 332618 297054 332854
rect 296434 315174 297054 332618
rect 296434 314938 296466 315174
rect 296702 314938 296786 315174
rect 297022 314938 297054 315174
rect 296434 314854 297054 314938
rect 296434 314618 296466 314854
rect 296702 314618 296786 314854
rect 297022 314618 297054 314854
rect 296434 297174 297054 314618
rect 296434 296938 296466 297174
rect 296702 296938 296786 297174
rect 297022 296938 297054 297174
rect 296434 296854 297054 296938
rect 296434 296618 296466 296854
rect 296702 296618 296786 296854
rect 297022 296618 297054 296854
rect 296434 279174 297054 296618
rect 296434 278938 296466 279174
rect 296702 278938 296786 279174
rect 297022 278938 297054 279174
rect 296434 278854 297054 278938
rect 296434 278618 296466 278854
rect 296702 278618 296786 278854
rect 297022 278618 297054 278854
rect 296434 261174 297054 278618
rect 296434 260938 296466 261174
rect 296702 260938 296786 261174
rect 297022 260938 297054 261174
rect 296434 260854 297054 260938
rect 296434 260618 296466 260854
rect 296702 260618 296786 260854
rect 297022 260618 297054 260854
rect 296434 243174 297054 260618
rect 296434 242938 296466 243174
rect 296702 242938 296786 243174
rect 297022 242938 297054 243174
rect 296434 242854 297054 242938
rect 296434 242618 296466 242854
rect 296702 242618 296786 242854
rect 297022 242618 297054 242854
rect 296434 225174 297054 242618
rect 296434 224938 296466 225174
rect 296702 224938 296786 225174
rect 297022 224938 297054 225174
rect 296434 224854 297054 224938
rect 296434 224618 296466 224854
rect 296702 224618 296786 224854
rect 297022 224618 297054 224854
rect 296434 207174 297054 224618
rect 296434 206938 296466 207174
rect 296702 206938 296786 207174
rect 297022 206938 297054 207174
rect 296434 206854 297054 206938
rect 296434 206618 296466 206854
rect 296702 206618 296786 206854
rect 297022 206618 297054 206854
rect 296434 189174 297054 206618
rect 296434 188938 296466 189174
rect 296702 188938 296786 189174
rect 297022 188938 297054 189174
rect 296434 188854 297054 188938
rect 296434 188618 296466 188854
rect 296702 188618 296786 188854
rect 297022 188618 297054 188854
rect 296434 171174 297054 188618
rect 296434 170938 296466 171174
rect 296702 170938 296786 171174
rect 297022 170938 297054 171174
rect 296434 170854 297054 170938
rect 296434 170618 296466 170854
rect 296702 170618 296786 170854
rect 297022 170618 297054 170854
rect 296434 153174 297054 170618
rect 296434 152938 296466 153174
rect 296702 152938 296786 153174
rect 297022 152938 297054 153174
rect 296434 152854 297054 152938
rect 296434 152618 296466 152854
rect 296702 152618 296786 152854
rect 297022 152618 297054 152854
rect 296434 135174 297054 152618
rect 296434 134938 296466 135174
rect 296702 134938 296786 135174
rect 297022 134938 297054 135174
rect 296434 134854 297054 134938
rect 296434 134618 296466 134854
rect 296702 134618 296786 134854
rect 297022 134618 297054 134854
rect 296434 117174 297054 134618
rect 296434 116938 296466 117174
rect 296702 116938 296786 117174
rect 297022 116938 297054 117174
rect 296434 116854 297054 116938
rect 296434 116618 296466 116854
rect 296702 116618 296786 116854
rect 297022 116618 297054 116854
rect 296434 99174 297054 116618
rect 296434 98938 296466 99174
rect 296702 98938 296786 99174
rect 297022 98938 297054 99174
rect 296434 98854 297054 98938
rect 296434 98618 296466 98854
rect 296702 98618 296786 98854
rect 297022 98618 297054 98854
rect 296434 81174 297054 98618
rect 296434 80938 296466 81174
rect 296702 80938 296786 81174
rect 297022 80938 297054 81174
rect 296434 80854 297054 80938
rect 296434 80618 296466 80854
rect 296702 80618 296786 80854
rect 297022 80618 297054 80854
rect 296434 63174 297054 80618
rect 296434 62938 296466 63174
rect 296702 62938 296786 63174
rect 297022 62938 297054 63174
rect 296434 62854 297054 62938
rect 296434 62618 296466 62854
rect 296702 62618 296786 62854
rect 297022 62618 297054 62854
rect 296434 45174 297054 62618
rect 296434 44938 296466 45174
rect 296702 44938 296786 45174
rect 297022 44938 297054 45174
rect 296434 44854 297054 44938
rect 296434 44618 296466 44854
rect 296702 44618 296786 44854
rect 297022 44618 297054 44854
rect 296434 27174 297054 44618
rect 296434 26938 296466 27174
rect 296702 26938 296786 27174
rect 297022 26938 297054 27174
rect 296434 26854 297054 26938
rect 296434 26618 296466 26854
rect 296702 26618 296786 26854
rect 297022 26618 297054 26854
rect 296434 9174 297054 26618
rect 296434 8938 296466 9174
rect 296702 8938 296786 9174
rect 297022 8938 297054 9174
rect 296434 8854 297054 8938
rect 296434 8618 296466 8854
rect 296702 8618 296786 8854
rect 297022 8618 297054 8854
rect 296434 -1816 297054 8618
rect 296434 -2052 296466 -1816
rect 296702 -2052 296786 -1816
rect 297022 -2052 297054 -1816
rect 296434 -2136 297054 -2052
rect 296434 -2372 296466 -2136
rect 296702 -2372 296786 -2136
rect 297022 -2372 297054 -2136
rect 296434 -4324 297054 -2372
rect 300154 463012 300774 464004
rect 300154 462776 300186 463012
rect 300422 462776 300506 463012
rect 300742 462776 300774 463012
rect 300154 462692 300774 462776
rect 300154 462456 300186 462692
rect 300422 462456 300506 462692
rect 300742 462456 300774 462692
rect 300154 444894 300774 462456
rect 300154 444658 300186 444894
rect 300422 444658 300506 444894
rect 300742 444658 300774 444894
rect 300154 444574 300774 444658
rect 300154 444338 300186 444574
rect 300422 444338 300506 444574
rect 300742 444338 300774 444574
rect 300154 426894 300774 444338
rect 300154 426658 300186 426894
rect 300422 426658 300506 426894
rect 300742 426658 300774 426894
rect 300154 426574 300774 426658
rect 300154 426338 300186 426574
rect 300422 426338 300506 426574
rect 300742 426338 300774 426574
rect 300154 408894 300774 426338
rect 300154 408658 300186 408894
rect 300422 408658 300506 408894
rect 300742 408658 300774 408894
rect 300154 408574 300774 408658
rect 300154 408338 300186 408574
rect 300422 408338 300506 408574
rect 300742 408338 300774 408574
rect 300154 390894 300774 408338
rect 300154 390658 300186 390894
rect 300422 390658 300506 390894
rect 300742 390658 300774 390894
rect 300154 390574 300774 390658
rect 300154 390338 300186 390574
rect 300422 390338 300506 390574
rect 300742 390338 300774 390574
rect 300154 372894 300774 390338
rect 300154 372658 300186 372894
rect 300422 372658 300506 372894
rect 300742 372658 300774 372894
rect 300154 372574 300774 372658
rect 300154 372338 300186 372574
rect 300422 372338 300506 372574
rect 300742 372338 300774 372574
rect 300154 354894 300774 372338
rect 300154 354658 300186 354894
rect 300422 354658 300506 354894
rect 300742 354658 300774 354894
rect 300154 354574 300774 354658
rect 300154 354338 300186 354574
rect 300422 354338 300506 354574
rect 300742 354338 300774 354574
rect 300154 336894 300774 354338
rect 300154 336658 300186 336894
rect 300422 336658 300506 336894
rect 300742 336658 300774 336894
rect 300154 336574 300774 336658
rect 300154 336338 300186 336574
rect 300422 336338 300506 336574
rect 300742 336338 300774 336574
rect 300154 318894 300774 336338
rect 300154 318658 300186 318894
rect 300422 318658 300506 318894
rect 300742 318658 300774 318894
rect 300154 318574 300774 318658
rect 300154 318338 300186 318574
rect 300422 318338 300506 318574
rect 300742 318338 300774 318574
rect 300154 300894 300774 318338
rect 300154 300658 300186 300894
rect 300422 300658 300506 300894
rect 300742 300658 300774 300894
rect 300154 300574 300774 300658
rect 300154 300338 300186 300574
rect 300422 300338 300506 300574
rect 300742 300338 300774 300574
rect 300154 282894 300774 300338
rect 300154 282658 300186 282894
rect 300422 282658 300506 282894
rect 300742 282658 300774 282894
rect 300154 282574 300774 282658
rect 300154 282338 300186 282574
rect 300422 282338 300506 282574
rect 300742 282338 300774 282574
rect 300154 264894 300774 282338
rect 300154 264658 300186 264894
rect 300422 264658 300506 264894
rect 300742 264658 300774 264894
rect 300154 264574 300774 264658
rect 300154 264338 300186 264574
rect 300422 264338 300506 264574
rect 300742 264338 300774 264574
rect 300154 246894 300774 264338
rect 300154 246658 300186 246894
rect 300422 246658 300506 246894
rect 300742 246658 300774 246894
rect 300154 246574 300774 246658
rect 300154 246338 300186 246574
rect 300422 246338 300506 246574
rect 300742 246338 300774 246574
rect 300154 228894 300774 246338
rect 300154 228658 300186 228894
rect 300422 228658 300506 228894
rect 300742 228658 300774 228894
rect 300154 228574 300774 228658
rect 300154 228338 300186 228574
rect 300422 228338 300506 228574
rect 300742 228338 300774 228574
rect 300154 210894 300774 228338
rect 300154 210658 300186 210894
rect 300422 210658 300506 210894
rect 300742 210658 300774 210894
rect 300154 210574 300774 210658
rect 300154 210338 300186 210574
rect 300422 210338 300506 210574
rect 300742 210338 300774 210574
rect 300154 192894 300774 210338
rect 300154 192658 300186 192894
rect 300422 192658 300506 192894
rect 300742 192658 300774 192894
rect 300154 192574 300774 192658
rect 300154 192338 300186 192574
rect 300422 192338 300506 192574
rect 300742 192338 300774 192574
rect 300154 174894 300774 192338
rect 300154 174658 300186 174894
rect 300422 174658 300506 174894
rect 300742 174658 300774 174894
rect 300154 174574 300774 174658
rect 300154 174338 300186 174574
rect 300422 174338 300506 174574
rect 300742 174338 300774 174574
rect 300154 156894 300774 174338
rect 300154 156658 300186 156894
rect 300422 156658 300506 156894
rect 300742 156658 300774 156894
rect 300154 156574 300774 156658
rect 300154 156338 300186 156574
rect 300422 156338 300506 156574
rect 300742 156338 300774 156574
rect 300154 138894 300774 156338
rect 300154 138658 300186 138894
rect 300422 138658 300506 138894
rect 300742 138658 300774 138894
rect 300154 138574 300774 138658
rect 300154 138338 300186 138574
rect 300422 138338 300506 138574
rect 300742 138338 300774 138574
rect 300154 120894 300774 138338
rect 300154 120658 300186 120894
rect 300422 120658 300506 120894
rect 300742 120658 300774 120894
rect 300154 120574 300774 120658
rect 300154 120338 300186 120574
rect 300422 120338 300506 120574
rect 300742 120338 300774 120574
rect 300154 102894 300774 120338
rect 300154 102658 300186 102894
rect 300422 102658 300506 102894
rect 300742 102658 300774 102894
rect 300154 102574 300774 102658
rect 300154 102338 300186 102574
rect 300422 102338 300506 102574
rect 300742 102338 300774 102574
rect 300154 84894 300774 102338
rect 300154 84658 300186 84894
rect 300422 84658 300506 84894
rect 300742 84658 300774 84894
rect 300154 84574 300774 84658
rect 300154 84338 300186 84574
rect 300422 84338 300506 84574
rect 300742 84338 300774 84574
rect 300154 66894 300774 84338
rect 300154 66658 300186 66894
rect 300422 66658 300506 66894
rect 300742 66658 300774 66894
rect 300154 66574 300774 66658
rect 300154 66338 300186 66574
rect 300422 66338 300506 66574
rect 300742 66338 300774 66574
rect 300154 48894 300774 66338
rect 300154 48658 300186 48894
rect 300422 48658 300506 48894
rect 300742 48658 300774 48894
rect 300154 48574 300774 48658
rect 300154 48338 300186 48574
rect 300422 48338 300506 48574
rect 300742 48338 300774 48574
rect 300154 30894 300774 48338
rect 300154 30658 300186 30894
rect 300422 30658 300506 30894
rect 300742 30658 300774 30894
rect 300154 30574 300774 30658
rect 300154 30338 300186 30574
rect 300422 30338 300506 30574
rect 300742 30338 300774 30574
rect 300154 12894 300774 30338
rect 300154 12658 300186 12894
rect 300422 12658 300506 12894
rect 300742 12658 300774 12894
rect 300154 12574 300774 12658
rect 300154 12338 300186 12574
rect 300422 12338 300506 12574
rect 300742 12338 300774 12574
rect 300154 -2776 300774 12338
rect 300154 -3012 300186 -2776
rect 300422 -3012 300506 -2776
rect 300742 -3012 300774 -2776
rect 300154 -3096 300774 -3012
rect 300154 -3332 300186 -3096
rect 300422 -3332 300506 -3096
rect 300742 -3332 300774 -3096
rect 300154 -4324 300774 -3332
rect 303874 463972 304494 464004
rect 303874 463736 303906 463972
rect 304142 463736 304226 463972
rect 304462 463736 304494 463972
rect 303874 463652 304494 463736
rect 303874 463416 303906 463652
rect 304142 463416 304226 463652
rect 304462 463416 304494 463652
rect 303874 448614 304494 463416
rect 303874 448378 303906 448614
rect 304142 448378 304226 448614
rect 304462 448378 304494 448614
rect 303874 448294 304494 448378
rect 303874 448058 303906 448294
rect 304142 448058 304226 448294
rect 304462 448058 304494 448294
rect 303874 430614 304494 448058
rect 303874 430378 303906 430614
rect 304142 430378 304226 430614
rect 304462 430378 304494 430614
rect 303874 430294 304494 430378
rect 303874 430058 303906 430294
rect 304142 430058 304226 430294
rect 304462 430058 304494 430294
rect 303874 412614 304494 430058
rect 303874 412378 303906 412614
rect 304142 412378 304226 412614
rect 304462 412378 304494 412614
rect 303874 412294 304494 412378
rect 303874 412058 303906 412294
rect 304142 412058 304226 412294
rect 304462 412058 304494 412294
rect 303874 394614 304494 412058
rect 303874 394378 303906 394614
rect 304142 394378 304226 394614
rect 304462 394378 304494 394614
rect 303874 394294 304494 394378
rect 303874 394058 303906 394294
rect 304142 394058 304226 394294
rect 304462 394058 304494 394294
rect 303874 376614 304494 394058
rect 303874 376378 303906 376614
rect 304142 376378 304226 376614
rect 304462 376378 304494 376614
rect 303874 376294 304494 376378
rect 303874 376058 303906 376294
rect 304142 376058 304226 376294
rect 304462 376058 304494 376294
rect 303874 358614 304494 376058
rect 303874 358378 303906 358614
rect 304142 358378 304226 358614
rect 304462 358378 304494 358614
rect 303874 358294 304494 358378
rect 303874 358058 303906 358294
rect 304142 358058 304226 358294
rect 304462 358058 304494 358294
rect 303874 340614 304494 358058
rect 303874 340378 303906 340614
rect 304142 340378 304226 340614
rect 304462 340378 304494 340614
rect 303874 340294 304494 340378
rect 303874 340058 303906 340294
rect 304142 340058 304226 340294
rect 304462 340058 304494 340294
rect 303874 322614 304494 340058
rect 303874 322378 303906 322614
rect 304142 322378 304226 322614
rect 304462 322378 304494 322614
rect 303874 322294 304494 322378
rect 303874 322058 303906 322294
rect 304142 322058 304226 322294
rect 304462 322058 304494 322294
rect 303874 304614 304494 322058
rect 303874 304378 303906 304614
rect 304142 304378 304226 304614
rect 304462 304378 304494 304614
rect 303874 304294 304494 304378
rect 303874 304058 303906 304294
rect 304142 304058 304226 304294
rect 304462 304058 304494 304294
rect 303874 286614 304494 304058
rect 303874 286378 303906 286614
rect 304142 286378 304226 286614
rect 304462 286378 304494 286614
rect 303874 286294 304494 286378
rect 303874 286058 303906 286294
rect 304142 286058 304226 286294
rect 304462 286058 304494 286294
rect 303874 268614 304494 286058
rect 303874 268378 303906 268614
rect 304142 268378 304226 268614
rect 304462 268378 304494 268614
rect 303874 268294 304494 268378
rect 303874 268058 303906 268294
rect 304142 268058 304226 268294
rect 304462 268058 304494 268294
rect 303874 250614 304494 268058
rect 303874 250378 303906 250614
rect 304142 250378 304226 250614
rect 304462 250378 304494 250614
rect 303874 250294 304494 250378
rect 303874 250058 303906 250294
rect 304142 250058 304226 250294
rect 304462 250058 304494 250294
rect 303874 232614 304494 250058
rect 303874 232378 303906 232614
rect 304142 232378 304226 232614
rect 304462 232378 304494 232614
rect 303874 232294 304494 232378
rect 303874 232058 303906 232294
rect 304142 232058 304226 232294
rect 304462 232058 304494 232294
rect 303874 214614 304494 232058
rect 303874 214378 303906 214614
rect 304142 214378 304226 214614
rect 304462 214378 304494 214614
rect 303874 214294 304494 214378
rect 303874 214058 303906 214294
rect 304142 214058 304226 214294
rect 304462 214058 304494 214294
rect 303874 196614 304494 214058
rect 303874 196378 303906 196614
rect 304142 196378 304226 196614
rect 304462 196378 304494 196614
rect 303874 196294 304494 196378
rect 303874 196058 303906 196294
rect 304142 196058 304226 196294
rect 304462 196058 304494 196294
rect 303874 178614 304494 196058
rect 303874 178378 303906 178614
rect 304142 178378 304226 178614
rect 304462 178378 304494 178614
rect 303874 178294 304494 178378
rect 303874 178058 303906 178294
rect 304142 178058 304226 178294
rect 304462 178058 304494 178294
rect 303874 160614 304494 178058
rect 303874 160378 303906 160614
rect 304142 160378 304226 160614
rect 304462 160378 304494 160614
rect 303874 160294 304494 160378
rect 303874 160058 303906 160294
rect 304142 160058 304226 160294
rect 304462 160058 304494 160294
rect 303874 142614 304494 160058
rect 303874 142378 303906 142614
rect 304142 142378 304226 142614
rect 304462 142378 304494 142614
rect 303874 142294 304494 142378
rect 303874 142058 303906 142294
rect 304142 142058 304226 142294
rect 304462 142058 304494 142294
rect 303874 124614 304494 142058
rect 303874 124378 303906 124614
rect 304142 124378 304226 124614
rect 304462 124378 304494 124614
rect 303874 124294 304494 124378
rect 303874 124058 303906 124294
rect 304142 124058 304226 124294
rect 304462 124058 304494 124294
rect 303874 106614 304494 124058
rect 303874 106378 303906 106614
rect 304142 106378 304226 106614
rect 304462 106378 304494 106614
rect 303874 106294 304494 106378
rect 303874 106058 303906 106294
rect 304142 106058 304226 106294
rect 304462 106058 304494 106294
rect 303874 88614 304494 106058
rect 303874 88378 303906 88614
rect 304142 88378 304226 88614
rect 304462 88378 304494 88614
rect 303874 88294 304494 88378
rect 303874 88058 303906 88294
rect 304142 88058 304226 88294
rect 304462 88058 304494 88294
rect 303874 70614 304494 88058
rect 303874 70378 303906 70614
rect 304142 70378 304226 70614
rect 304462 70378 304494 70614
rect 303874 70294 304494 70378
rect 303874 70058 303906 70294
rect 304142 70058 304226 70294
rect 304462 70058 304494 70294
rect 303874 52614 304494 70058
rect 303874 52378 303906 52614
rect 304142 52378 304226 52614
rect 304462 52378 304494 52614
rect 303874 52294 304494 52378
rect 303874 52058 303906 52294
rect 304142 52058 304226 52294
rect 304462 52058 304494 52294
rect 303874 34614 304494 52058
rect 303874 34378 303906 34614
rect 304142 34378 304226 34614
rect 304462 34378 304494 34614
rect 303874 34294 304494 34378
rect 303874 34058 303906 34294
rect 304142 34058 304226 34294
rect 304462 34058 304494 34294
rect 303874 16614 304494 34058
rect 303874 16378 303906 16614
rect 304142 16378 304226 16614
rect 304462 16378 304494 16614
rect 303874 16294 304494 16378
rect 303874 16058 303906 16294
rect 304142 16058 304226 16294
rect 304462 16058 304494 16294
rect 303874 -3736 304494 16058
rect 303874 -3972 303906 -3736
rect 304142 -3972 304226 -3736
rect 304462 -3972 304494 -3736
rect 303874 -4056 304494 -3972
rect 303874 -4292 303906 -4056
rect 304142 -4292 304226 -4056
rect 304462 -4292 304494 -4056
rect 303874 -4324 304494 -4292
rect 310714 461092 311334 464004
rect 310714 460856 310746 461092
rect 310982 460856 311066 461092
rect 311302 460856 311334 461092
rect 310714 460772 311334 460856
rect 310714 460536 310746 460772
rect 310982 460536 311066 460772
rect 311302 460536 311334 460772
rect 310714 455454 311334 460536
rect 310714 455218 310746 455454
rect 310982 455218 311066 455454
rect 311302 455218 311334 455454
rect 310714 455134 311334 455218
rect 310714 454898 310746 455134
rect 310982 454898 311066 455134
rect 311302 454898 311334 455134
rect 310714 437454 311334 454898
rect 310714 437218 310746 437454
rect 310982 437218 311066 437454
rect 311302 437218 311334 437454
rect 310714 437134 311334 437218
rect 310714 436898 310746 437134
rect 310982 436898 311066 437134
rect 311302 436898 311334 437134
rect 310714 419454 311334 436898
rect 310714 419218 310746 419454
rect 310982 419218 311066 419454
rect 311302 419218 311334 419454
rect 310714 419134 311334 419218
rect 310714 418898 310746 419134
rect 310982 418898 311066 419134
rect 311302 418898 311334 419134
rect 310714 401454 311334 418898
rect 310714 401218 310746 401454
rect 310982 401218 311066 401454
rect 311302 401218 311334 401454
rect 310714 401134 311334 401218
rect 310714 400898 310746 401134
rect 310982 400898 311066 401134
rect 311302 400898 311334 401134
rect 310714 383454 311334 400898
rect 310714 383218 310746 383454
rect 310982 383218 311066 383454
rect 311302 383218 311334 383454
rect 310714 383134 311334 383218
rect 310714 382898 310746 383134
rect 310982 382898 311066 383134
rect 311302 382898 311334 383134
rect 310714 365454 311334 382898
rect 310714 365218 310746 365454
rect 310982 365218 311066 365454
rect 311302 365218 311334 365454
rect 310714 365134 311334 365218
rect 310714 364898 310746 365134
rect 310982 364898 311066 365134
rect 311302 364898 311334 365134
rect 310714 347454 311334 364898
rect 310714 347218 310746 347454
rect 310982 347218 311066 347454
rect 311302 347218 311334 347454
rect 310714 347134 311334 347218
rect 310714 346898 310746 347134
rect 310982 346898 311066 347134
rect 311302 346898 311334 347134
rect 310714 329454 311334 346898
rect 310714 329218 310746 329454
rect 310982 329218 311066 329454
rect 311302 329218 311334 329454
rect 310714 329134 311334 329218
rect 310714 328898 310746 329134
rect 310982 328898 311066 329134
rect 311302 328898 311334 329134
rect 310714 311454 311334 328898
rect 310714 311218 310746 311454
rect 310982 311218 311066 311454
rect 311302 311218 311334 311454
rect 310714 311134 311334 311218
rect 310714 310898 310746 311134
rect 310982 310898 311066 311134
rect 311302 310898 311334 311134
rect 310714 293454 311334 310898
rect 310714 293218 310746 293454
rect 310982 293218 311066 293454
rect 311302 293218 311334 293454
rect 310714 293134 311334 293218
rect 310714 292898 310746 293134
rect 310982 292898 311066 293134
rect 311302 292898 311334 293134
rect 310714 275454 311334 292898
rect 310714 275218 310746 275454
rect 310982 275218 311066 275454
rect 311302 275218 311334 275454
rect 310714 275134 311334 275218
rect 310714 274898 310746 275134
rect 310982 274898 311066 275134
rect 311302 274898 311334 275134
rect 310714 257454 311334 274898
rect 310714 257218 310746 257454
rect 310982 257218 311066 257454
rect 311302 257218 311334 257454
rect 310714 257134 311334 257218
rect 310714 256898 310746 257134
rect 310982 256898 311066 257134
rect 311302 256898 311334 257134
rect 310714 239454 311334 256898
rect 310714 239218 310746 239454
rect 310982 239218 311066 239454
rect 311302 239218 311334 239454
rect 310714 239134 311334 239218
rect 310714 238898 310746 239134
rect 310982 238898 311066 239134
rect 311302 238898 311334 239134
rect 310714 221454 311334 238898
rect 310714 221218 310746 221454
rect 310982 221218 311066 221454
rect 311302 221218 311334 221454
rect 310714 221134 311334 221218
rect 310714 220898 310746 221134
rect 310982 220898 311066 221134
rect 311302 220898 311334 221134
rect 310714 203454 311334 220898
rect 310714 203218 310746 203454
rect 310982 203218 311066 203454
rect 311302 203218 311334 203454
rect 310714 203134 311334 203218
rect 310714 202898 310746 203134
rect 310982 202898 311066 203134
rect 311302 202898 311334 203134
rect 310714 185454 311334 202898
rect 310714 185218 310746 185454
rect 310982 185218 311066 185454
rect 311302 185218 311334 185454
rect 310714 185134 311334 185218
rect 310714 184898 310746 185134
rect 310982 184898 311066 185134
rect 311302 184898 311334 185134
rect 310714 167454 311334 184898
rect 310714 167218 310746 167454
rect 310982 167218 311066 167454
rect 311302 167218 311334 167454
rect 310714 167134 311334 167218
rect 310714 166898 310746 167134
rect 310982 166898 311066 167134
rect 311302 166898 311334 167134
rect 310714 149454 311334 166898
rect 310714 149218 310746 149454
rect 310982 149218 311066 149454
rect 311302 149218 311334 149454
rect 310714 149134 311334 149218
rect 310714 148898 310746 149134
rect 310982 148898 311066 149134
rect 311302 148898 311334 149134
rect 310714 131454 311334 148898
rect 310714 131218 310746 131454
rect 310982 131218 311066 131454
rect 311302 131218 311334 131454
rect 310714 131134 311334 131218
rect 310714 130898 310746 131134
rect 310982 130898 311066 131134
rect 311302 130898 311334 131134
rect 310714 113454 311334 130898
rect 310714 113218 310746 113454
rect 310982 113218 311066 113454
rect 311302 113218 311334 113454
rect 310714 113134 311334 113218
rect 310714 112898 310746 113134
rect 310982 112898 311066 113134
rect 311302 112898 311334 113134
rect 310714 95454 311334 112898
rect 310714 95218 310746 95454
rect 310982 95218 311066 95454
rect 311302 95218 311334 95454
rect 310714 95134 311334 95218
rect 310714 94898 310746 95134
rect 310982 94898 311066 95134
rect 311302 94898 311334 95134
rect 310714 77454 311334 94898
rect 310714 77218 310746 77454
rect 310982 77218 311066 77454
rect 311302 77218 311334 77454
rect 310714 77134 311334 77218
rect 310714 76898 310746 77134
rect 310982 76898 311066 77134
rect 311302 76898 311334 77134
rect 310714 59454 311334 76898
rect 310714 59218 310746 59454
rect 310982 59218 311066 59454
rect 311302 59218 311334 59454
rect 310714 59134 311334 59218
rect 310714 58898 310746 59134
rect 310982 58898 311066 59134
rect 311302 58898 311334 59134
rect 310714 41454 311334 58898
rect 310714 41218 310746 41454
rect 310982 41218 311066 41454
rect 311302 41218 311334 41454
rect 310714 41134 311334 41218
rect 310714 40898 310746 41134
rect 310982 40898 311066 41134
rect 311302 40898 311334 41134
rect 310714 23454 311334 40898
rect 310714 23218 310746 23454
rect 310982 23218 311066 23454
rect 311302 23218 311334 23454
rect 310714 23134 311334 23218
rect 310714 22898 310746 23134
rect 310982 22898 311066 23134
rect 311302 22898 311334 23134
rect 310714 5454 311334 22898
rect 310714 5218 310746 5454
rect 310982 5218 311066 5454
rect 311302 5218 311334 5454
rect 310714 5134 311334 5218
rect 310714 4898 310746 5134
rect 310982 4898 311066 5134
rect 311302 4898 311334 5134
rect 310714 -856 311334 4898
rect 310714 -1092 310746 -856
rect 310982 -1092 311066 -856
rect 311302 -1092 311334 -856
rect 310714 -1176 311334 -1092
rect 310714 -1412 310746 -1176
rect 310982 -1412 311066 -1176
rect 311302 -1412 311334 -1176
rect 310714 -4324 311334 -1412
rect 314434 462052 315054 464004
rect 314434 461816 314466 462052
rect 314702 461816 314786 462052
rect 315022 461816 315054 462052
rect 314434 461732 315054 461816
rect 314434 461496 314466 461732
rect 314702 461496 314786 461732
rect 315022 461496 315054 461732
rect 314434 441174 315054 461496
rect 314434 440938 314466 441174
rect 314702 440938 314786 441174
rect 315022 440938 315054 441174
rect 314434 440854 315054 440938
rect 314434 440618 314466 440854
rect 314702 440618 314786 440854
rect 315022 440618 315054 440854
rect 314434 423174 315054 440618
rect 314434 422938 314466 423174
rect 314702 422938 314786 423174
rect 315022 422938 315054 423174
rect 314434 422854 315054 422938
rect 314434 422618 314466 422854
rect 314702 422618 314786 422854
rect 315022 422618 315054 422854
rect 314434 405174 315054 422618
rect 314434 404938 314466 405174
rect 314702 404938 314786 405174
rect 315022 404938 315054 405174
rect 314434 404854 315054 404938
rect 314434 404618 314466 404854
rect 314702 404618 314786 404854
rect 315022 404618 315054 404854
rect 314434 387174 315054 404618
rect 314434 386938 314466 387174
rect 314702 386938 314786 387174
rect 315022 386938 315054 387174
rect 314434 386854 315054 386938
rect 314434 386618 314466 386854
rect 314702 386618 314786 386854
rect 315022 386618 315054 386854
rect 314434 369174 315054 386618
rect 314434 368938 314466 369174
rect 314702 368938 314786 369174
rect 315022 368938 315054 369174
rect 314434 368854 315054 368938
rect 314434 368618 314466 368854
rect 314702 368618 314786 368854
rect 315022 368618 315054 368854
rect 314434 351174 315054 368618
rect 314434 350938 314466 351174
rect 314702 350938 314786 351174
rect 315022 350938 315054 351174
rect 314434 350854 315054 350938
rect 314434 350618 314466 350854
rect 314702 350618 314786 350854
rect 315022 350618 315054 350854
rect 314434 333174 315054 350618
rect 314434 332938 314466 333174
rect 314702 332938 314786 333174
rect 315022 332938 315054 333174
rect 314434 332854 315054 332938
rect 314434 332618 314466 332854
rect 314702 332618 314786 332854
rect 315022 332618 315054 332854
rect 314434 315174 315054 332618
rect 314434 314938 314466 315174
rect 314702 314938 314786 315174
rect 315022 314938 315054 315174
rect 314434 314854 315054 314938
rect 314434 314618 314466 314854
rect 314702 314618 314786 314854
rect 315022 314618 315054 314854
rect 314434 297174 315054 314618
rect 314434 296938 314466 297174
rect 314702 296938 314786 297174
rect 315022 296938 315054 297174
rect 314434 296854 315054 296938
rect 314434 296618 314466 296854
rect 314702 296618 314786 296854
rect 315022 296618 315054 296854
rect 314434 279174 315054 296618
rect 314434 278938 314466 279174
rect 314702 278938 314786 279174
rect 315022 278938 315054 279174
rect 314434 278854 315054 278938
rect 314434 278618 314466 278854
rect 314702 278618 314786 278854
rect 315022 278618 315054 278854
rect 314434 261174 315054 278618
rect 314434 260938 314466 261174
rect 314702 260938 314786 261174
rect 315022 260938 315054 261174
rect 314434 260854 315054 260938
rect 314434 260618 314466 260854
rect 314702 260618 314786 260854
rect 315022 260618 315054 260854
rect 314434 243174 315054 260618
rect 314434 242938 314466 243174
rect 314702 242938 314786 243174
rect 315022 242938 315054 243174
rect 314434 242854 315054 242938
rect 314434 242618 314466 242854
rect 314702 242618 314786 242854
rect 315022 242618 315054 242854
rect 314434 225174 315054 242618
rect 314434 224938 314466 225174
rect 314702 224938 314786 225174
rect 315022 224938 315054 225174
rect 314434 224854 315054 224938
rect 314434 224618 314466 224854
rect 314702 224618 314786 224854
rect 315022 224618 315054 224854
rect 314434 207174 315054 224618
rect 314434 206938 314466 207174
rect 314702 206938 314786 207174
rect 315022 206938 315054 207174
rect 314434 206854 315054 206938
rect 314434 206618 314466 206854
rect 314702 206618 314786 206854
rect 315022 206618 315054 206854
rect 314434 189174 315054 206618
rect 314434 188938 314466 189174
rect 314702 188938 314786 189174
rect 315022 188938 315054 189174
rect 314434 188854 315054 188938
rect 314434 188618 314466 188854
rect 314702 188618 314786 188854
rect 315022 188618 315054 188854
rect 314434 171174 315054 188618
rect 314434 170938 314466 171174
rect 314702 170938 314786 171174
rect 315022 170938 315054 171174
rect 314434 170854 315054 170938
rect 314434 170618 314466 170854
rect 314702 170618 314786 170854
rect 315022 170618 315054 170854
rect 314434 153174 315054 170618
rect 314434 152938 314466 153174
rect 314702 152938 314786 153174
rect 315022 152938 315054 153174
rect 314434 152854 315054 152938
rect 314434 152618 314466 152854
rect 314702 152618 314786 152854
rect 315022 152618 315054 152854
rect 314434 135174 315054 152618
rect 314434 134938 314466 135174
rect 314702 134938 314786 135174
rect 315022 134938 315054 135174
rect 314434 134854 315054 134938
rect 314434 134618 314466 134854
rect 314702 134618 314786 134854
rect 315022 134618 315054 134854
rect 314434 117174 315054 134618
rect 314434 116938 314466 117174
rect 314702 116938 314786 117174
rect 315022 116938 315054 117174
rect 314434 116854 315054 116938
rect 314434 116618 314466 116854
rect 314702 116618 314786 116854
rect 315022 116618 315054 116854
rect 314434 99174 315054 116618
rect 314434 98938 314466 99174
rect 314702 98938 314786 99174
rect 315022 98938 315054 99174
rect 314434 98854 315054 98938
rect 314434 98618 314466 98854
rect 314702 98618 314786 98854
rect 315022 98618 315054 98854
rect 314434 81174 315054 98618
rect 314434 80938 314466 81174
rect 314702 80938 314786 81174
rect 315022 80938 315054 81174
rect 314434 80854 315054 80938
rect 314434 80618 314466 80854
rect 314702 80618 314786 80854
rect 315022 80618 315054 80854
rect 314434 63174 315054 80618
rect 314434 62938 314466 63174
rect 314702 62938 314786 63174
rect 315022 62938 315054 63174
rect 314434 62854 315054 62938
rect 314434 62618 314466 62854
rect 314702 62618 314786 62854
rect 315022 62618 315054 62854
rect 314434 45174 315054 62618
rect 314434 44938 314466 45174
rect 314702 44938 314786 45174
rect 315022 44938 315054 45174
rect 314434 44854 315054 44938
rect 314434 44618 314466 44854
rect 314702 44618 314786 44854
rect 315022 44618 315054 44854
rect 314434 27174 315054 44618
rect 314434 26938 314466 27174
rect 314702 26938 314786 27174
rect 315022 26938 315054 27174
rect 314434 26854 315054 26938
rect 314434 26618 314466 26854
rect 314702 26618 314786 26854
rect 315022 26618 315054 26854
rect 314434 9174 315054 26618
rect 314434 8938 314466 9174
rect 314702 8938 314786 9174
rect 315022 8938 315054 9174
rect 314434 8854 315054 8938
rect 314434 8618 314466 8854
rect 314702 8618 314786 8854
rect 315022 8618 315054 8854
rect 314434 -1816 315054 8618
rect 314434 -2052 314466 -1816
rect 314702 -2052 314786 -1816
rect 315022 -2052 315054 -1816
rect 314434 -2136 315054 -2052
rect 314434 -2372 314466 -2136
rect 314702 -2372 314786 -2136
rect 315022 -2372 315054 -2136
rect 314434 -4324 315054 -2372
rect 318154 463012 318774 464004
rect 318154 462776 318186 463012
rect 318422 462776 318506 463012
rect 318742 462776 318774 463012
rect 318154 462692 318774 462776
rect 318154 462456 318186 462692
rect 318422 462456 318506 462692
rect 318742 462456 318774 462692
rect 318154 444894 318774 462456
rect 318154 444658 318186 444894
rect 318422 444658 318506 444894
rect 318742 444658 318774 444894
rect 318154 444574 318774 444658
rect 318154 444338 318186 444574
rect 318422 444338 318506 444574
rect 318742 444338 318774 444574
rect 318154 426894 318774 444338
rect 318154 426658 318186 426894
rect 318422 426658 318506 426894
rect 318742 426658 318774 426894
rect 318154 426574 318774 426658
rect 318154 426338 318186 426574
rect 318422 426338 318506 426574
rect 318742 426338 318774 426574
rect 318154 408894 318774 426338
rect 318154 408658 318186 408894
rect 318422 408658 318506 408894
rect 318742 408658 318774 408894
rect 318154 408574 318774 408658
rect 318154 408338 318186 408574
rect 318422 408338 318506 408574
rect 318742 408338 318774 408574
rect 318154 390894 318774 408338
rect 318154 390658 318186 390894
rect 318422 390658 318506 390894
rect 318742 390658 318774 390894
rect 318154 390574 318774 390658
rect 318154 390338 318186 390574
rect 318422 390338 318506 390574
rect 318742 390338 318774 390574
rect 318154 372894 318774 390338
rect 318154 372658 318186 372894
rect 318422 372658 318506 372894
rect 318742 372658 318774 372894
rect 318154 372574 318774 372658
rect 318154 372338 318186 372574
rect 318422 372338 318506 372574
rect 318742 372338 318774 372574
rect 318154 354894 318774 372338
rect 318154 354658 318186 354894
rect 318422 354658 318506 354894
rect 318742 354658 318774 354894
rect 318154 354574 318774 354658
rect 318154 354338 318186 354574
rect 318422 354338 318506 354574
rect 318742 354338 318774 354574
rect 318154 336894 318774 354338
rect 318154 336658 318186 336894
rect 318422 336658 318506 336894
rect 318742 336658 318774 336894
rect 318154 336574 318774 336658
rect 318154 336338 318186 336574
rect 318422 336338 318506 336574
rect 318742 336338 318774 336574
rect 318154 318894 318774 336338
rect 318154 318658 318186 318894
rect 318422 318658 318506 318894
rect 318742 318658 318774 318894
rect 318154 318574 318774 318658
rect 318154 318338 318186 318574
rect 318422 318338 318506 318574
rect 318742 318338 318774 318574
rect 318154 300894 318774 318338
rect 318154 300658 318186 300894
rect 318422 300658 318506 300894
rect 318742 300658 318774 300894
rect 318154 300574 318774 300658
rect 318154 300338 318186 300574
rect 318422 300338 318506 300574
rect 318742 300338 318774 300574
rect 318154 282894 318774 300338
rect 318154 282658 318186 282894
rect 318422 282658 318506 282894
rect 318742 282658 318774 282894
rect 318154 282574 318774 282658
rect 318154 282338 318186 282574
rect 318422 282338 318506 282574
rect 318742 282338 318774 282574
rect 318154 264894 318774 282338
rect 318154 264658 318186 264894
rect 318422 264658 318506 264894
rect 318742 264658 318774 264894
rect 318154 264574 318774 264658
rect 318154 264338 318186 264574
rect 318422 264338 318506 264574
rect 318742 264338 318774 264574
rect 318154 246894 318774 264338
rect 318154 246658 318186 246894
rect 318422 246658 318506 246894
rect 318742 246658 318774 246894
rect 318154 246574 318774 246658
rect 318154 246338 318186 246574
rect 318422 246338 318506 246574
rect 318742 246338 318774 246574
rect 318154 228894 318774 246338
rect 318154 228658 318186 228894
rect 318422 228658 318506 228894
rect 318742 228658 318774 228894
rect 318154 228574 318774 228658
rect 318154 228338 318186 228574
rect 318422 228338 318506 228574
rect 318742 228338 318774 228574
rect 318154 210894 318774 228338
rect 318154 210658 318186 210894
rect 318422 210658 318506 210894
rect 318742 210658 318774 210894
rect 318154 210574 318774 210658
rect 318154 210338 318186 210574
rect 318422 210338 318506 210574
rect 318742 210338 318774 210574
rect 318154 192894 318774 210338
rect 318154 192658 318186 192894
rect 318422 192658 318506 192894
rect 318742 192658 318774 192894
rect 318154 192574 318774 192658
rect 318154 192338 318186 192574
rect 318422 192338 318506 192574
rect 318742 192338 318774 192574
rect 318154 174894 318774 192338
rect 318154 174658 318186 174894
rect 318422 174658 318506 174894
rect 318742 174658 318774 174894
rect 318154 174574 318774 174658
rect 318154 174338 318186 174574
rect 318422 174338 318506 174574
rect 318742 174338 318774 174574
rect 318154 156894 318774 174338
rect 318154 156658 318186 156894
rect 318422 156658 318506 156894
rect 318742 156658 318774 156894
rect 318154 156574 318774 156658
rect 318154 156338 318186 156574
rect 318422 156338 318506 156574
rect 318742 156338 318774 156574
rect 318154 138894 318774 156338
rect 318154 138658 318186 138894
rect 318422 138658 318506 138894
rect 318742 138658 318774 138894
rect 318154 138574 318774 138658
rect 318154 138338 318186 138574
rect 318422 138338 318506 138574
rect 318742 138338 318774 138574
rect 318154 120894 318774 138338
rect 318154 120658 318186 120894
rect 318422 120658 318506 120894
rect 318742 120658 318774 120894
rect 318154 120574 318774 120658
rect 318154 120338 318186 120574
rect 318422 120338 318506 120574
rect 318742 120338 318774 120574
rect 318154 102894 318774 120338
rect 318154 102658 318186 102894
rect 318422 102658 318506 102894
rect 318742 102658 318774 102894
rect 318154 102574 318774 102658
rect 318154 102338 318186 102574
rect 318422 102338 318506 102574
rect 318742 102338 318774 102574
rect 318154 84894 318774 102338
rect 318154 84658 318186 84894
rect 318422 84658 318506 84894
rect 318742 84658 318774 84894
rect 318154 84574 318774 84658
rect 318154 84338 318186 84574
rect 318422 84338 318506 84574
rect 318742 84338 318774 84574
rect 318154 66894 318774 84338
rect 318154 66658 318186 66894
rect 318422 66658 318506 66894
rect 318742 66658 318774 66894
rect 318154 66574 318774 66658
rect 318154 66338 318186 66574
rect 318422 66338 318506 66574
rect 318742 66338 318774 66574
rect 318154 48894 318774 66338
rect 318154 48658 318186 48894
rect 318422 48658 318506 48894
rect 318742 48658 318774 48894
rect 318154 48574 318774 48658
rect 318154 48338 318186 48574
rect 318422 48338 318506 48574
rect 318742 48338 318774 48574
rect 318154 30894 318774 48338
rect 318154 30658 318186 30894
rect 318422 30658 318506 30894
rect 318742 30658 318774 30894
rect 318154 30574 318774 30658
rect 318154 30338 318186 30574
rect 318422 30338 318506 30574
rect 318742 30338 318774 30574
rect 318154 12894 318774 30338
rect 318154 12658 318186 12894
rect 318422 12658 318506 12894
rect 318742 12658 318774 12894
rect 318154 12574 318774 12658
rect 318154 12338 318186 12574
rect 318422 12338 318506 12574
rect 318742 12338 318774 12574
rect 318154 -2776 318774 12338
rect 318154 -3012 318186 -2776
rect 318422 -3012 318506 -2776
rect 318742 -3012 318774 -2776
rect 318154 -3096 318774 -3012
rect 318154 -3332 318186 -3096
rect 318422 -3332 318506 -3096
rect 318742 -3332 318774 -3096
rect 318154 -4324 318774 -3332
rect 321874 463972 322494 464004
rect 321874 463736 321906 463972
rect 322142 463736 322226 463972
rect 322462 463736 322494 463972
rect 321874 463652 322494 463736
rect 321874 463416 321906 463652
rect 322142 463416 322226 463652
rect 322462 463416 322494 463652
rect 321874 448614 322494 463416
rect 321874 448378 321906 448614
rect 322142 448378 322226 448614
rect 322462 448378 322494 448614
rect 321874 448294 322494 448378
rect 321874 448058 321906 448294
rect 322142 448058 322226 448294
rect 322462 448058 322494 448294
rect 321874 430614 322494 448058
rect 321874 430378 321906 430614
rect 322142 430378 322226 430614
rect 322462 430378 322494 430614
rect 321874 430294 322494 430378
rect 321874 430058 321906 430294
rect 322142 430058 322226 430294
rect 322462 430058 322494 430294
rect 321874 412614 322494 430058
rect 321874 412378 321906 412614
rect 322142 412378 322226 412614
rect 322462 412378 322494 412614
rect 321874 412294 322494 412378
rect 321874 412058 321906 412294
rect 322142 412058 322226 412294
rect 322462 412058 322494 412294
rect 321874 394614 322494 412058
rect 321874 394378 321906 394614
rect 322142 394378 322226 394614
rect 322462 394378 322494 394614
rect 321874 394294 322494 394378
rect 321874 394058 321906 394294
rect 322142 394058 322226 394294
rect 322462 394058 322494 394294
rect 321874 376614 322494 394058
rect 321874 376378 321906 376614
rect 322142 376378 322226 376614
rect 322462 376378 322494 376614
rect 321874 376294 322494 376378
rect 321874 376058 321906 376294
rect 322142 376058 322226 376294
rect 322462 376058 322494 376294
rect 321874 358614 322494 376058
rect 321874 358378 321906 358614
rect 322142 358378 322226 358614
rect 322462 358378 322494 358614
rect 321874 358294 322494 358378
rect 321874 358058 321906 358294
rect 322142 358058 322226 358294
rect 322462 358058 322494 358294
rect 321874 340614 322494 358058
rect 321874 340378 321906 340614
rect 322142 340378 322226 340614
rect 322462 340378 322494 340614
rect 321874 340294 322494 340378
rect 321874 340058 321906 340294
rect 322142 340058 322226 340294
rect 322462 340058 322494 340294
rect 321874 322614 322494 340058
rect 321874 322378 321906 322614
rect 322142 322378 322226 322614
rect 322462 322378 322494 322614
rect 321874 322294 322494 322378
rect 321874 322058 321906 322294
rect 322142 322058 322226 322294
rect 322462 322058 322494 322294
rect 321874 304614 322494 322058
rect 321874 304378 321906 304614
rect 322142 304378 322226 304614
rect 322462 304378 322494 304614
rect 321874 304294 322494 304378
rect 321874 304058 321906 304294
rect 322142 304058 322226 304294
rect 322462 304058 322494 304294
rect 321874 286614 322494 304058
rect 321874 286378 321906 286614
rect 322142 286378 322226 286614
rect 322462 286378 322494 286614
rect 321874 286294 322494 286378
rect 321874 286058 321906 286294
rect 322142 286058 322226 286294
rect 322462 286058 322494 286294
rect 321874 268614 322494 286058
rect 321874 268378 321906 268614
rect 322142 268378 322226 268614
rect 322462 268378 322494 268614
rect 321874 268294 322494 268378
rect 321874 268058 321906 268294
rect 322142 268058 322226 268294
rect 322462 268058 322494 268294
rect 321874 250614 322494 268058
rect 321874 250378 321906 250614
rect 322142 250378 322226 250614
rect 322462 250378 322494 250614
rect 321874 250294 322494 250378
rect 321874 250058 321906 250294
rect 322142 250058 322226 250294
rect 322462 250058 322494 250294
rect 321874 232614 322494 250058
rect 321874 232378 321906 232614
rect 322142 232378 322226 232614
rect 322462 232378 322494 232614
rect 321874 232294 322494 232378
rect 321874 232058 321906 232294
rect 322142 232058 322226 232294
rect 322462 232058 322494 232294
rect 321874 214614 322494 232058
rect 321874 214378 321906 214614
rect 322142 214378 322226 214614
rect 322462 214378 322494 214614
rect 321874 214294 322494 214378
rect 321874 214058 321906 214294
rect 322142 214058 322226 214294
rect 322462 214058 322494 214294
rect 321874 196614 322494 214058
rect 321874 196378 321906 196614
rect 322142 196378 322226 196614
rect 322462 196378 322494 196614
rect 321874 196294 322494 196378
rect 321874 196058 321906 196294
rect 322142 196058 322226 196294
rect 322462 196058 322494 196294
rect 321874 178614 322494 196058
rect 321874 178378 321906 178614
rect 322142 178378 322226 178614
rect 322462 178378 322494 178614
rect 321874 178294 322494 178378
rect 321874 178058 321906 178294
rect 322142 178058 322226 178294
rect 322462 178058 322494 178294
rect 321874 160614 322494 178058
rect 321874 160378 321906 160614
rect 322142 160378 322226 160614
rect 322462 160378 322494 160614
rect 321874 160294 322494 160378
rect 321874 160058 321906 160294
rect 322142 160058 322226 160294
rect 322462 160058 322494 160294
rect 321874 142614 322494 160058
rect 321874 142378 321906 142614
rect 322142 142378 322226 142614
rect 322462 142378 322494 142614
rect 321874 142294 322494 142378
rect 321874 142058 321906 142294
rect 322142 142058 322226 142294
rect 322462 142058 322494 142294
rect 321874 124614 322494 142058
rect 321874 124378 321906 124614
rect 322142 124378 322226 124614
rect 322462 124378 322494 124614
rect 321874 124294 322494 124378
rect 321874 124058 321906 124294
rect 322142 124058 322226 124294
rect 322462 124058 322494 124294
rect 321874 106614 322494 124058
rect 321874 106378 321906 106614
rect 322142 106378 322226 106614
rect 322462 106378 322494 106614
rect 321874 106294 322494 106378
rect 321874 106058 321906 106294
rect 322142 106058 322226 106294
rect 322462 106058 322494 106294
rect 321874 88614 322494 106058
rect 321874 88378 321906 88614
rect 322142 88378 322226 88614
rect 322462 88378 322494 88614
rect 321874 88294 322494 88378
rect 321874 88058 321906 88294
rect 322142 88058 322226 88294
rect 322462 88058 322494 88294
rect 321874 70614 322494 88058
rect 321874 70378 321906 70614
rect 322142 70378 322226 70614
rect 322462 70378 322494 70614
rect 321874 70294 322494 70378
rect 321874 70058 321906 70294
rect 322142 70058 322226 70294
rect 322462 70058 322494 70294
rect 321874 52614 322494 70058
rect 321874 52378 321906 52614
rect 322142 52378 322226 52614
rect 322462 52378 322494 52614
rect 321874 52294 322494 52378
rect 321874 52058 321906 52294
rect 322142 52058 322226 52294
rect 322462 52058 322494 52294
rect 321874 34614 322494 52058
rect 321874 34378 321906 34614
rect 322142 34378 322226 34614
rect 322462 34378 322494 34614
rect 321874 34294 322494 34378
rect 321874 34058 321906 34294
rect 322142 34058 322226 34294
rect 322462 34058 322494 34294
rect 321874 16614 322494 34058
rect 321874 16378 321906 16614
rect 322142 16378 322226 16614
rect 322462 16378 322494 16614
rect 321874 16294 322494 16378
rect 321874 16058 321906 16294
rect 322142 16058 322226 16294
rect 322462 16058 322494 16294
rect 321874 -3736 322494 16058
rect 321874 -3972 321906 -3736
rect 322142 -3972 322226 -3736
rect 322462 -3972 322494 -3736
rect 321874 -4056 322494 -3972
rect 321874 -4292 321906 -4056
rect 322142 -4292 322226 -4056
rect 322462 -4292 322494 -4056
rect 321874 -4324 322494 -4292
rect 328714 461092 329334 464004
rect 328714 460856 328746 461092
rect 328982 460856 329066 461092
rect 329302 460856 329334 461092
rect 328714 460772 329334 460856
rect 328714 460536 328746 460772
rect 328982 460536 329066 460772
rect 329302 460536 329334 460772
rect 328714 455454 329334 460536
rect 354154 463012 354774 464004
rect 354154 462776 354186 463012
rect 354422 462776 354506 463012
rect 354742 462776 354774 463012
rect 354154 462692 354774 462776
rect 354154 462456 354186 462692
rect 354422 462456 354506 462692
rect 354742 462456 354774 462692
rect 333993 459700 334121 460000
rect 334505 459700 334633 460000
rect 335017 459700 335145 460000
rect 335529 459700 335657 460000
rect 336041 459700 336169 460000
rect 336553 459700 336681 460000
rect 337065 459700 337193 460000
rect 337577 459700 337705 460000
rect 338089 459700 338217 460000
rect 338601 459700 338729 460000
rect 339113 459700 339241 460000
rect 339625 459700 339753 460000
rect 340137 459700 340265 460000
rect 340649 459700 340777 460000
rect 341161 459700 341289 460000
rect 341673 459700 341801 460000
rect 342185 459700 342313 460000
rect 342697 459700 342825 460000
rect 343209 459700 343337 460000
rect 343721 459700 343849 460000
rect 344233 459700 344361 460000
rect 344745 459700 344873 460000
rect 345257 459700 345385 460000
rect 345769 459700 345897 460000
rect 346281 459700 346409 460000
rect 346793 459700 346921 460000
rect 347305 459700 347433 460000
rect 347817 459700 347945 460000
rect 348329 459700 348457 460000
rect 348841 459700 348969 460000
rect 349353 459700 349481 460000
rect 349865 459700 349993 460000
rect 350377 459700 350505 460000
rect 328714 455218 328746 455454
rect 328982 455218 329066 455454
rect 329302 455218 329334 455454
rect 328714 455134 329334 455218
rect 328714 454898 328746 455134
rect 328982 454898 329066 455134
rect 329302 454898 329334 455134
rect 328714 437454 329334 454898
rect 328714 437218 328746 437454
rect 328982 437218 329066 437454
rect 329302 437218 329334 437454
rect 328714 437134 329334 437218
rect 328714 436898 328746 437134
rect 328982 436898 329066 437134
rect 329302 436898 329334 437134
rect 328714 419454 329334 436898
rect 328714 419218 328746 419454
rect 328982 419218 329066 419454
rect 329302 419218 329334 419454
rect 328714 419134 329334 419218
rect 328714 418898 328746 419134
rect 328982 418898 329066 419134
rect 329302 418898 329334 419134
rect 328714 401454 329334 418898
rect 328714 401218 328746 401454
rect 328982 401218 329066 401454
rect 329302 401218 329334 401454
rect 328714 401134 329334 401218
rect 328714 400898 328746 401134
rect 328982 400898 329066 401134
rect 329302 400898 329334 401134
rect 328714 383454 329334 400898
rect 328714 383218 328746 383454
rect 328982 383218 329066 383454
rect 329302 383218 329334 383454
rect 328714 383134 329334 383218
rect 328714 382898 328746 383134
rect 328982 382898 329066 383134
rect 329302 382898 329334 383134
rect 328714 365454 329334 382898
rect 328714 365218 328746 365454
rect 328982 365218 329066 365454
rect 329302 365218 329334 365454
rect 328714 365134 329334 365218
rect 328714 364898 328746 365134
rect 328982 364898 329066 365134
rect 329302 364898 329334 365134
rect 328714 347454 329334 364898
rect 328714 347218 328746 347454
rect 328982 347218 329066 347454
rect 329302 347218 329334 347454
rect 328714 347134 329334 347218
rect 328714 346898 328746 347134
rect 328982 346898 329066 347134
rect 329302 346898 329334 347134
rect 328714 329454 329334 346898
rect 328714 329218 328746 329454
rect 328982 329218 329066 329454
rect 329302 329218 329334 329454
rect 328714 329134 329334 329218
rect 328714 328898 328746 329134
rect 328982 328898 329066 329134
rect 329302 328898 329334 329134
rect 328714 311454 329334 328898
rect 328714 311218 328746 311454
rect 328982 311218 329066 311454
rect 329302 311218 329334 311454
rect 328714 311134 329334 311218
rect 328714 310898 328746 311134
rect 328982 310898 329066 311134
rect 329302 310898 329334 311134
rect 328714 293454 329334 310898
rect 328714 293218 328746 293454
rect 328982 293218 329066 293454
rect 329302 293218 329334 293454
rect 328714 293134 329334 293218
rect 328714 292898 328746 293134
rect 328982 292898 329066 293134
rect 329302 292898 329334 293134
rect 328714 275454 329334 292898
rect 328714 275218 328746 275454
rect 328982 275218 329066 275454
rect 329302 275218 329334 275454
rect 328714 275134 329334 275218
rect 328714 274898 328746 275134
rect 328982 274898 329066 275134
rect 329302 274898 329334 275134
rect 328714 257454 329334 274898
rect 328714 257218 328746 257454
rect 328982 257218 329066 257454
rect 329302 257218 329334 257454
rect 328714 257134 329334 257218
rect 328714 256898 328746 257134
rect 328982 256898 329066 257134
rect 329302 256898 329334 257134
rect 328714 239454 329334 256898
rect 328714 239218 328746 239454
rect 328982 239218 329066 239454
rect 329302 239218 329334 239454
rect 328714 239134 329334 239218
rect 328714 238898 328746 239134
rect 328982 238898 329066 239134
rect 329302 238898 329334 239134
rect 328714 221454 329334 238898
rect 328714 221218 328746 221454
rect 328982 221218 329066 221454
rect 329302 221218 329334 221454
rect 328714 221134 329334 221218
rect 328714 220898 328746 221134
rect 328982 220898 329066 221134
rect 329302 220898 329334 221134
rect 328714 203454 329334 220898
rect 328714 203218 328746 203454
rect 328982 203218 329066 203454
rect 329302 203218 329334 203454
rect 328714 203134 329334 203218
rect 328714 202898 328746 203134
rect 328982 202898 329066 203134
rect 329302 202898 329334 203134
rect 328714 185454 329334 202898
rect 328714 185218 328746 185454
rect 328982 185218 329066 185454
rect 329302 185218 329334 185454
rect 328714 185134 329334 185218
rect 328714 184898 328746 185134
rect 328982 184898 329066 185134
rect 329302 184898 329334 185134
rect 328714 167454 329334 184898
rect 328714 167218 328746 167454
rect 328982 167218 329066 167454
rect 329302 167218 329334 167454
rect 328714 167134 329334 167218
rect 328714 166898 328746 167134
rect 328982 166898 329066 167134
rect 329302 166898 329334 167134
rect 328714 149454 329334 166898
rect 328714 149218 328746 149454
rect 328982 149218 329066 149454
rect 329302 149218 329334 149454
rect 328714 149134 329334 149218
rect 328714 148898 328746 149134
rect 328982 148898 329066 149134
rect 329302 148898 329334 149134
rect 328714 131454 329334 148898
rect 328714 131218 328746 131454
rect 328982 131218 329066 131454
rect 329302 131218 329334 131454
rect 328714 131134 329334 131218
rect 328714 130898 328746 131134
rect 328982 130898 329066 131134
rect 329302 130898 329334 131134
rect 328714 113454 329334 130898
rect 328714 113218 328746 113454
rect 328982 113218 329066 113454
rect 329302 113218 329334 113454
rect 328714 113134 329334 113218
rect 328714 112898 328746 113134
rect 328982 112898 329066 113134
rect 329302 112898 329334 113134
rect 328714 95454 329334 112898
rect 328714 95218 328746 95454
rect 328982 95218 329066 95454
rect 329302 95218 329334 95454
rect 328714 95134 329334 95218
rect 328714 94898 328746 95134
rect 328982 94898 329066 95134
rect 329302 94898 329334 95134
rect 328714 77454 329334 94898
rect 328714 77218 328746 77454
rect 328982 77218 329066 77454
rect 329302 77218 329334 77454
rect 328714 77134 329334 77218
rect 328714 76898 328746 77134
rect 328982 76898 329066 77134
rect 329302 76898 329334 77134
rect 328714 59454 329334 76898
rect 328714 59218 328746 59454
rect 328982 59218 329066 59454
rect 329302 59218 329334 59454
rect 328714 59134 329334 59218
rect 328714 58898 328746 59134
rect 328982 58898 329066 59134
rect 329302 58898 329334 59134
rect 328714 41454 329334 58898
rect 328714 41218 328746 41454
rect 328982 41218 329066 41454
rect 329302 41218 329334 41454
rect 328714 41134 329334 41218
rect 328714 40898 328746 41134
rect 328982 40898 329066 41134
rect 329302 40898 329334 41134
rect 328714 23454 329334 40898
rect 328714 23218 328746 23454
rect 328982 23218 329066 23454
rect 329302 23218 329334 23454
rect 328714 23134 329334 23218
rect 328714 22898 328746 23134
rect 328982 22898 329066 23134
rect 329302 22898 329334 23134
rect 328714 5454 329334 22898
rect 328714 5218 328746 5454
rect 328982 5218 329066 5454
rect 329302 5218 329334 5454
rect 328714 5134 329334 5218
rect 328714 4898 328746 5134
rect 328982 4898 329066 5134
rect 329302 4898 329334 5134
rect 328714 -856 329334 4898
rect 328714 -1092 328746 -856
rect 328982 -1092 329066 -856
rect 329302 -1092 329334 -856
rect 328714 -1176 329334 -1092
rect 328714 -1412 328746 -1176
rect 328982 -1412 329066 -1176
rect 329302 -1412 329334 -1176
rect 328714 -4324 329334 -1412
rect 332434 441174 333054 458520
rect 332434 440938 332466 441174
rect 332702 440938 332786 441174
rect 333022 440938 333054 441174
rect 332434 440854 333054 440938
rect 332434 440618 332466 440854
rect 332702 440618 332786 440854
rect 333022 440618 333054 440854
rect 332434 423174 333054 440618
rect 332434 422938 332466 423174
rect 332702 422938 332786 423174
rect 333022 422938 333054 423174
rect 332434 422854 333054 422938
rect 332434 422618 332466 422854
rect 332702 422618 332786 422854
rect 333022 422618 333054 422854
rect 332434 405174 333054 422618
rect 332434 404938 332466 405174
rect 332702 404938 332786 405174
rect 333022 404938 333054 405174
rect 332434 404854 333054 404938
rect 332434 404618 332466 404854
rect 332702 404618 332786 404854
rect 333022 404618 333054 404854
rect 332434 387174 333054 404618
rect 332434 386938 332466 387174
rect 332702 386938 332786 387174
rect 333022 386938 333054 387174
rect 332434 386854 333054 386938
rect 332434 386618 332466 386854
rect 332702 386618 332786 386854
rect 333022 386618 333054 386854
rect 332434 369174 333054 386618
rect 332434 368938 332466 369174
rect 332702 368938 332786 369174
rect 333022 368938 333054 369174
rect 332434 368854 333054 368938
rect 332434 368618 332466 368854
rect 332702 368618 332786 368854
rect 333022 368618 333054 368854
rect 332434 351174 333054 368618
rect 332434 350938 332466 351174
rect 332702 350938 332786 351174
rect 333022 350938 333054 351174
rect 332434 350854 333054 350938
rect 332434 350618 332466 350854
rect 332702 350618 332786 350854
rect 333022 350618 333054 350854
rect 332434 333174 333054 350618
rect 332434 332938 332466 333174
rect 332702 332938 332786 333174
rect 333022 332938 333054 333174
rect 332434 332854 333054 332938
rect 332434 332618 332466 332854
rect 332702 332618 332786 332854
rect 333022 332618 333054 332854
rect 332434 315174 333054 332618
rect 332434 314938 332466 315174
rect 332702 314938 332786 315174
rect 333022 314938 333054 315174
rect 332434 314854 333054 314938
rect 332434 314618 332466 314854
rect 332702 314618 332786 314854
rect 333022 314618 333054 314854
rect 332434 297174 333054 314618
rect 332434 296938 332466 297174
rect 332702 296938 332786 297174
rect 333022 296938 333054 297174
rect 332434 296854 333054 296938
rect 332434 296618 332466 296854
rect 332702 296618 332786 296854
rect 333022 296618 333054 296854
rect 332434 279174 333054 296618
rect 332434 278938 332466 279174
rect 332702 278938 332786 279174
rect 333022 278938 333054 279174
rect 332434 278854 333054 278938
rect 332434 278618 332466 278854
rect 332702 278618 332786 278854
rect 333022 278618 333054 278854
rect 332434 261174 333054 278618
rect 332434 260938 332466 261174
rect 332702 260938 332786 261174
rect 333022 260938 333054 261174
rect 332434 260854 333054 260938
rect 332434 260618 332466 260854
rect 332702 260618 332786 260854
rect 333022 260618 333054 260854
rect 332434 243174 333054 260618
rect 332434 242938 332466 243174
rect 332702 242938 332786 243174
rect 333022 242938 333054 243174
rect 332434 242854 333054 242938
rect 332434 242618 332466 242854
rect 332702 242618 332786 242854
rect 333022 242618 333054 242854
rect 332434 225174 333054 242618
rect 332434 224938 332466 225174
rect 332702 224938 332786 225174
rect 333022 224938 333054 225174
rect 332434 224854 333054 224938
rect 332434 224618 332466 224854
rect 332702 224618 332786 224854
rect 333022 224618 333054 224854
rect 332434 207174 333054 224618
rect 332434 206938 332466 207174
rect 332702 206938 332786 207174
rect 333022 206938 333054 207174
rect 332434 206854 333054 206938
rect 332434 206618 332466 206854
rect 332702 206618 332786 206854
rect 333022 206618 333054 206854
rect 332434 189174 333054 206618
rect 332434 188938 332466 189174
rect 332702 188938 332786 189174
rect 333022 188938 333054 189174
rect 332434 188854 333054 188938
rect 332434 188618 332466 188854
rect 332702 188618 332786 188854
rect 333022 188618 333054 188854
rect 332434 171174 333054 188618
rect 332434 170938 332466 171174
rect 332702 170938 332786 171174
rect 333022 170938 333054 171174
rect 332434 170854 333054 170938
rect 332434 170618 332466 170854
rect 332702 170618 332786 170854
rect 333022 170618 333054 170854
rect 332434 153174 333054 170618
rect 332434 152938 332466 153174
rect 332702 152938 332786 153174
rect 333022 152938 333054 153174
rect 332434 152854 333054 152938
rect 332434 152618 332466 152854
rect 332702 152618 332786 152854
rect 333022 152618 333054 152854
rect 332434 135174 333054 152618
rect 332434 134938 332466 135174
rect 332702 134938 332786 135174
rect 333022 134938 333054 135174
rect 332434 134854 333054 134938
rect 332434 134618 332466 134854
rect 332702 134618 332786 134854
rect 333022 134618 333054 134854
rect 332434 117174 333054 134618
rect 332434 116938 332466 117174
rect 332702 116938 332786 117174
rect 333022 116938 333054 117174
rect 332434 116854 333054 116938
rect 332434 116618 332466 116854
rect 332702 116618 332786 116854
rect 333022 116618 333054 116854
rect 332434 99174 333054 116618
rect 332434 98938 332466 99174
rect 332702 98938 332786 99174
rect 333022 98938 333054 99174
rect 332434 98854 333054 98938
rect 332434 98618 332466 98854
rect 332702 98618 332786 98854
rect 333022 98618 333054 98854
rect 332434 81174 333054 98618
rect 332434 80938 332466 81174
rect 332702 80938 332786 81174
rect 333022 80938 333054 81174
rect 332434 80854 333054 80938
rect 332434 80618 332466 80854
rect 332702 80618 332786 80854
rect 333022 80618 333054 80854
rect 332434 63174 333054 80618
rect 332434 62938 332466 63174
rect 332702 62938 332786 63174
rect 333022 62938 333054 63174
rect 332434 62854 333054 62938
rect 332434 62618 332466 62854
rect 332702 62618 332786 62854
rect 333022 62618 333054 62854
rect 332434 45174 333054 62618
rect 332434 44938 332466 45174
rect 332702 44938 332786 45174
rect 333022 44938 333054 45174
rect 332434 44854 333054 44938
rect 332434 44618 332466 44854
rect 332702 44618 332786 44854
rect 333022 44618 333054 44854
rect 332434 27174 333054 44618
rect 332434 26938 332466 27174
rect 332702 26938 332786 27174
rect 333022 26938 333054 27174
rect 332434 26854 333054 26938
rect 332434 26618 332466 26854
rect 332702 26618 332786 26854
rect 333022 26618 333054 26854
rect 332434 9174 333054 26618
rect 332434 8938 332466 9174
rect 332702 8938 332786 9174
rect 333022 8938 333054 9174
rect 332434 8854 333054 8938
rect 332434 8618 332466 8854
rect 332702 8618 332786 8854
rect 333022 8618 333054 8854
rect 332434 -1816 333054 8618
rect 332434 -2052 332466 -1816
rect 332702 -2052 332786 -1816
rect 333022 -2052 333054 -1816
rect 332434 -2136 333054 -2052
rect 332434 -2372 332466 -2136
rect 332702 -2372 332786 -2136
rect 333022 -2372 333054 -2136
rect 332434 -4324 333054 -2372
rect 336154 444894 336774 458520
rect 336154 444658 336186 444894
rect 336422 444658 336506 444894
rect 336742 444658 336774 444894
rect 336154 444574 336774 444658
rect 336154 444338 336186 444574
rect 336422 444338 336506 444574
rect 336742 444338 336774 444574
rect 336154 426894 336774 444338
rect 336154 426658 336186 426894
rect 336422 426658 336506 426894
rect 336742 426658 336774 426894
rect 336154 426574 336774 426658
rect 336154 426338 336186 426574
rect 336422 426338 336506 426574
rect 336742 426338 336774 426574
rect 336154 408894 336774 426338
rect 336154 408658 336186 408894
rect 336422 408658 336506 408894
rect 336742 408658 336774 408894
rect 336154 408574 336774 408658
rect 336154 408338 336186 408574
rect 336422 408338 336506 408574
rect 336742 408338 336774 408574
rect 336154 390894 336774 408338
rect 336154 390658 336186 390894
rect 336422 390658 336506 390894
rect 336742 390658 336774 390894
rect 336154 390574 336774 390658
rect 336154 390338 336186 390574
rect 336422 390338 336506 390574
rect 336742 390338 336774 390574
rect 336154 372894 336774 390338
rect 336154 372658 336186 372894
rect 336422 372658 336506 372894
rect 336742 372658 336774 372894
rect 336154 372574 336774 372658
rect 336154 372338 336186 372574
rect 336422 372338 336506 372574
rect 336742 372338 336774 372574
rect 336154 354894 336774 372338
rect 336154 354658 336186 354894
rect 336422 354658 336506 354894
rect 336742 354658 336774 354894
rect 336154 354574 336774 354658
rect 336154 354338 336186 354574
rect 336422 354338 336506 354574
rect 336742 354338 336774 354574
rect 336154 336894 336774 354338
rect 336154 336658 336186 336894
rect 336422 336658 336506 336894
rect 336742 336658 336774 336894
rect 336154 336574 336774 336658
rect 336154 336338 336186 336574
rect 336422 336338 336506 336574
rect 336742 336338 336774 336574
rect 336154 318894 336774 336338
rect 336154 318658 336186 318894
rect 336422 318658 336506 318894
rect 336742 318658 336774 318894
rect 336154 318574 336774 318658
rect 336154 318338 336186 318574
rect 336422 318338 336506 318574
rect 336742 318338 336774 318574
rect 336154 300894 336774 318338
rect 336154 300658 336186 300894
rect 336422 300658 336506 300894
rect 336742 300658 336774 300894
rect 336154 300574 336774 300658
rect 336154 300338 336186 300574
rect 336422 300338 336506 300574
rect 336742 300338 336774 300574
rect 336154 282894 336774 300338
rect 336154 282658 336186 282894
rect 336422 282658 336506 282894
rect 336742 282658 336774 282894
rect 336154 282574 336774 282658
rect 336154 282338 336186 282574
rect 336422 282338 336506 282574
rect 336742 282338 336774 282574
rect 336154 264894 336774 282338
rect 336154 264658 336186 264894
rect 336422 264658 336506 264894
rect 336742 264658 336774 264894
rect 336154 264574 336774 264658
rect 336154 264338 336186 264574
rect 336422 264338 336506 264574
rect 336742 264338 336774 264574
rect 336154 246894 336774 264338
rect 336154 246658 336186 246894
rect 336422 246658 336506 246894
rect 336742 246658 336774 246894
rect 336154 246574 336774 246658
rect 336154 246338 336186 246574
rect 336422 246338 336506 246574
rect 336742 246338 336774 246574
rect 336154 228894 336774 246338
rect 336154 228658 336186 228894
rect 336422 228658 336506 228894
rect 336742 228658 336774 228894
rect 336154 228574 336774 228658
rect 336154 228338 336186 228574
rect 336422 228338 336506 228574
rect 336742 228338 336774 228574
rect 336154 210894 336774 228338
rect 336154 210658 336186 210894
rect 336422 210658 336506 210894
rect 336742 210658 336774 210894
rect 336154 210574 336774 210658
rect 336154 210338 336186 210574
rect 336422 210338 336506 210574
rect 336742 210338 336774 210574
rect 336154 192894 336774 210338
rect 336154 192658 336186 192894
rect 336422 192658 336506 192894
rect 336742 192658 336774 192894
rect 336154 192574 336774 192658
rect 336154 192338 336186 192574
rect 336422 192338 336506 192574
rect 336742 192338 336774 192574
rect 336154 174894 336774 192338
rect 336154 174658 336186 174894
rect 336422 174658 336506 174894
rect 336742 174658 336774 174894
rect 336154 174574 336774 174658
rect 336154 174338 336186 174574
rect 336422 174338 336506 174574
rect 336742 174338 336774 174574
rect 336154 156894 336774 174338
rect 336154 156658 336186 156894
rect 336422 156658 336506 156894
rect 336742 156658 336774 156894
rect 336154 156574 336774 156658
rect 336154 156338 336186 156574
rect 336422 156338 336506 156574
rect 336742 156338 336774 156574
rect 336154 138894 336774 156338
rect 336154 138658 336186 138894
rect 336422 138658 336506 138894
rect 336742 138658 336774 138894
rect 336154 138574 336774 138658
rect 336154 138338 336186 138574
rect 336422 138338 336506 138574
rect 336742 138338 336774 138574
rect 336154 120894 336774 138338
rect 336154 120658 336186 120894
rect 336422 120658 336506 120894
rect 336742 120658 336774 120894
rect 336154 120574 336774 120658
rect 336154 120338 336186 120574
rect 336422 120338 336506 120574
rect 336742 120338 336774 120574
rect 336154 102894 336774 120338
rect 336154 102658 336186 102894
rect 336422 102658 336506 102894
rect 336742 102658 336774 102894
rect 336154 102574 336774 102658
rect 336154 102338 336186 102574
rect 336422 102338 336506 102574
rect 336742 102338 336774 102574
rect 336154 84894 336774 102338
rect 336154 84658 336186 84894
rect 336422 84658 336506 84894
rect 336742 84658 336774 84894
rect 336154 84574 336774 84658
rect 336154 84338 336186 84574
rect 336422 84338 336506 84574
rect 336742 84338 336774 84574
rect 336154 66894 336774 84338
rect 336154 66658 336186 66894
rect 336422 66658 336506 66894
rect 336742 66658 336774 66894
rect 336154 66574 336774 66658
rect 336154 66338 336186 66574
rect 336422 66338 336506 66574
rect 336742 66338 336774 66574
rect 336154 48894 336774 66338
rect 336154 48658 336186 48894
rect 336422 48658 336506 48894
rect 336742 48658 336774 48894
rect 336154 48574 336774 48658
rect 336154 48338 336186 48574
rect 336422 48338 336506 48574
rect 336742 48338 336774 48574
rect 336154 30894 336774 48338
rect 336154 30658 336186 30894
rect 336422 30658 336506 30894
rect 336742 30658 336774 30894
rect 336154 30574 336774 30658
rect 336154 30338 336186 30574
rect 336422 30338 336506 30574
rect 336742 30338 336774 30574
rect 336154 12894 336774 30338
rect 336154 12658 336186 12894
rect 336422 12658 336506 12894
rect 336742 12658 336774 12894
rect 336154 12574 336774 12658
rect 336154 12338 336186 12574
rect 336422 12338 336506 12574
rect 336742 12338 336774 12574
rect 336154 -2776 336774 12338
rect 336154 -3012 336186 -2776
rect 336422 -3012 336506 -2776
rect 336742 -3012 336774 -2776
rect 336154 -3096 336774 -3012
rect 336154 -3332 336186 -3096
rect 336422 -3332 336506 -3096
rect 336742 -3332 336774 -3096
rect 336154 -4324 336774 -3332
rect 339874 448614 340494 458520
rect 339874 448378 339906 448614
rect 340142 448378 340226 448614
rect 340462 448378 340494 448614
rect 339874 448294 340494 448378
rect 339874 448058 339906 448294
rect 340142 448058 340226 448294
rect 340462 448058 340494 448294
rect 339874 430614 340494 448058
rect 339874 430378 339906 430614
rect 340142 430378 340226 430614
rect 340462 430378 340494 430614
rect 339874 430294 340494 430378
rect 339874 430058 339906 430294
rect 340142 430058 340226 430294
rect 340462 430058 340494 430294
rect 339874 412614 340494 430058
rect 339874 412378 339906 412614
rect 340142 412378 340226 412614
rect 340462 412378 340494 412614
rect 339874 412294 340494 412378
rect 339874 412058 339906 412294
rect 340142 412058 340226 412294
rect 340462 412058 340494 412294
rect 339874 394614 340494 412058
rect 339874 394378 339906 394614
rect 340142 394378 340226 394614
rect 340462 394378 340494 394614
rect 339874 394294 340494 394378
rect 339874 394058 339906 394294
rect 340142 394058 340226 394294
rect 340462 394058 340494 394294
rect 339874 376614 340494 394058
rect 339874 376378 339906 376614
rect 340142 376378 340226 376614
rect 340462 376378 340494 376614
rect 339874 376294 340494 376378
rect 339874 376058 339906 376294
rect 340142 376058 340226 376294
rect 340462 376058 340494 376294
rect 339874 358614 340494 376058
rect 339874 358378 339906 358614
rect 340142 358378 340226 358614
rect 340462 358378 340494 358614
rect 339874 358294 340494 358378
rect 339874 358058 339906 358294
rect 340142 358058 340226 358294
rect 340462 358058 340494 358294
rect 339874 340614 340494 358058
rect 339874 340378 339906 340614
rect 340142 340378 340226 340614
rect 340462 340378 340494 340614
rect 339874 340294 340494 340378
rect 339874 340058 339906 340294
rect 340142 340058 340226 340294
rect 340462 340058 340494 340294
rect 339874 322614 340494 340058
rect 339874 322378 339906 322614
rect 340142 322378 340226 322614
rect 340462 322378 340494 322614
rect 339874 322294 340494 322378
rect 339874 322058 339906 322294
rect 340142 322058 340226 322294
rect 340462 322058 340494 322294
rect 339874 304614 340494 322058
rect 339874 304378 339906 304614
rect 340142 304378 340226 304614
rect 340462 304378 340494 304614
rect 339874 304294 340494 304378
rect 339874 304058 339906 304294
rect 340142 304058 340226 304294
rect 340462 304058 340494 304294
rect 339874 286614 340494 304058
rect 339874 286378 339906 286614
rect 340142 286378 340226 286614
rect 340462 286378 340494 286614
rect 339874 286294 340494 286378
rect 339874 286058 339906 286294
rect 340142 286058 340226 286294
rect 340462 286058 340494 286294
rect 339874 268614 340494 286058
rect 339874 268378 339906 268614
rect 340142 268378 340226 268614
rect 340462 268378 340494 268614
rect 339874 268294 340494 268378
rect 339874 268058 339906 268294
rect 340142 268058 340226 268294
rect 340462 268058 340494 268294
rect 339874 250614 340494 268058
rect 339874 250378 339906 250614
rect 340142 250378 340226 250614
rect 340462 250378 340494 250614
rect 339874 250294 340494 250378
rect 339874 250058 339906 250294
rect 340142 250058 340226 250294
rect 340462 250058 340494 250294
rect 339874 232614 340494 250058
rect 339874 232378 339906 232614
rect 340142 232378 340226 232614
rect 340462 232378 340494 232614
rect 339874 232294 340494 232378
rect 339874 232058 339906 232294
rect 340142 232058 340226 232294
rect 340462 232058 340494 232294
rect 339874 214614 340494 232058
rect 339874 214378 339906 214614
rect 340142 214378 340226 214614
rect 340462 214378 340494 214614
rect 339874 214294 340494 214378
rect 339874 214058 339906 214294
rect 340142 214058 340226 214294
rect 340462 214058 340494 214294
rect 339874 196614 340494 214058
rect 339874 196378 339906 196614
rect 340142 196378 340226 196614
rect 340462 196378 340494 196614
rect 339874 196294 340494 196378
rect 339874 196058 339906 196294
rect 340142 196058 340226 196294
rect 340462 196058 340494 196294
rect 339874 178614 340494 196058
rect 339874 178378 339906 178614
rect 340142 178378 340226 178614
rect 340462 178378 340494 178614
rect 339874 178294 340494 178378
rect 339874 178058 339906 178294
rect 340142 178058 340226 178294
rect 340462 178058 340494 178294
rect 339874 160614 340494 178058
rect 339874 160378 339906 160614
rect 340142 160378 340226 160614
rect 340462 160378 340494 160614
rect 339874 160294 340494 160378
rect 339874 160058 339906 160294
rect 340142 160058 340226 160294
rect 340462 160058 340494 160294
rect 339874 142614 340494 160058
rect 339874 142378 339906 142614
rect 340142 142378 340226 142614
rect 340462 142378 340494 142614
rect 339874 142294 340494 142378
rect 339874 142058 339906 142294
rect 340142 142058 340226 142294
rect 340462 142058 340494 142294
rect 339874 124614 340494 142058
rect 339874 124378 339906 124614
rect 340142 124378 340226 124614
rect 340462 124378 340494 124614
rect 339874 124294 340494 124378
rect 339874 124058 339906 124294
rect 340142 124058 340226 124294
rect 340462 124058 340494 124294
rect 339874 106614 340494 124058
rect 339874 106378 339906 106614
rect 340142 106378 340226 106614
rect 340462 106378 340494 106614
rect 339874 106294 340494 106378
rect 339874 106058 339906 106294
rect 340142 106058 340226 106294
rect 340462 106058 340494 106294
rect 339874 88614 340494 106058
rect 339874 88378 339906 88614
rect 340142 88378 340226 88614
rect 340462 88378 340494 88614
rect 339874 88294 340494 88378
rect 339874 88058 339906 88294
rect 340142 88058 340226 88294
rect 340462 88058 340494 88294
rect 339874 70614 340494 88058
rect 339874 70378 339906 70614
rect 340142 70378 340226 70614
rect 340462 70378 340494 70614
rect 339874 70294 340494 70378
rect 339874 70058 339906 70294
rect 340142 70058 340226 70294
rect 340462 70058 340494 70294
rect 339874 52614 340494 70058
rect 339874 52378 339906 52614
rect 340142 52378 340226 52614
rect 340462 52378 340494 52614
rect 339874 52294 340494 52378
rect 339874 52058 339906 52294
rect 340142 52058 340226 52294
rect 340462 52058 340494 52294
rect 339874 34614 340494 52058
rect 339874 34378 339906 34614
rect 340142 34378 340226 34614
rect 340462 34378 340494 34614
rect 339874 34294 340494 34378
rect 339874 34058 339906 34294
rect 340142 34058 340226 34294
rect 340462 34058 340494 34294
rect 339874 16614 340494 34058
rect 339874 16378 339906 16614
rect 340142 16378 340226 16614
rect 340462 16378 340494 16614
rect 339874 16294 340494 16378
rect 339874 16058 339906 16294
rect 340142 16058 340226 16294
rect 340462 16058 340494 16294
rect 339874 -3736 340494 16058
rect 339874 -3972 339906 -3736
rect 340142 -3972 340226 -3736
rect 340462 -3972 340494 -3736
rect 339874 -4056 340494 -3972
rect 339874 -4292 339906 -4056
rect 340142 -4292 340226 -4056
rect 340462 -4292 340494 -4056
rect 339874 -4324 340494 -4292
rect 346714 455454 347334 458520
rect 346714 455218 346746 455454
rect 346982 455218 347066 455454
rect 347302 455218 347334 455454
rect 346714 455134 347334 455218
rect 346714 454898 346746 455134
rect 346982 454898 347066 455134
rect 347302 454898 347334 455134
rect 346714 437454 347334 454898
rect 346714 437218 346746 437454
rect 346982 437218 347066 437454
rect 347302 437218 347334 437454
rect 346714 437134 347334 437218
rect 346714 436898 346746 437134
rect 346982 436898 347066 437134
rect 347302 436898 347334 437134
rect 346714 419454 347334 436898
rect 346714 419218 346746 419454
rect 346982 419218 347066 419454
rect 347302 419218 347334 419454
rect 346714 419134 347334 419218
rect 346714 418898 346746 419134
rect 346982 418898 347066 419134
rect 347302 418898 347334 419134
rect 346714 401454 347334 418898
rect 346714 401218 346746 401454
rect 346982 401218 347066 401454
rect 347302 401218 347334 401454
rect 346714 401134 347334 401218
rect 346714 400898 346746 401134
rect 346982 400898 347066 401134
rect 347302 400898 347334 401134
rect 346714 383454 347334 400898
rect 346714 383218 346746 383454
rect 346982 383218 347066 383454
rect 347302 383218 347334 383454
rect 346714 383134 347334 383218
rect 346714 382898 346746 383134
rect 346982 382898 347066 383134
rect 347302 382898 347334 383134
rect 346714 365454 347334 382898
rect 346714 365218 346746 365454
rect 346982 365218 347066 365454
rect 347302 365218 347334 365454
rect 346714 365134 347334 365218
rect 346714 364898 346746 365134
rect 346982 364898 347066 365134
rect 347302 364898 347334 365134
rect 346714 347454 347334 364898
rect 346714 347218 346746 347454
rect 346982 347218 347066 347454
rect 347302 347218 347334 347454
rect 346714 347134 347334 347218
rect 346714 346898 346746 347134
rect 346982 346898 347066 347134
rect 347302 346898 347334 347134
rect 346714 329454 347334 346898
rect 346714 329218 346746 329454
rect 346982 329218 347066 329454
rect 347302 329218 347334 329454
rect 346714 329134 347334 329218
rect 346714 328898 346746 329134
rect 346982 328898 347066 329134
rect 347302 328898 347334 329134
rect 346714 311454 347334 328898
rect 346714 311218 346746 311454
rect 346982 311218 347066 311454
rect 347302 311218 347334 311454
rect 346714 311134 347334 311218
rect 346714 310898 346746 311134
rect 346982 310898 347066 311134
rect 347302 310898 347334 311134
rect 346714 293454 347334 310898
rect 346714 293218 346746 293454
rect 346982 293218 347066 293454
rect 347302 293218 347334 293454
rect 346714 293134 347334 293218
rect 346714 292898 346746 293134
rect 346982 292898 347066 293134
rect 347302 292898 347334 293134
rect 346714 275454 347334 292898
rect 346714 275218 346746 275454
rect 346982 275218 347066 275454
rect 347302 275218 347334 275454
rect 346714 275134 347334 275218
rect 346714 274898 346746 275134
rect 346982 274898 347066 275134
rect 347302 274898 347334 275134
rect 346714 257454 347334 274898
rect 346714 257218 346746 257454
rect 346982 257218 347066 257454
rect 347302 257218 347334 257454
rect 346714 257134 347334 257218
rect 346714 256898 346746 257134
rect 346982 256898 347066 257134
rect 347302 256898 347334 257134
rect 346714 239454 347334 256898
rect 346714 239218 346746 239454
rect 346982 239218 347066 239454
rect 347302 239218 347334 239454
rect 346714 239134 347334 239218
rect 346714 238898 346746 239134
rect 346982 238898 347066 239134
rect 347302 238898 347334 239134
rect 346714 221454 347334 238898
rect 346714 221218 346746 221454
rect 346982 221218 347066 221454
rect 347302 221218 347334 221454
rect 346714 221134 347334 221218
rect 346714 220898 346746 221134
rect 346982 220898 347066 221134
rect 347302 220898 347334 221134
rect 346714 203454 347334 220898
rect 346714 203218 346746 203454
rect 346982 203218 347066 203454
rect 347302 203218 347334 203454
rect 346714 203134 347334 203218
rect 346714 202898 346746 203134
rect 346982 202898 347066 203134
rect 347302 202898 347334 203134
rect 346714 185454 347334 202898
rect 346714 185218 346746 185454
rect 346982 185218 347066 185454
rect 347302 185218 347334 185454
rect 346714 185134 347334 185218
rect 346714 184898 346746 185134
rect 346982 184898 347066 185134
rect 347302 184898 347334 185134
rect 346714 167454 347334 184898
rect 346714 167218 346746 167454
rect 346982 167218 347066 167454
rect 347302 167218 347334 167454
rect 346714 167134 347334 167218
rect 346714 166898 346746 167134
rect 346982 166898 347066 167134
rect 347302 166898 347334 167134
rect 346714 149454 347334 166898
rect 346714 149218 346746 149454
rect 346982 149218 347066 149454
rect 347302 149218 347334 149454
rect 346714 149134 347334 149218
rect 346714 148898 346746 149134
rect 346982 148898 347066 149134
rect 347302 148898 347334 149134
rect 346714 131454 347334 148898
rect 346714 131218 346746 131454
rect 346982 131218 347066 131454
rect 347302 131218 347334 131454
rect 346714 131134 347334 131218
rect 346714 130898 346746 131134
rect 346982 130898 347066 131134
rect 347302 130898 347334 131134
rect 346714 113454 347334 130898
rect 346714 113218 346746 113454
rect 346982 113218 347066 113454
rect 347302 113218 347334 113454
rect 346714 113134 347334 113218
rect 346714 112898 346746 113134
rect 346982 112898 347066 113134
rect 347302 112898 347334 113134
rect 346714 95454 347334 112898
rect 346714 95218 346746 95454
rect 346982 95218 347066 95454
rect 347302 95218 347334 95454
rect 346714 95134 347334 95218
rect 346714 94898 346746 95134
rect 346982 94898 347066 95134
rect 347302 94898 347334 95134
rect 346714 77454 347334 94898
rect 346714 77218 346746 77454
rect 346982 77218 347066 77454
rect 347302 77218 347334 77454
rect 346714 77134 347334 77218
rect 346714 76898 346746 77134
rect 346982 76898 347066 77134
rect 347302 76898 347334 77134
rect 346714 59454 347334 76898
rect 346714 59218 346746 59454
rect 346982 59218 347066 59454
rect 347302 59218 347334 59454
rect 346714 59134 347334 59218
rect 346714 58898 346746 59134
rect 346982 58898 347066 59134
rect 347302 58898 347334 59134
rect 346714 41454 347334 58898
rect 346714 41218 346746 41454
rect 346982 41218 347066 41454
rect 347302 41218 347334 41454
rect 346714 41134 347334 41218
rect 346714 40898 346746 41134
rect 346982 40898 347066 41134
rect 347302 40898 347334 41134
rect 346714 23454 347334 40898
rect 346714 23218 346746 23454
rect 346982 23218 347066 23454
rect 347302 23218 347334 23454
rect 346714 23134 347334 23218
rect 346714 22898 346746 23134
rect 346982 22898 347066 23134
rect 347302 22898 347334 23134
rect 346714 5454 347334 22898
rect 346714 5218 346746 5454
rect 346982 5218 347066 5454
rect 347302 5218 347334 5454
rect 346714 5134 347334 5218
rect 346714 4898 346746 5134
rect 346982 4898 347066 5134
rect 347302 4898 347334 5134
rect 346714 -856 347334 4898
rect 346714 -1092 346746 -856
rect 346982 -1092 347066 -856
rect 347302 -1092 347334 -856
rect 346714 -1176 347334 -1092
rect 346714 -1412 346746 -1176
rect 346982 -1412 347066 -1176
rect 347302 -1412 347334 -1176
rect 346714 -4324 347334 -1412
rect 350434 441174 351054 458520
rect 350434 440938 350466 441174
rect 350702 440938 350786 441174
rect 351022 440938 351054 441174
rect 350434 440854 351054 440938
rect 350434 440618 350466 440854
rect 350702 440618 350786 440854
rect 351022 440618 351054 440854
rect 350434 423174 351054 440618
rect 350434 422938 350466 423174
rect 350702 422938 350786 423174
rect 351022 422938 351054 423174
rect 350434 422854 351054 422938
rect 350434 422618 350466 422854
rect 350702 422618 350786 422854
rect 351022 422618 351054 422854
rect 350434 405174 351054 422618
rect 350434 404938 350466 405174
rect 350702 404938 350786 405174
rect 351022 404938 351054 405174
rect 350434 404854 351054 404938
rect 350434 404618 350466 404854
rect 350702 404618 350786 404854
rect 351022 404618 351054 404854
rect 350434 387174 351054 404618
rect 350434 386938 350466 387174
rect 350702 386938 350786 387174
rect 351022 386938 351054 387174
rect 350434 386854 351054 386938
rect 350434 386618 350466 386854
rect 350702 386618 350786 386854
rect 351022 386618 351054 386854
rect 350434 369174 351054 386618
rect 350434 368938 350466 369174
rect 350702 368938 350786 369174
rect 351022 368938 351054 369174
rect 350434 368854 351054 368938
rect 350434 368618 350466 368854
rect 350702 368618 350786 368854
rect 351022 368618 351054 368854
rect 350434 351174 351054 368618
rect 350434 350938 350466 351174
rect 350702 350938 350786 351174
rect 351022 350938 351054 351174
rect 350434 350854 351054 350938
rect 350434 350618 350466 350854
rect 350702 350618 350786 350854
rect 351022 350618 351054 350854
rect 350434 333174 351054 350618
rect 350434 332938 350466 333174
rect 350702 332938 350786 333174
rect 351022 332938 351054 333174
rect 350434 332854 351054 332938
rect 350434 332618 350466 332854
rect 350702 332618 350786 332854
rect 351022 332618 351054 332854
rect 350434 315174 351054 332618
rect 350434 314938 350466 315174
rect 350702 314938 350786 315174
rect 351022 314938 351054 315174
rect 350434 314854 351054 314938
rect 350434 314618 350466 314854
rect 350702 314618 350786 314854
rect 351022 314618 351054 314854
rect 350434 297174 351054 314618
rect 350434 296938 350466 297174
rect 350702 296938 350786 297174
rect 351022 296938 351054 297174
rect 350434 296854 351054 296938
rect 350434 296618 350466 296854
rect 350702 296618 350786 296854
rect 351022 296618 351054 296854
rect 350434 279174 351054 296618
rect 350434 278938 350466 279174
rect 350702 278938 350786 279174
rect 351022 278938 351054 279174
rect 350434 278854 351054 278938
rect 350434 278618 350466 278854
rect 350702 278618 350786 278854
rect 351022 278618 351054 278854
rect 350434 261174 351054 278618
rect 350434 260938 350466 261174
rect 350702 260938 350786 261174
rect 351022 260938 351054 261174
rect 350434 260854 351054 260938
rect 350434 260618 350466 260854
rect 350702 260618 350786 260854
rect 351022 260618 351054 260854
rect 350434 243174 351054 260618
rect 350434 242938 350466 243174
rect 350702 242938 350786 243174
rect 351022 242938 351054 243174
rect 350434 242854 351054 242938
rect 350434 242618 350466 242854
rect 350702 242618 350786 242854
rect 351022 242618 351054 242854
rect 350434 225174 351054 242618
rect 350434 224938 350466 225174
rect 350702 224938 350786 225174
rect 351022 224938 351054 225174
rect 350434 224854 351054 224938
rect 350434 224618 350466 224854
rect 350702 224618 350786 224854
rect 351022 224618 351054 224854
rect 350434 207174 351054 224618
rect 350434 206938 350466 207174
rect 350702 206938 350786 207174
rect 351022 206938 351054 207174
rect 350434 206854 351054 206938
rect 350434 206618 350466 206854
rect 350702 206618 350786 206854
rect 351022 206618 351054 206854
rect 350434 189174 351054 206618
rect 350434 188938 350466 189174
rect 350702 188938 350786 189174
rect 351022 188938 351054 189174
rect 350434 188854 351054 188938
rect 350434 188618 350466 188854
rect 350702 188618 350786 188854
rect 351022 188618 351054 188854
rect 350434 171174 351054 188618
rect 350434 170938 350466 171174
rect 350702 170938 350786 171174
rect 351022 170938 351054 171174
rect 350434 170854 351054 170938
rect 350434 170618 350466 170854
rect 350702 170618 350786 170854
rect 351022 170618 351054 170854
rect 350434 153174 351054 170618
rect 350434 152938 350466 153174
rect 350702 152938 350786 153174
rect 351022 152938 351054 153174
rect 350434 152854 351054 152938
rect 350434 152618 350466 152854
rect 350702 152618 350786 152854
rect 351022 152618 351054 152854
rect 350434 135174 351054 152618
rect 350434 134938 350466 135174
rect 350702 134938 350786 135174
rect 351022 134938 351054 135174
rect 350434 134854 351054 134938
rect 350434 134618 350466 134854
rect 350702 134618 350786 134854
rect 351022 134618 351054 134854
rect 350434 117174 351054 134618
rect 350434 116938 350466 117174
rect 350702 116938 350786 117174
rect 351022 116938 351054 117174
rect 350434 116854 351054 116938
rect 350434 116618 350466 116854
rect 350702 116618 350786 116854
rect 351022 116618 351054 116854
rect 350434 99174 351054 116618
rect 350434 98938 350466 99174
rect 350702 98938 350786 99174
rect 351022 98938 351054 99174
rect 350434 98854 351054 98938
rect 350434 98618 350466 98854
rect 350702 98618 350786 98854
rect 351022 98618 351054 98854
rect 350434 81174 351054 98618
rect 350434 80938 350466 81174
rect 350702 80938 350786 81174
rect 351022 80938 351054 81174
rect 350434 80854 351054 80938
rect 350434 80618 350466 80854
rect 350702 80618 350786 80854
rect 351022 80618 351054 80854
rect 350434 63174 351054 80618
rect 350434 62938 350466 63174
rect 350702 62938 350786 63174
rect 351022 62938 351054 63174
rect 350434 62854 351054 62938
rect 350434 62618 350466 62854
rect 350702 62618 350786 62854
rect 351022 62618 351054 62854
rect 350434 45174 351054 62618
rect 350434 44938 350466 45174
rect 350702 44938 350786 45174
rect 351022 44938 351054 45174
rect 350434 44854 351054 44938
rect 350434 44618 350466 44854
rect 350702 44618 350786 44854
rect 351022 44618 351054 44854
rect 350434 27174 351054 44618
rect 350434 26938 350466 27174
rect 350702 26938 350786 27174
rect 351022 26938 351054 27174
rect 350434 26854 351054 26938
rect 350434 26618 350466 26854
rect 350702 26618 350786 26854
rect 351022 26618 351054 26854
rect 350434 9174 351054 26618
rect 350434 8938 350466 9174
rect 350702 8938 350786 9174
rect 351022 8938 351054 9174
rect 350434 8854 351054 8938
rect 350434 8618 350466 8854
rect 350702 8618 350786 8854
rect 351022 8618 351054 8854
rect 350434 -1816 351054 8618
rect 350434 -2052 350466 -1816
rect 350702 -2052 350786 -1816
rect 351022 -2052 351054 -1816
rect 350434 -2136 351054 -2052
rect 350434 -2372 350466 -2136
rect 350702 -2372 350786 -2136
rect 351022 -2372 351054 -2136
rect 350434 -4324 351054 -2372
rect 354154 444894 354774 462456
rect 354154 444658 354186 444894
rect 354422 444658 354506 444894
rect 354742 444658 354774 444894
rect 354154 444574 354774 444658
rect 354154 444338 354186 444574
rect 354422 444338 354506 444574
rect 354742 444338 354774 444574
rect 354154 426894 354774 444338
rect 354154 426658 354186 426894
rect 354422 426658 354506 426894
rect 354742 426658 354774 426894
rect 354154 426574 354774 426658
rect 354154 426338 354186 426574
rect 354422 426338 354506 426574
rect 354742 426338 354774 426574
rect 354154 408894 354774 426338
rect 354154 408658 354186 408894
rect 354422 408658 354506 408894
rect 354742 408658 354774 408894
rect 354154 408574 354774 408658
rect 354154 408338 354186 408574
rect 354422 408338 354506 408574
rect 354742 408338 354774 408574
rect 354154 390894 354774 408338
rect 354154 390658 354186 390894
rect 354422 390658 354506 390894
rect 354742 390658 354774 390894
rect 354154 390574 354774 390658
rect 354154 390338 354186 390574
rect 354422 390338 354506 390574
rect 354742 390338 354774 390574
rect 354154 372894 354774 390338
rect 354154 372658 354186 372894
rect 354422 372658 354506 372894
rect 354742 372658 354774 372894
rect 354154 372574 354774 372658
rect 354154 372338 354186 372574
rect 354422 372338 354506 372574
rect 354742 372338 354774 372574
rect 354154 354894 354774 372338
rect 354154 354658 354186 354894
rect 354422 354658 354506 354894
rect 354742 354658 354774 354894
rect 354154 354574 354774 354658
rect 354154 354338 354186 354574
rect 354422 354338 354506 354574
rect 354742 354338 354774 354574
rect 354154 336894 354774 354338
rect 354154 336658 354186 336894
rect 354422 336658 354506 336894
rect 354742 336658 354774 336894
rect 354154 336574 354774 336658
rect 354154 336338 354186 336574
rect 354422 336338 354506 336574
rect 354742 336338 354774 336574
rect 354154 318894 354774 336338
rect 354154 318658 354186 318894
rect 354422 318658 354506 318894
rect 354742 318658 354774 318894
rect 354154 318574 354774 318658
rect 354154 318338 354186 318574
rect 354422 318338 354506 318574
rect 354742 318338 354774 318574
rect 354154 300894 354774 318338
rect 354154 300658 354186 300894
rect 354422 300658 354506 300894
rect 354742 300658 354774 300894
rect 354154 300574 354774 300658
rect 354154 300338 354186 300574
rect 354422 300338 354506 300574
rect 354742 300338 354774 300574
rect 354154 282894 354774 300338
rect 354154 282658 354186 282894
rect 354422 282658 354506 282894
rect 354742 282658 354774 282894
rect 354154 282574 354774 282658
rect 354154 282338 354186 282574
rect 354422 282338 354506 282574
rect 354742 282338 354774 282574
rect 354154 264894 354774 282338
rect 354154 264658 354186 264894
rect 354422 264658 354506 264894
rect 354742 264658 354774 264894
rect 354154 264574 354774 264658
rect 354154 264338 354186 264574
rect 354422 264338 354506 264574
rect 354742 264338 354774 264574
rect 354154 246894 354774 264338
rect 354154 246658 354186 246894
rect 354422 246658 354506 246894
rect 354742 246658 354774 246894
rect 354154 246574 354774 246658
rect 354154 246338 354186 246574
rect 354422 246338 354506 246574
rect 354742 246338 354774 246574
rect 354154 228894 354774 246338
rect 354154 228658 354186 228894
rect 354422 228658 354506 228894
rect 354742 228658 354774 228894
rect 354154 228574 354774 228658
rect 354154 228338 354186 228574
rect 354422 228338 354506 228574
rect 354742 228338 354774 228574
rect 354154 210894 354774 228338
rect 354154 210658 354186 210894
rect 354422 210658 354506 210894
rect 354742 210658 354774 210894
rect 354154 210574 354774 210658
rect 354154 210338 354186 210574
rect 354422 210338 354506 210574
rect 354742 210338 354774 210574
rect 354154 192894 354774 210338
rect 354154 192658 354186 192894
rect 354422 192658 354506 192894
rect 354742 192658 354774 192894
rect 354154 192574 354774 192658
rect 354154 192338 354186 192574
rect 354422 192338 354506 192574
rect 354742 192338 354774 192574
rect 354154 174894 354774 192338
rect 354154 174658 354186 174894
rect 354422 174658 354506 174894
rect 354742 174658 354774 174894
rect 354154 174574 354774 174658
rect 354154 174338 354186 174574
rect 354422 174338 354506 174574
rect 354742 174338 354774 174574
rect 354154 156894 354774 174338
rect 354154 156658 354186 156894
rect 354422 156658 354506 156894
rect 354742 156658 354774 156894
rect 354154 156574 354774 156658
rect 354154 156338 354186 156574
rect 354422 156338 354506 156574
rect 354742 156338 354774 156574
rect 354154 138894 354774 156338
rect 354154 138658 354186 138894
rect 354422 138658 354506 138894
rect 354742 138658 354774 138894
rect 354154 138574 354774 138658
rect 354154 138338 354186 138574
rect 354422 138338 354506 138574
rect 354742 138338 354774 138574
rect 354154 120894 354774 138338
rect 354154 120658 354186 120894
rect 354422 120658 354506 120894
rect 354742 120658 354774 120894
rect 354154 120574 354774 120658
rect 354154 120338 354186 120574
rect 354422 120338 354506 120574
rect 354742 120338 354774 120574
rect 354154 102894 354774 120338
rect 354154 102658 354186 102894
rect 354422 102658 354506 102894
rect 354742 102658 354774 102894
rect 354154 102574 354774 102658
rect 354154 102338 354186 102574
rect 354422 102338 354506 102574
rect 354742 102338 354774 102574
rect 354154 84894 354774 102338
rect 354154 84658 354186 84894
rect 354422 84658 354506 84894
rect 354742 84658 354774 84894
rect 354154 84574 354774 84658
rect 354154 84338 354186 84574
rect 354422 84338 354506 84574
rect 354742 84338 354774 84574
rect 354154 66894 354774 84338
rect 354154 66658 354186 66894
rect 354422 66658 354506 66894
rect 354742 66658 354774 66894
rect 354154 66574 354774 66658
rect 354154 66338 354186 66574
rect 354422 66338 354506 66574
rect 354742 66338 354774 66574
rect 354154 48894 354774 66338
rect 354154 48658 354186 48894
rect 354422 48658 354506 48894
rect 354742 48658 354774 48894
rect 354154 48574 354774 48658
rect 354154 48338 354186 48574
rect 354422 48338 354506 48574
rect 354742 48338 354774 48574
rect 354154 30894 354774 48338
rect 354154 30658 354186 30894
rect 354422 30658 354506 30894
rect 354742 30658 354774 30894
rect 354154 30574 354774 30658
rect 354154 30338 354186 30574
rect 354422 30338 354506 30574
rect 354742 30338 354774 30574
rect 354154 12894 354774 30338
rect 354154 12658 354186 12894
rect 354422 12658 354506 12894
rect 354742 12658 354774 12894
rect 354154 12574 354774 12658
rect 354154 12338 354186 12574
rect 354422 12338 354506 12574
rect 354742 12338 354774 12574
rect 354154 -2776 354774 12338
rect 354154 -3012 354186 -2776
rect 354422 -3012 354506 -2776
rect 354742 -3012 354774 -2776
rect 354154 -3096 354774 -3012
rect 354154 -3332 354186 -3096
rect 354422 -3332 354506 -3096
rect 354742 -3332 354774 -3096
rect 354154 -4324 354774 -3332
rect 357874 463972 358494 464004
rect 357874 463736 357906 463972
rect 358142 463736 358226 463972
rect 358462 463736 358494 463972
rect 357874 463652 358494 463736
rect 357874 463416 357906 463652
rect 358142 463416 358226 463652
rect 358462 463416 358494 463652
rect 357874 448614 358494 463416
rect 357874 448378 357906 448614
rect 358142 448378 358226 448614
rect 358462 448378 358494 448614
rect 357874 448294 358494 448378
rect 357874 448058 357906 448294
rect 358142 448058 358226 448294
rect 358462 448058 358494 448294
rect 357874 430614 358494 448058
rect 357874 430378 357906 430614
rect 358142 430378 358226 430614
rect 358462 430378 358494 430614
rect 357874 430294 358494 430378
rect 357874 430058 357906 430294
rect 358142 430058 358226 430294
rect 358462 430058 358494 430294
rect 357874 412614 358494 430058
rect 357874 412378 357906 412614
rect 358142 412378 358226 412614
rect 358462 412378 358494 412614
rect 357874 412294 358494 412378
rect 357874 412058 357906 412294
rect 358142 412058 358226 412294
rect 358462 412058 358494 412294
rect 357874 394614 358494 412058
rect 357874 394378 357906 394614
rect 358142 394378 358226 394614
rect 358462 394378 358494 394614
rect 357874 394294 358494 394378
rect 357874 394058 357906 394294
rect 358142 394058 358226 394294
rect 358462 394058 358494 394294
rect 357874 376614 358494 394058
rect 357874 376378 357906 376614
rect 358142 376378 358226 376614
rect 358462 376378 358494 376614
rect 357874 376294 358494 376378
rect 357874 376058 357906 376294
rect 358142 376058 358226 376294
rect 358462 376058 358494 376294
rect 357874 358614 358494 376058
rect 357874 358378 357906 358614
rect 358142 358378 358226 358614
rect 358462 358378 358494 358614
rect 357874 358294 358494 358378
rect 357874 358058 357906 358294
rect 358142 358058 358226 358294
rect 358462 358058 358494 358294
rect 357874 340614 358494 358058
rect 357874 340378 357906 340614
rect 358142 340378 358226 340614
rect 358462 340378 358494 340614
rect 357874 340294 358494 340378
rect 357874 340058 357906 340294
rect 358142 340058 358226 340294
rect 358462 340058 358494 340294
rect 357874 322614 358494 340058
rect 357874 322378 357906 322614
rect 358142 322378 358226 322614
rect 358462 322378 358494 322614
rect 357874 322294 358494 322378
rect 357874 322058 357906 322294
rect 358142 322058 358226 322294
rect 358462 322058 358494 322294
rect 357874 304614 358494 322058
rect 357874 304378 357906 304614
rect 358142 304378 358226 304614
rect 358462 304378 358494 304614
rect 357874 304294 358494 304378
rect 357874 304058 357906 304294
rect 358142 304058 358226 304294
rect 358462 304058 358494 304294
rect 357874 286614 358494 304058
rect 357874 286378 357906 286614
rect 358142 286378 358226 286614
rect 358462 286378 358494 286614
rect 357874 286294 358494 286378
rect 357874 286058 357906 286294
rect 358142 286058 358226 286294
rect 358462 286058 358494 286294
rect 357874 268614 358494 286058
rect 357874 268378 357906 268614
rect 358142 268378 358226 268614
rect 358462 268378 358494 268614
rect 357874 268294 358494 268378
rect 357874 268058 357906 268294
rect 358142 268058 358226 268294
rect 358462 268058 358494 268294
rect 357874 250614 358494 268058
rect 357874 250378 357906 250614
rect 358142 250378 358226 250614
rect 358462 250378 358494 250614
rect 357874 250294 358494 250378
rect 357874 250058 357906 250294
rect 358142 250058 358226 250294
rect 358462 250058 358494 250294
rect 357874 232614 358494 250058
rect 357874 232378 357906 232614
rect 358142 232378 358226 232614
rect 358462 232378 358494 232614
rect 357874 232294 358494 232378
rect 357874 232058 357906 232294
rect 358142 232058 358226 232294
rect 358462 232058 358494 232294
rect 357874 214614 358494 232058
rect 357874 214378 357906 214614
rect 358142 214378 358226 214614
rect 358462 214378 358494 214614
rect 357874 214294 358494 214378
rect 357874 214058 357906 214294
rect 358142 214058 358226 214294
rect 358462 214058 358494 214294
rect 357874 196614 358494 214058
rect 357874 196378 357906 196614
rect 358142 196378 358226 196614
rect 358462 196378 358494 196614
rect 357874 196294 358494 196378
rect 357874 196058 357906 196294
rect 358142 196058 358226 196294
rect 358462 196058 358494 196294
rect 357874 178614 358494 196058
rect 357874 178378 357906 178614
rect 358142 178378 358226 178614
rect 358462 178378 358494 178614
rect 357874 178294 358494 178378
rect 357874 178058 357906 178294
rect 358142 178058 358226 178294
rect 358462 178058 358494 178294
rect 357874 160614 358494 178058
rect 357874 160378 357906 160614
rect 358142 160378 358226 160614
rect 358462 160378 358494 160614
rect 357874 160294 358494 160378
rect 357874 160058 357906 160294
rect 358142 160058 358226 160294
rect 358462 160058 358494 160294
rect 357874 142614 358494 160058
rect 357874 142378 357906 142614
rect 358142 142378 358226 142614
rect 358462 142378 358494 142614
rect 357874 142294 358494 142378
rect 357874 142058 357906 142294
rect 358142 142058 358226 142294
rect 358462 142058 358494 142294
rect 357874 124614 358494 142058
rect 357874 124378 357906 124614
rect 358142 124378 358226 124614
rect 358462 124378 358494 124614
rect 357874 124294 358494 124378
rect 357874 124058 357906 124294
rect 358142 124058 358226 124294
rect 358462 124058 358494 124294
rect 357874 106614 358494 124058
rect 357874 106378 357906 106614
rect 358142 106378 358226 106614
rect 358462 106378 358494 106614
rect 357874 106294 358494 106378
rect 357874 106058 357906 106294
rect 358142 106058 358226 106294
rect 358462 106058 358494 106294
rect 357874 88614 358494 106058
rect 357874 88378 357906 88614
rect 358142 88378 358226 88614
rect 358462 88378 358494 88614
rect 357874 88294 358494 88378
rect 357874 88058 357906 88294
rect 358142 88058 358226 88294
rect 358462 88058 358494 88294
rect 357874 70614 358494 88058
rect 357874 70378 357906 70614
rect 358142 70378 358226 70614
rect 358462 70378 358494 70614
rect 357874 70294 358494 70378
rect 357874 70058 357906 70294
rect 358142 70058 358226 70294
rect 358462 70058 358494 70294
rect 357874 52614 358494 70058
rect 357874 52378 357906 52614
rect 358142 52378 358226 52614
rect 358462 52378 358494 52614
rect 357874 52294 358494 52378
rect 357874 52058 357906 52294
rect 358142 52058 358226 52294
rect 358462 52058 358494 52294
rect 357874 34614 358494 52058
rect 357874 34378 357906 34614
rect 358142 34378 358226 34614
rect 358462 34378 358494 34614
rect 357874 34294 358494 34378
rect 357874 34058 357906 34294
rect 358142 34058 358226 34294
rect 358462 34058 358494 34294
rect 357874 16614 358494 34058
rect 357874 16378 357906 16614
rect 358142 16378 358226 16614
rect 358462 16378 358494 16614
rect 357874 16294 358494 16378
rect 357874 16058 357906 16294
rect 358142 16058 358226 16294
rect 358462 16058 358494 16294
rect 357874 -3736 358494 16058
rect 357874 -3972 357906 -3736
rect 358142 -3972 358226 -3736
rect 358462 -3972 358494 -3736
rect 357874 -4056 358494 -3972
rect 357874 -4292 357906 -4056
rect 358142 -4292 358226 -4056
rect 358462 -4292 358494 -4056
rect 357874 -4324 358494 -4292
rect 364714 461092 365334 464004
rect 364714 460856 364746 461092
rect 364982 460856 365066 461092
rect 365302 460856 365334 461092
rect 364714 460772 365334 460856
rect 364714 460536 364746 460772
rect 364982 460536 365066 460772
rect 365302 460536 365334 460772
rect 364714 455454 365334 460536
rect 364714 455218 364746 455454
rect 364982 455218 365066 455454
rect 365302 455218 365334 455454
rect 364714 455134 365334 455218
rect 364714 454898 364746 455134
rect 364982 454898 365066 455134
rect 365302 454898 365334 455134
rect 364714 437454 365334 454898
rect 364714 437218 364746 437454
rect 364982 437218 365066 437454
rect 365302 437218 365334 437454
rect 364714 437134 365334 437218
rect 364714 436898 364746 437134
rect 364982 436898 365066 437134
rect 365302 436898 365334 437134
rect 364714 419454 365334 436898
rect 364714 419218 364746 419454
rect 364982 419218 365066 419454
rect 365302 419218 365334 419454
rect 364714 419134 365334 419218
rect 364714 418898 364746 419134
rect 364982 418898 365066 419134
rect 365302 418898 365334 419134
rect 364714 401454 365334 418898
rect 364714 401218 364746 401454
rect 364982 401218 365066 401454
rect 365302 401218 365334 401454
rect 364714 401134 365334 401218
rect 364714 400898 364746 401134
rect 364982 400898 365066 401134
rect 365302 400898 365334 401134
rect 364714 383454 365334 400898
rect 364714 383218 364746 383454
rect 364982 383218 365066 383454
rect 365302 383218 365334 383454
rect 364714 383134 365334 383218
rect 364714 382898 364746 383134
rect 364982 382898 365066 383134
rect 365302 382898 365334 383134
rect 364714 365454 365334 382898
rect 364714 365218 364746 365454
rect 364982 365218 365066 365454
rect 365302 365218 365334 365454
rect 364714 365134 365334 365218
rect 364714 364898 364746 365134
rect 364982 364898 365066 365134
rect 365302 364898 365334 365134
rect 364714 347454 365334 364898
rect 364714 347218 364746 347454
rect 364982 347218 365066 347454
rect 365302 347218 365334 347454
rect 364714 347134 365334 347218
rect 364714 346898 364746 347134
rect 364982 346898 365066 347134
rect 365302 346898 365334 347134
rect 364714 329454 365334 346898
rect 364714 329218 364746 329454
rect 364982 329218 365066 329454
rect 365302 329218 365334 329454
rect 364714 329134 365334 329218
rect 364714 328898 364746 329134
rect 364982 328898 365066 329134
rect 365302 328898 365334 329134
rect 364714 311454 365334 328898
rect 364714 311218 364746 311454
rect 364982 311218 365066 311454
rect 365302 311218 365334 311454
rect 364714 311134 365334 311218
rect 364714 310898 364746 311134
rect 364982 310898 365066 311134
rect 365302 310898 365334 311134
rect 364714 293454 365334 310898
rect 364714 293218 364746 293454
rect 364982 293218 365066 293454
rect 365302 293218 365334 293454
rect 364714 293134 365334 293218
rect 364714 292898 364746 293134
rect 364982 292898 365066 293134
rect 365302 292898 365334 293134
rect 364714 275454 365334 292898
rect 364714 275218 364746 275454
rect 364982 275218 365066 275454
rect 365302 275218 365334 275454
rect 364714 275134 365334 275218
rect 364714 274898 364746 275134
rect 364982 274898 365066 275134
rect 365302 274898 365334 275134
rect 364714 257454 365334 274898
rect 364714 257218 364746 257454
rect 364982 257218 365066 257454
rect 365302 257218 365334 257454
rect 364714 257134 365334 257218
rect 364714 256898 364746 257134
rect 364982 256898 365066 257134
rect 365302 256898 365334 257134
rect 364714 239454 365334 256898
rect 364714 239218 364746 239454
rect 364982 239218 365066 239454
rect 365302 239218 365334 239454
rect 364714 239134 365334 239218
rect 364714 238898 364746 239134
rect 364982 238898 365066 239134
rect 365302 238898 365334 239134
rect 364714 221454 365334 238898
rect 364714 221218 364746 221454
rect 364982 221218 365066 221454
rect 365302 221218 365334 221454
rect 364714 221134 365334 221218
rect 364714 220898 364746 221134
rect 364982 220898 365066 221134
rect 365302 220898 365334 221134
rect 364714 203454 365334 220898
rect 364714 203218 364746 203454
rect 364982 203218 365066 203454
rect 365302 203218 365334 203454
rect 364714 203134 365334 203218
rect 364714 202898 364746 203134
rect 364982 202898 365066 203134
rect 365302 202898 365334 203134
rect 364714 185454 365334 202898
rect 364714 185218 364746 185454
rect 364982 185218 365066 185454
rect 365302 185218 365334 185454
rect 364714 185134 365334 185218
rect 364714 184898 364746 185134
rect 364982 184898 365066 185134
rect 365302 184898 365334 185134
rect 364714 167454 365334 184898
rect 364714 167218 364746 167454
rect 364982 167218 365066 167454
rect 365302 167218 365334 167454
rect 364714 167134 365334 167218
rect 364714 166898 364746 167134
rect 364982 166898 365066 167134
rect 365302 166898 365334 167134
rect 364714 149454 365334 166898
rect 364714 149218 364746 149454
rect 364982 149218 365066 149454
rect 365302 149218 365334 149454
rect 364714 149134 365334 149218
rect 364714 148898 364746 149134
rect 364982 148898 365066 149134
rect 365302 148898 365334 149134
rect 364714 131454 365334 148898
rect 364714 131218 364746 131454
rect 364982 131218 365066 131454
rect 365302 131218 365334 131454
rect 364714 131134 365334 131218
rect 364714 130898 364746 131134
rect 364982 130898 365066 131134
rect 365302 130898 365334 131134
rect 364714 113454 365334 130898
rect 364714 113218 364746 113454
rect 364982 113218 365066 113454
rect 365302 113218 365334 113454
rect 364714 113134 365334 113218
rect 364714 112898 364746 113134
rect 364982 112898 365066 113134
rect 365302 112898 365334 113134
rect 364714 95454 365334 112898
rect 364714 95218 364746 95454
rect 364982 95218 365066 95454
rect 365302 95218 365334 95454
rect 364714 95134 365334 95218
rect 364714 94898 364746 95134
rect 364982 94898 365066 95134
rect 365302 94898 365334 95134
rect 364714 77454 365334 94898
rect 364714 77218 364746 77454
rect 364982 77218 365066 77454
rect 365302 77218 365334 77454
rect 364714 77134 365334 77218
rect 364714 76898 364746 77134
rect 364982 76898 365066 77134
rect 365302 76898 365334 77134
rect 364714 59454 365334 76898
rect 364714 59218 364746 59454
rect 364982 59218 365066 59454
rect 365302 59218 365334 59454
rect 364714 59134 365334 59218
rect 364714 58898 364746 59134
rect 364982 58898 365066 59134
rect 365302 58898 365334 59134
rect 364714 41454 365334 58898
rect 364714 41218 364746 41454
rect 364982 41218 365066 41454
rect 365302 41218 365334 41454
rect 364714 41134 365334 41218
rect 364714 40898 364746 41134
rect 364982 40898 365066 41134
rect 365302 40898 365334 41134
rect 364714 23454 365334 40898
rect 364714 23218 364746 23454
rect 364982 23218 365066 23454
rect 365302 23218 365334 23454
rect 364714 23134 365334 23218
rect 364714 22898 364746 23134
rect 364982 22898 365066 23134
rect 365302 22898 365334 23134
rect 364714 5454 365334 22898
rect 364714 5218 364746 5454
rect 364982 5218 365066 5454
rect 365302 5218 365334 5454
rect 364714 5134 365334 5218
rect 364714 4898 364746 5134
rect 364982 4898 365066 5134
rect 365302 4898 365334 5134
rect 364714 -856 365334 4898
rect 364714 -1092 364746 -856
rect 364982 -1092 365066 -856
rect 365302 -1092 365334 -856
rect 364714 -1176 365334 -1092
rect 364714 -1412 364746 -1176
rect 364982 -1412 365066 -1176
rect 365302 -1412 365334 -1176
rect 364714 -4324 365334 -1412
rect 368434 462052 369054 464004
rect 368434 461816 368466 462052
rect 368702 461816 368786 462052
rect 369022 461816 369054 462052
rect 368434 461732 369054 461816
rect 368434 461496 368466 461732
rect 368702 461496 368786 461732
rect 369022 461496 369054 461732
rect 368434 441174 369054 461496
rect 368434 440938 368466 441174
rect 368702 440938 368786 441174
rect 369022 440938 369054 441174
rect 368434 440854 369054 440938
rect 368434 440618 368466 440854
rect 368702 440618 368786 440854
rect 369022 440618 369054 440854
rect 368434 423174 369054 440618
rect 368434 422938 368466 423174
rect 368702 422938 368786 423174
rect 369022 422938 369054 423174
rect 368434 422854 369054 422938
rect 368434 422618 368466 422854
rect 368702 422618 368786 422854
rect 369022 422618 369054 422854
rect 368434 405174 369054 422618
rect 368434 404938 368466 405174
rect 368702 404938 368786 405174
rect 369022 404938 369054 405174
rect 368434 404854 369054 404938
rect 368434 404618 368466 404854
rect 368702 404618 368786 404854
rect 369022 404618 369054 404854
rect 368434 387174 369054 404618
rect 368434 386938 368466 387174
rect 368702 386938 368786 387174
rect 369022 386938 369054 387174
rect 368434 386854 369054 386938
rect 368434 386618 368466 386854
rect 368702 386618 368786 386854
rect 369022 386618 369054 386854
rect 368434 369174 369054 386618
rect 368434 368938 368466 369174
rect 368702 368938 368786 369174
rect 369022 368938 369054 369174
rect 368434 368854 369054 368938
rect 368434 368618 368466 368854
rect 368702 368618 368786 368854
rect 369022 368618 369054 368854
rect 368434 351174 369054 368618
rect 368434 350938 368466 351174
rect 368702 350938 368786 351174
rect 369022 350938 369054 351174
rect 368434 350854 369054 350938
rect 368434 350618 368466 350854
rect 368702 350618 368786 350854
rect 369022 350618 369054 350854
rect 368434 333174 369054 350618
rect 368434 332938 368466 333174
rect 368702 332938 368786 333174
rect 369022 332938 369054 333174
rect 368434 332854 369054 332938
rect 368434 332618 368466 332854
rect 368702 332618 368786 332854
rect 369022 332618 369054 332854
rect 368434 315174 369054 332618
rect 368434 314938 368466 315174
rect 368702 314938 368786 315174
rect 369022 314938 369054 315174
rect 368434 314854 369054 314938
rect 368434 314618 368466 314854
rect 368702 314618 368786 314854
rect 369022 314618 369054 314854
rect 368434 297174 369054 314618
rect 368434 296938 368466 297174
rect 368702 296938 368786 297174
rect 369022 296938 369054 297174
rect 368434 296854 369054 296938
rect 368434 296618 368466 296854
rect 368702 296618 368786 296854
rect 369022 296618 369054 296854
rect 368434 279174 369054 296618
rect 368434 278938 368466 279174
rect 368702 278938 368786 279174
rect 369022 278938 369054 279174
rect 368434 278854 369054 278938
rect 368434 278618 368466 278854
rect 368702 278618 368786 278854
rect 369022 278618 369054 278854
rect 368434 261174 369054 278618
rect 368434 260938 368466 261174
rect 368702 260938 368786 261174
rect 369022 260938 369054 261174
rect 368434 260854 369054 260938
rect 368434 260618 368466 260854
rect 368702 260618 368786 260854
rect 369022 260618 369054 260854
rect 368434 243174 369054 260618
rect 368434 242938 368466 243174
rect 368702 242938 368786 243174
rect 369022 242938 369054 243174
rect 368434 242854 369054 242938
rect 368434 242618 368466 242854
rect 368702 242618 368786 242854
rect 369022 242618 369054 242854
rect 368434 225174 369054 242618
rect 368434 224938 368466 225174
rect 368702 224938 368786 225174
rect 369022 224938 369054 225174
rect 368434 224854 369054 224938
rect 368434 224618 368466 224854
rect 368702 224618 368786 224854
rect 369022 224618 369054 224854
rect 368434 207174 369054 224618
rect 368434 206938 368466 207174
rect 368702 206938 368786 207174
rect 369022 206938 369054 207174
rect 368434 206854 369054 206938
rect 368434 206618 368466 206854
rect 368702 206618 368786 206854
rect 369022 206618 369054 206854
rect 368434 189174 369054 206618
rect 368434 188938 368466 189174
rect 368702 188938 368786 189174
rect 369022 188938 369054 189174
rect 368434 188854 369054 188938
rect 368434 188618 368466 188854
rect 368702 188618 368786 188854
rect 369022 188618 369054 188854
rect 368434 171174 369054 188618
rect 368434 170938 368466 171174
rect 368702 170938 368786 171174
rect 369022 170938 369054 171174
rect 368434 170854 369054 170938
rect 368434 170618 368466 170854
rect 368702 170618 368786 170854
rect 369022 170618 369054 170854
rect 368434 153174 369054 170618
rect 368434 152938 368466 153174
rect 368702 152938 368786 153174
rect 369022 152938 369054 153174
rect 368434 152854 369054 152938
rect 368434 152618 368466 152854
rect 368702 152618 368786 152854
rect 369022 152618 369054 152854
rect 368434 135174 369054 152618
rect 368434 134938 368466 135174
rect 368702 134938 368786 135174
rect 369022 134938 369054 135174
rect 368434 134854 369054 134938
rect 368434 134618 368466 134854
rect 368702 134618 368786 134854
rect 369022 134618 369054 134854
rect 368434 117174 369054 134618
rect 368434 116938 368466 117174
rect 368702 116938 368786 117174
rect 369022 116938 369054 117174
rect 368434 116854 369054 116938
rect 368434 116618 368466 116854
rect 368702 116618 368786 116854
rect 369022 116618 369054 116854
rect 368434 99174 369054 116618
rect 368434 98938 368466 99174
rect 368702 98938 368786 99174
rect 369022 98938 369054 99174
rect 368434 98854 369054 98938
rect 368434 98618 368466 98854
rect 368702 98618 368786 98854
rect 369022 98618 369054 98854
rect 368434 81174 369054 98618
rect 368434 80938 368466 81174
rect 368702 80938 368786 81174
rect 369022 80938 369054 81174
rect 368434 80854 369054 80938
rect 368434 80618 368466 80854
rect 368702 80618 368786 80854
rect 369022 80618 369054 80854
rect 368434 63174 369054 80618
rect 368434 62938 368466 63174
rect 368702 62938 368786 63174
rect 369022 62938 369054 63174
rect 368434 62854 369054 62938
rect 368434 62618 368466 62854
rect 368702 62618 368786 62854
rect 369022 62618 369054 62854
rect 368434 45174 369054 62618
rect 368434 44938 368466 45174
rect 368702 44938 368786 45174
rect 369022 44938 369054 45174
rect 368434 44854 369054 44938
rect 368434 44618 368466 44854
rect 368702 44618 368786 44854
rect 369022 44618 369054 44854
rect 368434 27174 369054 44618
rect 368434 26938 368466 27174
rect 368702 26938 368786 27174
rect 369022 26938 369054 27174
rect 368434 26854 369054 26938
rect 368434 26618 368466 26854
rect 368702 26618 368786 26854
rect 369022 26618 369054 26854
rect 368434 9174 369054 26618
rect 368434 8938 368466 9174
rect 368702 8938 368786 9174
rect 369022 8938 369054 9174
rect 368434 8854 369054 8938
rect 368434 8618 368466 8854
rect 368702 8618 368786 8854
rect 369022 8618 369054 8854
rect 368434 -1816 369054 8618
rect 368434 -2052 368466 -1816
rect 368702 -2052 368786 -1816
rect 369022 -2052 369054 -1816
rect 368434 -2136 369054 -2052
rect 368434 -2372 368466 -2136
rect 368702 -2372 368786 -2136
rect 369022 -2372 369054 -2136
rect 368434 -4324 369054 -2372
rect 372154 463012 372774 464004
rect 372154 462776 372186 463012
rect 372422 462776 372506 463012
rect 372742 462776 372774 463012
rect 372154 462692 372774 462776
rect 372154 462456 372186 462692
rect 372422 462456 372506 462692
rect 372742 462456 372774 462692
rect 372154 444894 372774 462456
rect 372154 444658 372186 444894
rect 372422 444658 372506 444894
rect 372742 444658 372774 444894
rect 372154 444574 372774 444658
rect 372154 444338 372186 444574
rect 372422 444338 372506 444574
rect 372742 444338 372774 444574
rect 372154 426894 372774 444338
rect 372154 426658 372186 426894
rect 372422 426658 372506 426894
rect 372742 426658 372774 426894
rect 372154 426574 372774 426658
rect 372154 426338 372186 426574
rect 372422 426338 372506 426574
rect 372742 426338 372774 426574
rect 372154 408894 372774 426338
rect 372154 408658 372186 408894
rect 372422 408658 372506 408894
rect 372742 408658 372774 408894
rect 372154 408574 372774 408658
rect 372154 408338 372186 408574
rect 372422 408338 372506 408574
rect 372742 408338 372774 408574
rect 372154 390894 372774 408338
rect 372154 390658 372186 390894
rect 372422 390658 372506 390894
rect 372742 390658 372774 390894
rect 372154 390574 372774 390658
rect 372154 390338 372186 390574
rect 372422 390338 372506 390574
rect 372742 390338 372774 390574
rect 372154 372894 372774 390338
rect 372154 372658 372186 372894
rect 372422 372658 372506 372894
rect 372742 372658 372774 372894
rect 372154 372574 372774 372658
rect 372154 372338 372186 372574
rect 372422 372338 372506 372574
rect 372742 372338 372774 372574
rect 372154 354894 372774 372338
rect 372154 354658 372186 354894
rect 372422 354658 372506 354894
rect 372742 354658 372774 354894
rect 372154 354574 372774 354658
rect 372154 354338 372186 354574
rect 372422 354338 372506 354574
rect 372742 354338 372774 354574
rect 372154 336894 372774 354338
rect 372154 336658 372186 336894
rect 372422 336658 372506 336894
rect 372742 336658 372774 336894
rect 372154 336574 372774 336658
rect 372154 336338 372186 336574
rect 372422 336338 372506 336574
rect 372742 336338 372774 336574
rect 372154 318894 372774 336338
rect 372154 318658 372186 318894
rect 372422 318658 372506 318894
rect 372742 318658 372774 318894
rect 372154 318574 372774 318658
rect 372154 318338 372186 318574
rect 372422 318338 372506 318574
rect 372742 318338 372774 318574
rect 372154 300894 372774 318338
rect 372154 300658 372186 300894
rect 372422 300658 372506 300894
rect 372742 300658 372774 300894
rect 372154 300574 372774 300658
rect 372154 300338 372186 300574
rect 372422 300338 372506 300574
rect 372742 300338 372774 300574
rect 372154 282894 372774 300338
rect 372154 282658 372186 282894
rect 372422 282658 372506 282894
rect 372742 282658 372774 282894
rect 372154 282574 372774 282658
rect 372154 282338 372186 282574
rect 372422 282338 372506 282574
rect 372742 282338 372774 282574
rect 372154 264894 372774 282338
rect 372154 264658 372186 264894
rect 372422 264658 372506 264894
rect 372742 264658 372774 264894
rect 372154 264574 372774 264658
rect 372154 264338 372186 264574
rect 372422 264338 372506 264574
rect 372742 264338 372774 264574
rect 372154 246894 372774 264338
rect 372154 246658 372186 246894
rect 372422 246658 372506 246894
rect 372742 246658 372774 246894
rect 372154 246574 372774 246658
rect 372154 246338 372186 246574
rect 372422 246338 372506 246574
rect 372742 246338 372774 246574
rect 372154 228894 372774 246338
rect 372154 228658 372186 228894
rect 372422 228658 372506 228894
rect 372742 228658 372774 228894
rect 372154 228574 372774 228658
rect 372154 228338 372186 228574
rect 372422 228338 372506 228574
rect 372742 228338 372774 228574
rect 372154 210894 372774 228338
rect 372154 210658 372186 210894
rect 372422 210658 372506 210894
rect 372742 210658 372774 210894
rect 372154 210574 372774 210658
rect 372154 210338 372186 210574
rect 372422 210338 372506 210574
rect 372742 210338 372774 210574
rect 372154 192894 372774 210338
rect 372154 192658 372186 192894
rect 372422 192658 372506 192894
rect 372742 192658 372774 192894
rect 372154 192574 372774 192658
rect 372154 192338 372186 192574
rect 372422 192338 372506 192574
rect 372742 192338 372774 192574
rect 372154 174894 372774 192338
rect 372154 174658 372186 174894
rect 372422 174658 372506 174894
rect 372742 174658 372774 174894
rect 372154 174574 372774 174658
rect 372154 174338 372186 174574
rect 372422 174338 372506 174574
rect 372742 174338 372774 174574
rect 372154 156894 372774 174338
rect 372154 156658 372186 156894
rect 372422 156658 372506 156894
rect 372742 156658 372774 156894
rect 372154 156574 372774 156658
rect 372154 156338 372186 156574
rect 372422 156338 372506 156574
rect 372742 156338 372774 156574
rect 372154 138894 372774 156338
rect 372154 138658 372186 138894
rect 372422 138658 372506 138894
rect 372742 138658 372774 138894
rect 372154 138574 372774 138658
rect 372154 138338 372186 138574
rect 372422 138338 372506 138574
rect 372742 138338 372774 138574
rect 372154 120894 372774 138338
rect 372154 120658 372186 120894
rect 372422 120658 372506 120894
rect 372742 120658 372774 120894
rect 372154 120574 372774 120658
rect 372154 120338 372186 120574
rect 372422 120338 372506 120574
rect 372742 120338 372774 120574
rect 372154 102894 372774 120338
rect 372154 102658 372186 102894
rect 372422 102658 372506 102894
rect 372742 102658 372774 102894
rect 372154 102574 372774 102658
rect 372154 102338 372186 102574
rect 372422 102338 372506 102574
rect 372742 102338 372774 102574
rect 372154 84894 372774 102338
rect 372154 84658 372186 84894
rect 372422 84658 372506 84894
rect 372742 84658 372774 84894
rect 372154 84574 372774 84658
rect 372154 84338 372186 84574
rect 372422 84338 372506 84574
rect 372742 84338 372774 84574
rect 372154 66894 372774 84338
rect 372154 66658 372186 66894
rect 372422 66658 372506 66894
rect 372742 66658 372774 66894
rect 372154 66574 372774 66658
rect 372154 66338 372186 66574
rect 372422 66338 372506 66574
rect 372742 66338 372774 66574
rect 372154 48894 372774 66338
rect 372154 48658 372186 48894
rect 372422 48658 372506 48894
rect 372742 48658 372774 48894
rect 372154 48574 372774 48658
rect 372154 48338 372186 48574
rect 372422 48338 372506 48574
rect 372742 48338 372774 48574
rect 372154 30894 372774 48338
rect 372154 30658 372186 30894
rect 372422 30658 372506 30894
rect 372742 30658 372774 30894
rect 372154 30574 372774 30658
rect 372154 30338 372186 30574
rect 372422 30338 372506 30574
rect 372742 30338 372774 30574
rect 372154 12894 372774 30338
rect 372154 12658 372186 12894
rect 372422 12658 372506 12894
rect 372742 12658 372774 12894
rect 372154 12574 372774 12658
rect 372154 12338 372186 12574
rect 372422 12338 372506 12574
rect 372742 12338 372774 12574
rect 372154 -2776 372774 12338
rect 372154 -3012 372186 -2776
rect 372422 -3012 372506 -2776
rect 372742 -3012 372774 -2776
rect 372154 -3096 372774 -3012
rect 372154 -3332 372186 -3096
rect 372422 -3332 372506 -3096
rect 372742 -3332 372774 -3096
rect 372154 -4324 372774 -3332
rect 375874 463972 376494 464004
rect 375874 463736 375906 463972
rect 376142 463736 376226 463972
rect 376462 463736 376494 463972
rect 375874 463652 376494 463736
rect 375874 463416 375906 463652
rect 376142 463416 376226 463652
rect 376462 463416 376494 463652
rect 375874 448614 376494 463416
rect 375874 448378 375906 448614
rect 376142 448378 376226 448614
rect 376462 448378 376494 448614
rect 375874 448294 376494 448378
rect 375874 448058 375906 448294
rect 376142 448058 376226 448294
rect 376462 448058 376494 448294
rect 375874 430614 376494 448058
rect 375874 430378 375906 430614
rect 376142 430378 376226 430614
rect 376462 430378 376494 430614
rect 375874 430294 376494 430378
rect 375874 430058 375906 430294
rect 376142 430058 376226 430294
rect 376462 430058 376494 430294
rect 375874 412614 376494 430058
rect 375874 412378 375906 412614
rect 376142 412378 376226 412614
rect 376462 412378 376494 412614
rect 375874 412294 376494 412378
rect 375874 412058 375906 412294
rect 376142 412058 376226 412294
rect 376462 412058 376494 412294
rect 375874 394614 376494 412058
rect 375874 394378 375906 394614
rect 376142 394378 376226 394614
rect 376462 394378 376494 394614
rect 375874 394294 376494 394378
rect 375874 394058 375906 394294
rect 376142 394058 376226 394294
rect 376462 394058 376494 394294
rect 375874 376614 376494 394058
rect 375874 376378 375906 376614
rect 376142 376378 376226 376614
rect 376462 376378 376494 376614
rect 375874 376294 376494 376378
rect 375874 376058 375906 376294
rect 376142 376058 376226 376294
rect 376462 376058 376494 376294
rect 375874 358614 376494 376058
rect 375874 358378 375906 358614
rect 376142 358378 376226 358614
rect 376462 358378 376494 358614
rect 375874 358294 376494 358378
rect 375874 358058 375906 358294
rect 376142 358058 376226 358294
rect 376462 358058 376494 358294
rect 375874 340614 376494 358058
rect 375874 340378 375906 340614
rect 376142 340378 376226 340614
rect 376462 340378 376494 340614
rect 375874 340294 376494 340378
rect 375874 340058 375906 340294
rect 376142 340058 376226 340294
rect 376462 340058 376494 340294
rect 375874 322614 376494 340058
rect 375874 322378 375906 322614
rect 376142 322378 376226 322614
rect 376462 322378 376494 322614
rect 375874 322294 376494 322378
rect 375874 322058 375906 322294
rect 376142 322058 376226 322294
rect 376462 322058 376494 322294
rect 375874 304614 376494 322058
rect 375874 304378 375906 304614
rect 376142 304378 376226 304614
rect 376462 304378 376494 304614
rect 375874 304294 376494 304378
rect 375874 304058 375906 304294
rect 376142 304058 376226 304294
rect 376462 304058 376494 304294
rect 375874 286614 376494 304058
rect 375874 286378 375906 286614
rect 376142 286378 376226 286614
rect 376462 286378 376494 286614
rect 375874 286294 376494 286378
rect 375874 286058 375906 286294
rect 376142 286058 376226 286294
rect 376462 286058 376494 286294
rect 375874 268614 376494 286058
rect 375874 268378 375906 268614
rect 376142 268378 376226 268614
rect 376462 268378 376494 268614
rect 375874 268294 376494 268378
rect 375874 268058 375906 268294
rect 376142 268058 376226 268294
rect 376462 268058 376494 268294
rect 375874 250614 376494 268058
rect 375874 250378 375906 250614
rect 376142 250378 376226 250614
rect 376462 250378 376494 250614
rect 375874 250294 376494 250378
rect 375874 250058 375906 250294
rect 376142 250058 376226 250294
rect 376462 250058 376494 250294
rect 375874 232614 376494 250058
rect 375874 232378 375906 232614
rect 376142 232378 376226 232614
rect 376462 232378 376494 232614
rect 375874 232294 376494 232378
rect 375874 232058 375906 232294
rect 376142 232058 376226 232294
rect 376462 232058 376494 232294
rect 375874 214614 376494 232058
rect 375874 214378 375906 214614
rect 376142 214378 376226 214614
rect 376462 214378 376494 214614
rect 375874 214294 376494 214378
rect 375874 214058 375906 214294
rect 376142 214058 376226 214294
rect 376462 214058 376494 214294
rect 375874 196614 376494 214058
rect 375874 196378 375906 196614
rect 376142 196378 376226 196614
rect 376462 196378 376494 196614
rect 375874 196294 376494 196378
rect 375874 196058 375906 196294
rect 376142 196058 376226 196294
rect 376462 196058 376494 196294
rect 375874 178614 376494 196058
rect 375874 178378 375906 178614
rect 376142 178378 376226 178614
rect 376462 178378 376494 178614
rect 375874 178294 376494 178378
rect 375874 178058 375906 178294
rect 376142 178058 376226 178294
rect 376462 178058 376494 178294
rect 375874 160614 376494 178058
rect 375874 160378 375906 160614
rect 376142 160378 376226 160614
rect 376462 160378 376494 160614
rect 375874 160294 376494 160378
rect 375874 160058 375906 160294
rect 376142 160058 376226 160294
rect 376462 160058 376494 160294
rect 375874 142614 376494 160058
rect 375874 142378 375906 142614
rect 376142 142378 376226 142614
rect 376462 142378 376494 142614
rect 375874 142294 376494 142378
rect 375874 142058 375906 142294
rect 376142 142058 376226 142294
rect 376462 142058 376494 142294
rect 375874 124614 376494 142058
rect 375874 124378 375906 124614
rect 376142 124378 376226 124614
rect 376462 124378 376494 124614
rect 375874 124294 376494 124378
rect 375874 124058 375906 124294
rect 376142 124058 376226 124294
rect 376462 124058 376494 124294
rect 375874 106614 376494 124058
rect 375874 106378 375906 106614
rect 376142 106378 376226 106614
rect 376462 106378 376494 106614
rect 375874 106294 376494 106378
rect 375874 106058 375906 106294
rect 376142 106058 376226 106294
rect 376462 106058 376494 106294
rect 375874 88614 376494 106058
rect 375874 88378 375906 88614
rect 376142 88378 376226 88614
rect 376462 88378 376494 88614
rect 375874 88294 376494 88378
rect 375874 88058 375906 88294
rect 376142 88058 376226 88294
rect 376462 88058 376494 88294
rect 375874 70614 376494 88058
rect 375874 70378 375906 70614
rect 376142 70378 376226 70614
rect 376462 70378 376494 70614
rect 375874 70294 376494 70378
rect 375874 70058 375906 70294
rect 376142 70058 376226 70294
rect 376462 70058 376494 70294
rect 375874 52614 376494 70058
rect 375874 52378 375906 52614
rect 376142 52378 376226 52614
rect 376462 52378 376494 52614
rect 375874 52294 376494 52378
rect 375874 52058 375906 52294
rect 376142 52058 376226 52294
rect 376462 52058 376494 52294
rect 375874 34614 376494 52058
rect 375874 34378 375906 34614
rect 376142 34378 376226 34614
rect 376462 34378 376494 34614
rect 375874 34294 376494 34378
rect 375874 34058 375906 34294
rect 376142 34058 376226 34294
rect 376462 34058 376494 34294
rect 375874 16614 376494 34058
rect 375874 16378 375906 16614
rect 376142 16378 376226 16614
rect 376462 16378 376494 16614
rect 375874 16294 376494 16378
rect 375874 16058 375906 16294
rect 376142 16058 376226 16294
rect 376462 16058 376494 16294
rect 375874 -3736 376494 16058
rect 375874 -3972 375906 -3736
rect 376142 -3972 376226 -3736
rect 376462 -3972 376494 -3736
rect 375874 -4056 376494 -3972
rect 375874 -4292 375906 -4056
rect 376142 -4292 376226 -4056
rect 376462 -4292 376494 -4056
rect 375874 -4324 376494 -4292
rect 382714 461092 383334 464004
rect 382714 460856 382746 461092
rect 382982 460856 383066 461092
rect 383302 460856 383334 461092
rect 382714 460772 383334 460856
rect 382714 460536 382746 460772
rect 382982 460536 383066 460772
rect 383302 460536 383334 460772
rect 382714 455454 383334 460536
rect 382714 455218 382746 455454
rect 382982 455218 383066 455454
rect 383302 455218 383334 455454
rect 382714 455134 383334 455218
rect 382714 454898 382746 455134
rect 382982 454898 383066 455134
rect 383302 454898 383334 455134
rect 382714 437454 383334 454898
rect 382714 437218 382746 437454
rect 382982 437218 383066 437454
rect 383302 437218 383334 437454
rect 382714 437134 383334 437218
rect 382714 436898 382746 437134
rect 382982 436898 383066 437134
rect 383302 436898 383334 437134
rect 382714 419454 383334 436898
rect 382714 419218 382746 419454
rect 382982 419218 383066 419454
rect 383302 419218 383334 419454
rect 382714 419134 383334 419218
rect 382714 418898 382746 419134
rect 382982 418898 383066 419134
rect 383302 418898 383334 419134
rect 382714 401454 383334 418898
rect 382714 401218 382746 401454
rect 382982 401218 383066 401454
rect 383302 401218 383334 401454
rect 382714 401134 383334 401218
rect 382714 400898 382746 401134
rect 382982 400898 383066 401134
rect 383302 400898 383334 401134
rect 382714 383454 383334 400898
rect 382714 383218 382746 383454
rect 382982 383218 383066 383454
rect 383302 383218 383334 383454
rect 382714 383134 383334 383218
rect 382714 382898 382746 383134
rect 382982 382898 383066 383134
rect 383302 382898 383334 383134
rect 382714 365454 383334 382898
rect 382714 365218 382746 365454
rect 382982 365218 383066 365454
rect 383302 365218 383334 365454
rect 382714 365134 383334 365218
rect 382714 364898 382746 365134
rect 382982 364898 383066 365134
rect 383302 364898 383334 365134
rect 382714 347454 383334 364898
rect 382714 347218 382746 347454
rect 382982 347218 383066 347454
rect 383302 347218 383334 347454
rect 382714 347134 383334 347218
rect 382714 346898 382746 347134
rect 382982 346898 383066 347134
rect 383302 346898 383334 347134
rect 382714 329454 383334 346898
rect 382714 329218 382746 329454
rect 382982 329218 383066 329454
rect 383302 329218 383334 329454
rect 382714 329134 383334 329218
rect 382714 328898 382746 329134
rect 382982 328898 383066 329134
rect 383302 328898 383334 329134
rect 382714 311454 383334 328898
rect 382714 311218 382746 311454
rect 382982 311218 383066 311454
rect 383302 311218 383334 311454
rect 382714 311134 383334 311218
rect 382714 310898 382746 311134
rect 382982 310898 383066 311134
rect 383302 310898 383334 311134
rect 382714 293454 383334 310898
rect 382714 293218 382746 293454
rect 382982 293218 383066 293454
rect 383302 293218 383334 293454
rect 382714 293134 383334 293218
rect 382714 292898 382746 293134
rect 382982 292898 383066 293134
rect 383302 292898 383334 293134
rect 382714 275454 383334 292898
rect 382714 275218 382746 275454
rect 382982 275218 383066 275454
rect 383302 275218 383334 275454
rect 382714 275134 383334 275218
rect 382714 274898 382746 275134
rect 382982 274898 383066 275134
rect 383302 274898 383334 275134
rect 382714 257454 383334 274898
rect 382714 257218 382746 257454
rect 382982 257218 383066 257454
rect 383302 257218 383334 257454
rect 382714 257134 383334 257218
rect 382714 256898 382746 257134
rect 382982 256898 383066 257134
rect 383302 256898 383334 257134
rect 382714 239454 383334 256898
rect 382714 239218 382746 239454
rect 382982 239218 383066 239454
rect 383302 239218 383334 239454
rect 382714 239134 383334 239218
rect 382714 238898 382746 239134
rect 382982 238898 383066 239134
rect 383302 238898 383334 239134
rect 382714 221454 383334 238898
rect 382714 221218 382746 221454
rect 382982 221218 383066 221454
rect 383302 221218 383334 221454
rect 382714 221134 383334 221218
rect 382714 220898 382746 221134
rect 382982 220898 383066 221134
rect 383302 220898 383334 221134
rect 382714 203454 383334 220898
rect 382714 203218 382746 203454
rect 382982 203218 383066 203454
rect 383302 203218 383334 203454
rect 382714 203134 383334 203218
rect 382714 202898 382746 203134
rect 382982 202898 383066 203134
rect 383302 202898 383334 203134
rect 382714 185454 383334 202898
rect 382714 185218 382746 185454
rect 382982 185218 383066 185454
rect 383302 185218 383334 185454
rect 382714 185134 383334 185218
rect 382714 184898 382746 185134
rect 382982 184898 383066 185134
rect 383302 184898 383334 185134
rect 382714 167454 383334 184898
rect 382714 167218 382746 167454
rect 382982 167218 383066 167454
rect 383302 167218 383334 167454
rect 382714 167134 383334 167218
rect 382714 166898 382746 167134
rect 382982 166898 383066 167134
rect 383302 166898 383334 167134
rect 382714 149454 383334 166898
rect 382714 149218 382746 149454
rect 382982 149218 383066 149454
rect 383302 149218 383334 149454
rect 382714 149134 383334 149218
rect 382714 148898 382746 149134
rect 382982 148898 383066 149134
rect 383302 148898 383334 149134
rect 382714 131454 383334 148898
rect 382714 131218 382746 131454
rect 382982 131218 383066 131454
rect 383302 131218 383334 131454
rect 382714 131134 383334 131218
rect 382714 130898 382746 131134
rect 382982 130898 383066 131134
rect 383302 130898 383334 131134
rect 382714 113454 383334 130898
rect 382714 113218 382746 113454
rect 382982 113218 383066 113454
rect 383302 113218 383334 113454
rect 382714 113134 383334 113218
rect 382714 112898 382746 113134
rect 382982 112898 383066 113134
rect 383302 112898 383334 113134
rect 382714 95454 383334 112898
rect 382714 95218 382746 95454
rect 382982 95218 383066 95454
rect 383302 95218 383334 95454
rect 382714 95134 383334 95218
rect 382714 94898 382746 95134
rect 382982 94898 383066 95134
rect 383302 94898 383334 95134
rect 382714 77454 383334 94898
rect 382714 77218 382746 77454
rect 382982 77218 383066 77454
rect 383302 77218 383334 77454
rect 382714 77134 383334 77218
rect 382714 76898 382746 77134
rect 382982 76898 383066 77134
rect 383302 76898 383334 77134
rect 382714 59454 383334 76898
rect 382714 59218 382746 59454
rect 382982 59218 383066 59454
rect 383302 59218 383334 59454
rect 382714 59134 383334 59218
rect 382714 58898 382746 59134
rect 382982 58898 383066 59134
rect 383302 58898 383334 59134
rect 382714 41454 383334 58898
rect 382714 41218 382746 41454
rect 382982 41218 383066 41454
rect 383302 41218 383334 41454
rect 382714 41134 383334 41218
rect 382714 40898 382746 41134
rect 382982 40898 383066 41134
rect 383302 40898 383334 41134
rect 382714 23454 383334 40898
rect 382714 23218 382746 23454
rect 382982 23218 383066 23454
rect 383302 23218 383334 23454
rect 382714 23134 383334 23218
rect 382714 22898 382746 23134
rect 382982 22898 383066 23134
rect 383302 22898 383334 23134
rect 382714 5454 383334 22898
rect 382714 5218 382746 5454
rect 382982 5218 383066 5454
rect 383302 5218 383334 5454
rect 382714 5134 383334 5218
rect 382714 4898 382746 5134
rect 382982 4898 383066 5134
rect 383302 4898 383334 5134
rect 382714 -856 383334 4898
rect 382714 -1092 382746 -856
rect 382982 -1092 383066 -856
rect 383302 -1092 383334 -856
rect 382714 -1176 383334 -1092
rect 382714 -1412 382746 -1176
rect 382982 -1412 383066 -1176
rect 383302 -1412 383334 -1176
rect 382714 -4324 383334 -1412
rect 386434 462052 387054 464004
rect 386434 461816 386466 462052
rect 386702 461816 386786 462052
rect 387022 461816 387054 462052
rect 386434 461732 387054 461816
rect 386434 461496 386466 461732
rect 386702 461496 386786 461732
rect 387022 461496 387054 461732
rect 386434 441174 387054 461496
rect 386434 440938 386466 441174
rect 386702 440938 386786 441174
rect 387022 440938 387054 441174
rect 386434 440854 387054 440938
rect 386434 440618 386466 440854
rect 386702 440618 386786 440854
rect 387022 440618 387054 440854
rect 386434 423174 387054 440618
rect 386434 422938 386466 423174
rect 386702 422938 386786 423174
rect 387022 422938 387054 423174
rect 386434 422854 387054 422938
rect 386434 422618 386466 422854
rect 386702 422618 386786 422854
rect 387022 422618 387054 422854
rect 386434 405174 387054 422618
rect 386434 404938 386466 405174
rect 386702 404938 386786 405174
rect 387022 404938 387054 405174
rect 386434 404854 387054 404938
rect 386434 404618 386466 404854
rect 386702 404618 386786 404854
rect 387022 404618 387054 404854
rect 386434 387174 387054 404618
rect 386434 386938 386466 387174
rect 386702 386938 386786 387174
rect 387022 386938 387054 387174
rect 386434 386854 387054 386938
rect 386434 386618 386466 386854
rect 386702 386618 386786 386854
rect 387022 386618 387054 386854
rect 386434 369174 387054 386618
rect 386434 368938 386466 369174
rect 386702 368938 386786 369174
rect 387022 368938 387054 369174
rect 386434 368854 387054 368938
rect 386434 368618 386466 368854
rect 386702 368618 386786 368854
rect 387022 368618 387054 368854
rect 386434 351174 387054 368618
rect 386434 350938 386466 351174
rect 386702 350938 386786 351174
rect 387022 350938 387054 351174
rect 386434 350854 387054 350938
rect 386434 350618 386466 350854
rect 386702 350618 386786 350854
rect 387022 350618 387054 350854
rect 386434 333174 387054 350618
rect 386434 332938 386466 333174
rect 386702 332938 386786 333174
rect 387022 332938 387054 333174
rect 386434 332854 387054 332938
rect 386434 332618 386466 332854
rect 386702 332618 386786 332854
rect 387022 332618 387054 332854
rect 386434 315174 387054 332618
rect 386434 314938 386466 315174
rect 386702 314938 386786 315174
rect 387022 314938 387054 315174
rect 386434 314854 387054 314938
rect 386434 314618 386466 314854
rect 386702 314618 386786 314854
rect 387022 314618 387054 314854
rect 386434 297174 387054 314618
rect 386434 296938 386466 297174
rect 386702 296938 386786 297174
rect 387022 296938 387054 297174
rect 386434 296854 387054 296938
rect 386434 296618 386466 296854
rect 386702 296618 386786 296854
rect 387022 296618 387054 296854
rect 386434 279174 387054 296618
rect 386434 278938 386466 279174
rect 386702 278938 386786 279174
rect 387022 278938 387054 279174
rect 386434 278854 387054 278938
rect 386434 278618 386466 278854
rect 386702 278618 386786 278854
rect 387022 278618 387054 278854
rect 386434 261174 387054 278618
rect 386434 260938 386466 261174
rect 386702 260938 386786 261174
rect 387022 260938 387054 261174
rect 386434 260854 387054 260938
rect 386434 260618 386466 260854
rect 386702 260618 386786 260854
rect 387022 260618 387054 260854
rect 386434 243174 387054 260618
rect 386434 242938 386466 243174
rect 386702 242938 386786 243174
rect 387022 242938 387054 243174
rect 386434 242854 387054 242938
rect 386434 242618 386466 242854
rect 386702 242618 386786 242854
rect 387022 242618 387054 242854
rect 386434 225174 387054 242618
rect 386434 224938 386466 225174
rect 386702 224938 386786 225174
rect 387022 224938 387054 225174
rect 386434 224854 387054 224938
rect 386434 224618 386466 224854
rect 386702 224618 386786 224854
rect 387022 224618 387054 224854
rect 386434 207174 387054 224618
rect 386434 206938 386466 207174
rect 386702 206938 386786 207174
rect 387022 206938 387054 207174
rect 386434 206854 387054 206938
rect 386434 206618 386466 206854
rect 386702 206618 386786 206854
rect 387022 206618 387054 206854
rect 386434 189174 387054 206618
rect 386434 188938 386466 189174
rect 386702 188938 386786 189174
rect 387022 188938 387054 189174
rect 386434 188854 387054 188938
rect 386434 188618 386466 188854
rect 386702 188618 386786 188854
rect 387022 188618 387054 188854
rect 386434 171174 387054 188618
rect 386434 170938 386466 171174
rect 386702 170938 386786 171174
rect 387022 170938 387054 171174
rect 386434 170854 387054 170938
rect 386434 170618 386466 170854
rect 386702 170618 386786 170854
rect 387022 170618 387054 170854
rect 386434 153174 387054 170618
rect 386434 152938 386466 153174
rect 386702 152938 386786 153174
rect 387022 152938 387054 153174
rect 386434 152854 387054 152938
rect 386434 152618 386466 152854
rect 386702 152618 386786 152854
rect 387022 152618 387054 152854
rect 386434 135174 387054 152618
rect 386434 134938 386466 135174
rect 386702 134938 386786 135174
rect 387022 134938 387054 135174
rect 386434 134854 387054 134938
rect 386434 134618 386466 134854
rect 386702 134618 386786 134854
rect 387022 134618 387054 134854
rect 386434 117174 387054 134618
rect 386434 116938 386466 117174
rect 386702 116938 386786 117174
rect 387022 116938 387054 117174
rect 386434 116854 387054 116938
rect 386434 116618 386466 116854
rect 386702 116618 386786 116854
rect 387022 116618 387054 116854
rect 386434 99174 387054 116618
rect 386434 98938 386466 99174
rect 386702 98938 386786 99174
rect 387022 98938 387054 99174
rect 386434 98854 387054 98938
rect 386434 98618 386466 98854
rect 386702 98618 386786 98854
rect 387022 98618 387054 98854
rect 386434 81174 387054 98618
rect 386434 80938 386466 81174
rect 386702 80938 386786 81174
rect 387022 80938 387054 81174
rect 386434 80854 387054 80938
rect 386434 80618 386466 80854
rect 386702 80618 386786 80854
rect 387022 80618 387054 80854
rect 386434 63174 387054 80618
rect 386434 62938 386466 63174
rect 386702 62938 386786 63174
rect 387022 62938 387054 63174
rect 386434 62854 387054 62938
rect 386434 62618 386466 62854
rect 386702 62618 386786 62854
rect 387022 62618 387054 62854
rect 386434 45174 387054 62618
rect 386434 44938 386466 45174
rect 386702 44938 386786 45174
rect 387022 44938 387054 45174
rect 386434 44854 387054 44938
rect 386434 44618 386466 44854
rect 386702 44618 386786 44854
rect 387022 44618 387054 44854
rect 386434 27174 387054 44618
rect 386434 26938 386466 27174
rect 386702 26938 386786 27174
rect 387022 26938 387054 27174
rect 386434 26854 387054 26938
rect 386434 26618 386466 26854
rect 386702 26618 386786 26854
rect 387022 26618 387054 26854
rect 386434 9174 387054 26618
rect 386434 8938 386466 9174
rect 386702 8938 386786 9174
rect 387022 8938 387054 9174
rect 386434 8854 387054 8938
rect 386434 8618 386466 8854
rect 386702 8618 386786 8854
rect 387022 8618 387054 8854
rect 386434 -1816 387054 8618
rect 386434 -2052 386466 -1816
rect 386702 -2052 386786 -1816
rect 387022 -2052 387054 -1816
rect 386434 -2136 387054 -2052
rect 386434 -2372 386466 -2136
rect 386702 -2372 386786 -2136
rect 387022 -2372 387054 -2136
rect 386434 -4324 387054 -2372
rect 390154 463012 390774 464004
rect 390154 462776 390186 463012
rect 390422 462776 390506 463012
rect 390742 462776 390774 463012
rect 390154 462692 390774 462776
rect 390154 462456 390186 462692
rect 390422 462456 390506 462692
rect 390742 462456 390774 462692
rect 390154 444894 390774 462456
rect 390154 444658 390186 444894
rect 390422 444658 390506 444894
rect 390742 444658 390774 444894
rect 390154 444574 390774 444658
rect 390154 444338 390186 444574
rect 390422 444338 390506 444574
rect 390742 444338 390774 444574
rect 390154 426894 390774 444338
rect 390154 426658 390186 426894
rect 390422 426658 390506 426894
rect 390742 426658 390774 426894
rect 390154 426574 390774 426658
rect 390154 426338 390186 426574
rect 390422 426338 390506 426574
rect 390742 426338 390774 426574
rect 390154 408894 390774 426338
rect 390154 408658 390186 408894
rect 390422 408658 390506 408894
rect 390742 408658 390774 408894
rect 390154 408574 390774 408658
rect 390154 408338 390186 408574
rect 390422 408338 390506 408574
rect 390742 408338 390774 408574
rect 390154 390894 390774 408338
rect 390154 390658 390186 390894
rect 390422 390658 390506 390894
rect 390742 390658 390774 390894
rect 390154 390574 390774 390658
rect 390154 390338 390186 390574
rect 390422 390338 390506 390574
rect 390742 390338 390774 390574
rect 390154 372894 390774 390338
rect 390154 372658 390186 372894
rect 390422 372658 390506 372894
rect 390742 372658 390774 372894
rect 390154 372574 390774 372658
rect 390154 372338 390186 372574
rect 390422 372338 390506 372574
rect 390742 372338 390774 372574
rect 390154 354894 390774 372338
rect 390154 354658 390186 354894
rect 390422 354658 390506 354894
rect 390742 354658 390774 354894
rect 390154 354574 390774 354658
rect 390154 354338 390186 354574
rect 390422 354338 390506 354574
rect 390742 354338 390774 354574
rect 390154 336894 390774 354338
rect 390154 336658 390186 336894
rect 390422 336658 390506 336894
rect 390742 336658 390774 336894
rect 390154 336574 390774 336658
rect 390154 336338 390186 336574
rect 390422 336338 390506 336574
rect 390742 336338 390774 336574
rect 390154 318894 390774 336338
rect 390154 318658 390186 318894
rect 390422 318658 390506 318894
rect 390742 318658 390774 318894
rect 390154 318574 390774 318658
rect 390154 318338 390186 318574
rect 390422 318338 390506 318574
rect 390742 318338 390774 318574
rect 390154 300894 390774 318338
rect 390154 300658 390186 300894
rect 390422 300658 390506 300894
rect 390742 300658 390774 300894
rect 390154 300574 390774 300658
rect 390154 300338 390186 300574
rect 390422 300338 390506 300574
rect 390742 300338 390774 300574
rect 390154 282894 390774 300338
rect 390154 282658 390186 282894
rect 390422 282658 390506 282894
rect 390742 282658 390774 282894
rect 390154 282574 390774 282658
rect 390154 282338 390186 282574
rect 390422 282338 390506 282574
rect 390742 282338 390774 282574
rect 390154 264894 390774 282338
rect 390154 264658 390186 264894
rect 390422 264658 390506 264894
rect 390742 264658 390774 264894
rect 390154 264574 390774 264658
rect 390154 264338 390186 264574
rect 390422 264338 390506 264574
rect 390742 264338 390774 264574
rect 390154 246894 390774 264338
rect 390154 246658 390186 246894
rect 390422 246658 390506 246894
rect 390742 246658 390774 246894
rect 390154 246574 390774 246658
rect 390154 246338 390186 246574
rect 390422 246338 390506 246574
rect 390742 246338 390774 246574
rect 390154 228894 390774 246338
rect 390154 228658 390186 228894
rect 390422 228658 390506 228894
rect 390742 228658 390774 228894
rect 390154 228574 390774 228658
rect 390154 228338 390186 228574
rect 390422 228338 390506 228574
rect 390742 228338 390774 228574
rect 390154 210894 390774 228338
rect 390154 210658 390186 210894
rect 390422 210658 390506 210894
rect 390742 210658 390774 210894
rect 390154 210574 390774 210658
rect 390154 210338 390186 210574
rect 390422 210338 390506 210574
rect 390742 210338 390774 210574
rect 390154 192894 390774 210338
rect 390154 192658 390186 192894
rect 390422 192658 390506 192894
rect 390742 192658 390774 192894
rect 390154 192574 390774 192658
rect 390154 192338 390186 192574
rect 390422 192338 390506 192574
rect 390742 192338 390774 192574
rect 390154 174894 390774 192338
rect 390154 174658 390186 174894
rect 390422 174658 390506 174894
rect 390742 174658 390774 174894
rect 390154 174574 390774 174658
rect 390154 174338 390186 174574
rect 390422 174338 390506 174574
rect 390742 174338 390774 174574
rect 390154 156894 390774 174338
rect 390154 156658 390186 156894
rect 390422 156658 390506 156894
rect 390742 156658 390774 156894
rect 390154 156574 390774 156658
rect 390154 156338 390186 156574
rect 390422 156338 390506 156574
rect 390742 156338 390774 156574
rect 390154 138894 390774 156338
rect 390154 138658 390186 138894
rect 390422 138658 390506 138894
rect 390742 138658 390774 138894
rect 390154 138574 390774 138658
rect 390154 138338 390186 138574
rect 390422 138338 390506 138574
rect 390742 138338 390774 138574
rect 390154 120894 390774 138338
rect 390154 120658 390186 120894
rect 390422 120658 390506 120894
rect 390742 120658 390774 120894
rect 390154 120574 390774 120658
rect 390154 120338 390186 120574
rect 390422 120338 390506 120574
rect 390742 120338 390774 120574
rect 390154 102894 390774 120338
rect 390154 102658 390186 102894
rect 390422 102658 390506 102894
rect 390742 102658 390774 102894
rect 390154 102574 390774 102658
rect 390154 102338 390186 102574
rect 390422 102338 390506 102574
rect 390742 102338 390774 102574
rect 390154 84894 390774 102338
rect 390154 84658 390186 84894
rect 390422 84658 390506 84894
rect 390742 84658 390774 84894
rect 390154 84574 390774 84658
rect 390154 84338 390186 84574
rect 390422 84338 390506 84574
rect 390742 84338 390774 84574
rect 390154 66894 390774 84338
rect 390154 66658 390186 66894
rect 390422 66658 390506 66894
rect 390742 66658 390774 66894
rect 390154 66574 390774 66658
rect 390154 66338 390186 66574
rect 390422 66338 390506 66574
rect 390742 66338 390774 66574
rect 390154 48894 390774 66338
rect 390154 48658 390186 48894
rect 390422 48658 390506 48894
rect 390742 48658 390774 48894
rect 390154 48574 390774 48658
rect 390154 48338 390186 48574
rect 390422 48338 390506 48574
rect 390742 48338 390774 48574
rect 390154 30894 390774 48338
rect 390154 30658 390186 30894
rect 390422 30658 390506 30894
rect 390742 30658 390774 30894
rect 390154 30574 390774 30658
rect 390154 30338 390186 30574
rect 390422 30338 390506 30574
rect 390742 30338 390774 30574
rect 390154 12894 390774 30338
rect 390154 12658 390186 12894
rect 390422 12658 390506 12894
rect 390742 12658 390774 12894
rect 390154 12574 390774 12658
rect 390154 12338 390186 12574
rect 390422 12338 390506 12574
rect 390742 12338 390774 12574
rect 390154 -2776 390774 12338
rect 390154 -3012 390186 -2776
rect 390422 -3012 390506 -2776
rect 390742 -3012 390774 -2776
rect 390154 -3096 390774 -3012
rect 390154 -3332 390186 -3096
rect 390422 -3332 390506 -3096
rect 390742 -3332 390774 -3096
rect 390154 -4324 390774 -3332
rect 393874 463972 394494 464004
rect 393874 463736 393906 463972
rect 394142 463736 394226 463972
rect 394462 463736 394494 463972
rect 393874 463652 394494 463736
rect 393874 463416 393906 463652
rect 394142 463416 394226 463652
rect 394462 463416 394494 463652
rect 393874 448614 394494 463416
rect 393874 448378 393906 448614
rect 394142 448378 394226 448614
rect 394462 448378 394494 448614
rect 393874 448294 394494 448378
rect 393874 448058 393906 448294
rect 394142 448058 394226 448294
rect 394462 448058 394494 448294
rect 393874 430614 394494 448058
rect 393874 430378 393906 430614
rect 394142 430378 394226 430614
rect 394462 430378 394494 430614
rect 393874 430294 394494 430378
rect 393874 430058 393906 430294
rect 394142 430058 394226 430294
rect 394462 430058 394494 430294
rect 393874 412614 394494 430058
rect 393874 412378 393906 412614
rect 394142 412378 394226 412614
rect 394462 412378 394494 412614
rect 393874 412294 394494 412378
rect 393874 412058 393906 412294
rect 394142 412058 394226 412294
rect 394462 412058 394494 412294
rect 393874 394614 394494 412058
rect 393874 394378 393906 394614
rect 394142 394378 394226 394614
rect 394462 394378 394494 394614
rect 393874 394294 394494 394378
rect 393874 394058 393906 394294
rect 394142 394058 394226 394294
rect 394462 394058 394494 394294
rect 393874 376614 394494 394058
rect 393874 376378 393906 376614
rect 394142 376378 394226 376614
rect 394462 376378 394494 376614
rect 393874 376294 394494 376378
rect 393874 376058 393906 376294
rect 394142 376058 394226 376294
rect 394462 376058 394494 376294
rect 393874 358614 394494 376058
rect 393874 358378 393906 358614
rect 394142 358378 394226 358614
rect 394462 358378 394494 358614
rect 393874 358294 394494 358378
rect 393874 358058 393906 358294
rect 394142 358058 394226 358294
rect 394462 358058 394494 358294
rect 393874 340614 394494 358058
rect 393874 340378 393906 340614
rect 394142 340378 394226 340614
rect 394462 340378 394494 340614
rect 393874 340294 394494 340378
rect 393874 340058 393906 340294
rect 394142 340058 394226 340294
rect 394462 340058 394494 340294
rect 393874 322614 394494 340058
rect 393874 322378 393906 322614
rect 394142 322378 394226 322614
rect 394462 322378 394494 322614
rect 393874 322294 394494 322378
rect 393874 322058 393906 322294
rect 394142 322058 394226 322294
rect 394462 322058 394494 322294
rect 393874 304614 394494 322058
rect 393874 304378 393906 304614
rect 394142 304378 394226 304614
rect 394462 304378 394494 304614
rect 393874 304294 394494 304378
rect 393874 304058 393906 304294
rect 394142 304058 394226 304294
rect 394462 304058 394494 304294
rect 393874 286614 394494 304058
rect 393874 286378 393906 286614
rect 394142 286378 394226 286614
rect 394462 286378 394494 286614
rect 393874 286294 394494 286378
rect 393874 286058 393906 286294
rect 394142 286058 394226 286294
rect 394462 286058 394494 286294
rect 393874 268614 394494 286058
rect 393874 268378 393906 268614
rect 394142 268378 394226 268614
rect 394462 268378 394494 268614
rect 393874 268294 394494 268378
rect 393874 268058 393906 268294
rect 394142 268058 394226 268294
rect 394462 268058 394494 268294
rect 393874 250614 394494 268058
rect 393874 250378 393906 250614
rect 394142 250378 394226 250614
rect 394462 250378 394494 250614
rect 393874 250294 394494 250378
rect 393874 250058 393906 250294
rect 394142 250058 394226 250294
rect 394462 250058 394494 250294
rect 393874 232614 394494 250058
rect 393874 232378 393906 232614
rect 394142 232378 394226 232614
rect 394462 232378 394494 232614
rect 393874 232294 394494 232378
rect 393874 232058 393906 232294
rect 394142 232058 394226 232294
rect 394462 232058 394494 232294
rect 393874 214614 394494 232058
rect 393874 214378 393906 214614
rect 394142 214378 394226 214614
rect 394462 214378 394494 214614
rect 393874 214294 394494 214378
rect 393874 214058 393906 214294
rect 394142 214058 394226 214294
rect 394462 214058 394494 214294
rect 393874 196614 394494 214058
rect 393874 196378 393906 196614
rect 394142 196378 394226 196614
rect 394462 196378 394494 196614
rect 393874 196294 394494 196378
rect 393874 196058 393906 196294
rect 394142 196058 394226 196294
rect 394462 196058 394494 196294
rect 393874 178614 394494 196058
rect 393874 178378 393906 178614
rect 394142 178378 394226 178614
rect 394462 178378 394494 178614
rect 393874 178294 394494 178378
rect 393874 178058 393906 178294
rect 394142 178058 394226 178294
rect 394462 178058 394494 178294
rect 393874 160614 394494 178058
rect 393874 160378 393906 160614
rect 394142 160378 394226 160614
rect 394462 160378 394494 160614
rect 393874 160294 394494 160378
rect 393874 160058 393906 160294
rect 394142 160058 394226 160294
rect 394462 160058 394494 160294
rect 393874 142614 394494 160058
rect 393874 142378 393906 142614
rect 394142 142378 394226 142614
rect 394462 142378 394494 142614
rect 393874 142294 394494 142378
rect 393874 142058 393906 142294
rect 394142 142058 394226 142294
rect 394462 142058 394494 142294
rect 393874 124614 394494 142058
rect 393874 124378 393906 124614
rect 394142 124378 394226 124614
rect 394462 124378 394494 124614
rect 393874 124294 394494 124378
rect 393874 124058 393906 124294
rect 394142 124058 394226 124294
rect 394462 124058 394494 124294
rect 393874 106614 394494 124058
rect 393874 106378 393906 106614
rect 394142 106378 394226 106614
rect 394462 106378 394494 106614
rect 393874 106294 394494 106378
rect 393874 106058 393906 106294
rect 394142 106058 394226 106294
rect 394462 106058 394494 106294
rect 393874 88614 394494 106058
rect 393874 88378 393906 88614
rect 394142 88378 394226 88614
rect 394462 88378 394494 88614
rect 393874 88294 394494 88378
rect 393874 88058 393906 88294
rect 394142 88058 394226 88294
rect 394462 88058 394494 88294
rect 393874 70614 394494 88058
rect 393874 70378 393906 70614
rect 394142 70378 394226 70614
rect 394462 70378 394494 70614
rect 393874 70294 394494 70378
rect 393874 70058 393906 70294
rect 394142 70058 394226 70294
rect 394462 70058 394494 70294
rect 393874 52614 394494 70058
rect 393874 52378 393906 52614
rect 394142 52378 394226 52614
rect 394462 52378 394494 52614
rect 393874 52294 394494 52378
rect 393874 52058 393906 52294
rect 394142 52058 394226 52294
rect 394462 52058 394494 52294
rect 393874 34614 394494 52058
rect 393874 34378 393906 34614
rect 394142 34378 394226 34614
rect 394462 34378 394494 34614
rect 393874 34294 394494 34378
rect 393874 34058 393906 34294
rect 394142 34058 394226 34294
rect 394462 34058 394494 34294
rect 393874 16614 394494 34058
rect 393874 16378 393906 16614
rect 394142 16378 394226 16614
rect 394462 16378 394494 16614
rect 393874 16294 394494 16378
rect 393874 16058 393906 16294
rect 394142 16058 394226 16294
rect 394462 16058 394494 16294
rect 393874 -3736 394494 16058
rect 393874 -3972 393906 -3736
rect 394142 -3972 394226 -3736
rect 394462 -3972 394494 -3736
rect 393874 -4056 394494 -3972
rect 393874 -4292 393906 -4056
rect 394142 -4292 394226 -4056
rect 394462 -4292 394494 -4056
rect 393874 -4324 394494 -4292
rect 400714 461092 401334 464004
rect 400714 460856 400746 461092
rect 400982 460856 401066 461092
rect 401302 460856 401334 461092
rect 400714 460772 401334 460856
rect 400714 460536 400746 460772
rect 400982 460536 401066 460772
rect 401302 460536 401334 460772
rect 400714 455454 401334 460536
rect 400714 455218 400746 455454
rect 400982 455218 401066 455454
rect 401302 455218 401334 455454
rect 400714 455134 401334 455218
rect 400714 454898 400746 455134
rect 400982 454898 401066 455134
rect 401302 454898 401334 455134
rect 400714 437454 401334 454898
rect 400714 437218 400746 437454
rect 400982 437218 401066 437454
rect 401302 437218 401334 437454
rect 400714 437134 401334 437218
rect 400714 436898 400746 437134
rect 400982 436898 401066 437134
rect 401302 436898 401334 437134
rect 400714 419454 401334 436898
rect 400714 419218 400746 419454
rect 400982 419218 401066 419454
rect 401302 419218 401334 419454
rect 400714 419134 401334 419218
rect 400714 418898 400746 419134
rect 400982 418898 401066 419134
rect 401302 418898 401334 419134
rect 400714 401454 401334 418898
rect 400714 401218 400746 401454
rect 400982 401218 401066 401454
rect 401302 401218 401334 401454
rect 400714 401134 401334 401218
rect 400714 400898 400746 401134
rect 400982 400898 401066 401134
rect 401302 400898 401334 401134
rect 400714 383454 401334 400898
rect 400714 383218 400746 383454
rect 400982 383218 401066 383454
rect 401302 383218 401334 383454
rect 400714 383134 401334 383218
rect 400714 382898 400746 383134
rect 400982 382898 401066 383134
rect 401302 382898 401334 383134
rect 400714 365454 401334 382898
rect 400714 365218 400746 365454
rect 400982 365218 401066 365454
rect 401302 365218 401334 365454
rect 400714 365134 401334 365218
rect 400714 364898 400746 365134
rect 400982 364898 401066 365134
rect 401302 364898 401334 365134
rect 400714 347454 401334 364898
rect 400714 347218 400746 347454
rect 400982 347218 401066 347454
rect 401302 347218 401334 347454
rect 400714 347134 401334 347218
rect 400714 346898 400746 347134
rect 400982 346898 401066 347134
rect 401302 346898 401334 347134
rect 400714 329454 401334 346898
rect 400714 329218 400746 329454
rect 400982 329218 401066 329454
rect 401302 329218 401334 329454
rect 400714 329134 401334 329218
rect 400714 328898 400746 329134
rect 400982 328898 401066 329134
rect 401302 328898 401334 329134
rect 400714 311454 401334 328898
rect 400714 311218 400746 311454
rect 400982 311218 401066 311454
rect 401302 311218 401334 311454
rect 400714 311134 401334 311218
rect 400714 310898 400746 311134
rect 400982 310898 401066 311134
rect 401302 310898 401334 311134
rect 400714 293454 401334 310898
rect 400714 293218 400746 293454
rect 400982 293218 401066 293454
rect 401302 293218 401334 293454
rect 400714 293134 401334 293218
rect 400714 292898 400746 293134
rect 400982 292898 401066 293134
rect 401302 292898 401334 293134
rect 400714 275454 401334 292898
rect 400714 275218 400746 275454
rect 400982 275218 401066 275454
rect 401302 275218 401334 275454
rect 400714 275134 401334 275218
rect 400714 274898 400746 275134
rect 400982 274898 401066 275134
rect 401302 274898 401334 275134
rect 400714 257454 401334 274898
rect 400714 257218 400746 257454
rect 400982 257218 401066 257454
rect 401302 257218 401334 257454
rect 400714 257134 401334 257218
rect 400714 256898 400746 257134
rect 400982 256898 401066 257134
rect 401302 256898 401334 257134
rect 400714 239454 401334 256898
rect 400714 239218 400746 239454
rect 400982 239218 401066 239454
rect 401302 239218 401334 239454
rect 400714 239134 401334 239218
rect 400714 238898 400746 239134
rect 400982 238898 401066 239134
rect 401302 238898 401334 239134
rect 400714 221454 401334 238898
rect 400714 221218 400746 221454
rect 400982 221218 401066 221454
rect 401302 221218 401334 221454
rect 400714 221134 401334 221218
rect 400714 220898 400746 221134
rect 400982 220898 401066 221134
rect 401302 220898 401334 221134
rect 400714 203454 401334 220898
rect 400714 203218 400746 203454
rect 400982 203218 401066 203454
rect 401302 203218 401334 203454
rect 400714 203134 401334 203218
rect 400714 202898 400746 203134
rect 400982 202898 401066 203134
rect 401302 202898 401334 203134
rect 400714 185454 401334 202898
rect 400714 185218 400746 185454
rect 400982 185218 401066 185454
rect 401302 185218 401334 185454
rect 400714 185134 401334 185218
rect 400714 184898 400746 185134
rect 400982 184898 401066 185134
rect 401302 184898 401334 185134
rect 400714 167454 401334 184898
rect 400714 167218 400746 167454
rect 400982 167218 401066 167454
rect 401302 167218 401334 167454
rect 400714 167134 401334 167218
rect 400714 166898 400746 167134
rect 400982 166898 401066 167134
rect 401302 166898 401334 167134
rect 400714 149454 401334 166898
rect 400714 149218 400746 149454
rect 400982 149218 401066 149454
rect 401302 149218 401334 149454
rect 400714 149134 401334 149218
rect 400714 148898 400746 149134
rect 400982 148898 401066 149134
rect 401302 148898 401334 149134
rect 400714 131454 401334 148898
rect 400714 131218 400746 131454
rect 400982 131218 401066 131454
rect 401302 131218 401334 131454
rect 400714 131134 401334 131218
rect 400714 130898 400746 131134
rect 400982 130898 401066 131134
rect 401302 130898 401334 131134
rect 400714 113454 401334 130898
rect 400714 113218 400746 113454
rect 400982 113218 401066 113454
rect 401302 113218 401334 113454
rect 400714 113134 401334 113218
rect 400714 112898 400746 113134
rect 400982 112898 401066 113134
rect 401302 112898 401334 113134
rect 400714 95454 401334 112898
rect 400714 95218 400746 95454
rect 400982 95218 401066 95454
rect 401302 95218 401334 95454
rect 400714 95134 401334 95218
rect 400714 94898 400746 95134
rect 400982 94898 401066 95134
rect 401302 94898 401334 95134
rect 400714 77454 401334 94898
rect 400714 77218 400746 77454
rect 400982 77218 401066 77454
rect 401302 77218 401334 77454
rect 400714 77134 401334 77218
rect 400714 76898 400746 77134
rect 400982 76898 401066 77134
rect 401302 76898 401334 77134
rect 400714 59454 401334 76898
rect 400714 59218 400746 59454
rect 400982 59218 401066 59454
rect 401302 59218 401334 59454
rect 400714 59134 401334 59218
rect 400714 58898 400746 59134
rect 400982 58898 401066 59134
rect 401302 58898 401334 59134
rect 400714 41454 401334 58898
rect 400714 41218 400746 41454
rect 400982 41218 401066 41454
rect 401302 41218 401334 41454
rect 400714 41134 401334 41218
rect 400714 40898 400746 41134
rect 400982 40898 401066 41134
rect 401302 40898 401334 41134
rect 400714 23454 401334 40898
rect 400714 23218 400746 23454
rect 400982 23218 401066 23454
rect 401302 23218 401334 23454
rect 400714 23134 401334 23218
rect 400714 22898 400746 23134
rect 400982 22898 401066 23134
rect 401302 22898 401334 23134
rect 400714 5454 401334 22898
rect 400714 5218 400746 5454
rect 400982 5218 401066 5454
rect 401302 5218 401334 5454
rect 400714 5134 401334 5218
rect 400714 4898 400746 5134
rect 400982 4898 401066 5134
rect 401302 4898 401334 5134
rect 400714 -856 401334 4898
rect 400714 -1092 400746 -856
rect 400982 -1092 401066 -856
rect 401302 -1092 401334 -856
rect 400714 -1176 401334 -1092
rect 400714 -1412 400746 -1176
rect 400982 -1412 401066 -1176
rect 401302 -1412 401334 -1176
rect 400714 -4324 401334 -1412
rect 404434 462052 405054 464004
rect 404434 461816 404466 462052
rect 404702 461816 404786 462052
rect 405022 461816 405054 462052
rect 404434 461732 405054 461816
rect 404434 461496 404466 461732
rect 404702 461496 404786 461732
rect 405022 461496 405054 461732
rect 404434 441174 405054 461496
rect 404434 440938 404466 441174
rect 404702 440938 404786 441174
rect 405022 440938 405054 441174
rect 404434 440854 405054 440938
rect 404434 440618 404466 440854
rect 404702 440618 404786 440854
rect 405022 440618 405054 440854
rect 404434 423174 405054 440618
rect 404434 422938 404466 423174
rect 404702 422938 404786 423174
rect 405022 422938 405054 423174
rect 404434 422854 405054 422938
rect 404434 422618 404466 422854
rect 404702 422618 404786 422854
rect 405022 422618 405054 422854
rect 404434 405174 405054 422618
rect 404434 404938 404466 405174
rect 404702 404938 404786 405174
rect 405022 404938 405054 405174
rect 404434 404854 405054 404938
rect 404434 404618 404466 404854
rect 404702 404618 404786 404854
rect 405022 404618 405054 404854
rect 404434 387174 405054 404618
rect 404434 386938 404466 387174
rect 404702 386938 404786 387174
rect 405022 386938 405054 387174
rect 404434 386854 405054 386938
rect 404434 386618 404466 386854
rect 404702 386618 404786 386854
rect 405022 386618 405054 386854
rect 404434 369174 405054 386618
rect 404434 368938 404466 369174
rect 404702 368938 404786 369174
rect 405022 368938 405054 369174
rect 404434 368854 405054 368938
rect 404434 368618 404466 368854
rect 404702 368618 404786 368854
rect 405022 368618 405054 368854
rect 404434 351174 405054 368618
rect 404434 350938 404466 351174
rect 404702 350938 404786 351174
rect 405022 350938 405054 351174
rect 404434 350854 405054 350938
rect 404434 350618 404466 350854
rect 404702 350618 404786 350854
rect 405022 350618 405054 350854
rect 404434 333174 405054 350618
rect 404434 332938 404466 333174
rect 404702 332938 404786 333174
rect 405022 332938 405054 333174
rect 404434 332854 405054 332938
rect 404434 332618 404466 332854
rect 404702 332618 404786 332854
rect 405022 332618 405054 332854
rect 404434 315174 405054 332618
rect 404434 314938 404466 315174
rect 404702 314938 404786 315174
rect 405022 314938 405054 315174
rect 404434 314854 405054 314938
rect 404434 314618 404466 314854
rect 404702 314618 404786 314854
rect 405022 314618 405054 314854
rect 404434 297174 405054 314618
rect 404434 296938 404466 297174
rect 404702 296938 404786 297174
rect 405022 296938 405054 297174
rect 404434 296854 405054 296938
rect 404434 296618 404466 296854
rect 404702 296618 404786 296854
rect 405022 296618 405054 296854
rect 404434 279174 405054 296618
rect 404434 278938 404466 279174
rect 404702 278938 404786 279174
rect 405022 278938 405054 279174
rect 404434 278854 405054 278938
rect 404434 278618 404466 278854
rect 404702 278618 404786 278854
rect 405022 278618 405054 278854
rect 404434 261174 405054 278618
rect 404434 260938 404466 261174
rect 404702 260938 404786 261174
rect 405022 260938 405054 261174
rect 404434 260854 405054 260938
rect 404434 260618 404466 260854
rect 404702 260618 404786 260854
rect 405022 260618 405054 260854
rect 404434 243174 405054 260618
rect 404434 242938 404466 243174
rect 404702 242938 404786 243174
rect 405022 242938 405054 243174
rect 404434 242854 405054 242938
rect 404434 242618 404466 242854
rect 404702 242618 404786 242854
rect 405022 242618 405054 242854
rect 404434 225174 405054 242618
rect 404434 224938 404466 225174
rect 404702 224938 404786 225174
rect 405022 224938 405054 225174
rect 404434 224854 405054 224938
rect 404434 224618 404466 224854
rect 404702 224618 404786 224854
rect 405022 224618 405054 224854
rect 404434 207174 405054 224618
rect 404434 206938 404466 207174
rect 404702 206938 404786 207174
rect 405022 206938 405054 207174
rect 404434 206854 405054 206938
rect 404434 206618 404466 206854
rect 404702 206618 404786 206854
rect 405022 206618 405054 206854
rect 404434 189174 405054 206618
rect 404434 188938 404466 189174
rect 404702 188938 404786 189174
rect 405022 188938 405054 189174
rect 404434 188854 405054 188938
rect 404434 188618 404466 188854
rect 404702 188618 404786 188854
rect 405022 188618 405054 188854
rect 404434 171174 405054 188618
rect 404434 170938 404466 171174
rect 404702 170938 404786 171174
rect 405022 170938 405054 171174
rect 404434 170854 405054 170938
rect 404434 170618 404466 170854
rect 404702 170618 404786 170854
rect 405022 170618 405054 170854
rect 404434 153174 405054 170618
rect 404434 152938 404466 153174
rect 404702 152938 404786 153174
rect 405022 152938 405054 153174
rect 404434 152854 405054 152938
rect 404434 152618 404466 152854
rect 404702 152618 404786 152854
rect 405022 152618 405054 152854
rect 404434 135174 405054 152618
rect 404434 134938 404466 135174
rect 404702 134938 404786 135174
rect 405022 134938 405054 135174
rect 404434 134854 405054 134938
rect 404434 134618 404466 134854
rect 404702 134618 404786 134854
rect 405022 134618 405054 134854
rect 404434 117174 405054 134618
rect 404434 116938 404466 117174
rect 404702 116938 404786 117174
rect 405022 116938 405054 117174
rect 404434 116854 405054 116938
rect 404434 116618 404466 116854
rect 404702 116618 404786 116854
rect 405022 116618 405054 116854
rect 404434 99174 405054 116618
rect 404434 98938 404466 99174
rect 404702 98938 404786 99174
rect 405022 98938 405054 99174
rect 404434 98854 405054 98938
rect 404434 98618 404466 98854
rect 404702 98618 404786 98854
rect 405022 98618 405054 98854
rect 404434 81174 405054 98618
rect 404434 80938 404466 81174
rect 404702 80938 404786 81174
rect 405022 80938 405054 81174
rect 404434 80854 405054 80938
rect 404434 80618 404466 80854
rect 404702 80618 404786 80854
rect 405022 80618 405054 80854
rect 404434 63174 405054 80618
rect 404434 62938 404466 63174
rect 404702 62938 404786 63174
rect 405022 62938 405054 63174
rect 404434 62854 405054 62938
rect 404434 62618 404466 62854
rect 404702 62618 404786 62854
rect 405022 62618 405054 62854
rect 404434 45174 405054 62618
rect 404434 44938 404466 45174
rect 404702 44938 404786 45174
rect 405022 44938 405054 45174
rect 404434 44854 405054 44938
rect 404434 44618 404466 44854
rect 404702 44618 404786 44854
rect 405022 44618 405054 44854
rect 404434 27174 405054 44618
rect 404434 26938 404466 27174
rect 404702 26938 404786 27174
rect 405022 26938 405054 27174
rect 404434 26854 405054 26938
rect 404434 26618 404466 26854
rect 404702 26618 404786 26854
rect 405022 26618 405054 26854
rect 404434 9174 405054 26618
rect 404434 8938 404466 9174
rect 404702 8938 404786 9174
rect 405022 8938 405054 9174
rect 404434 8854 405054 8938
rect 404434 8618 404466 8854
rect 404702 8618 404786 8854
rect 405022 8618 405054 8854
rect 404434 -1816 405054 8618
rect 404434 -2052 404466 -1816
rect 404702 -2052 404786 -1816
rect 405022 -2052 405054 -1816
rect 404434 -2136 405054 -2052
rect 404434 -2372 404466 -2136
rect 404702 -2372 404786 -2136
rect 405022 -2372 405054 -2136
rect 404434 -4324 405054 -2372
rect 408154 463012 408774 464004
rect 408154 462776 408186 463012
rect 408422 462776 408506 463012
rect 408742 462776 408774 463012
rect 408154 462692 408774 462776
rect 408154 462456 408186 462692
rect 408422 462456 408506 462692
rect 408742 462456 408774 462692
rect 408154 444894 408774 462456
rect 408154 444658 408186 444894
rect 408422 444658 408506 444894
rect 408742 444658 408774 444894
rect 408154 444574 408774 444658
rect 408154 444338 408186 444574
rect 408422 444338 408506 444574
rect 408742 444338 408774 444574
rect 408154 426894 408774 444338
rect 408154 426658 408186 426894
rect 408422 426658 408506 426894
rect 408742 426658 408774 426894
rect 408154 426574 408774 426658
rect 408154 426338 408186 426574
rect 408422 426338 408506 426574
rect 408742 426338 408774 426574
rect 408154 408894 408774 426338
rect 408154 408658 408186 408894
rect 408422 408658 408506 408894
rect 408742 408658 408774 408894
rect 408154 408574 408774 408658
rect 408154 408338 408186 408574
rect 408422 408338 408506 408574
rect 408742 408338 408774 408574
rect 408154 390894 408774 408338
rect 408154 390658 408186 390894
rect 408422 390658 408506 390894
rect 408742 390658 408774 390894
rect 408154 390574 408774 390658
rect 408154 390338 408186 390574
rect 408422 390338 408506 390574
rect 408742 390338 408774 390574
rect 408154 372894 408774 390338
rect 408154 372658 408186 372894
rect 408422 372658 408506 372894
rect 408742 372658 408774 372894
rect 408154 372574 408774 372658
rect 408154 372338 408186 372574
rect 408422 372338 408506 372574
rect 408742 372338 408774 372574
rect 408154 354894 408774 372338
rect 408154 354658 408186 354894
rect 408422 354658 408506 354894
rect 408742 354658 408774 354894
rect 408154 354574 408774 354658
rect 408154 354338 408186 354574
rect 408422 354338 408506 354574
rect 408742 354338 408774 354574
rect 408154 336894 408774 354338
rect 408154 336658 408186 336894
rect 408422 336658 408506 336894
rect 408742 336658 408774 336894
rect 408154 336574 408774 336658
rect 408154 336338 408186 336574
rect 408422 336338 408506 336574
rect 408742 336338 408774 336574
rect 408154 318894 408774 336338
rect 408154 318658 408186 318894
rect 408422 318658 408506 318894
rect 408742 318658 408774 318894
rect 408154 318574 408774 318658
rect 408154 318338 408186 318574
rect 408422 318338 408506 318574
rect 408742 318338 408774 318574
rect 408154 300894 408774 318338
rect 408154 300658 408186 300894
rect 408422 300658 408506 300894
rect 408742 300658 408774 300894
rect 408154 300574 408774 300658
rect 408154 300338 408186 300574
rect 408422 300338 408506 300574
rect 408742 300338 408774 300574
rect 408154 282894 408774 300338
rect 408154 282658 408186 282894
rect 408422 282658 408506 282894
rect 408742 282658 408774 282894
rect 408154 282574 408774 282658
rect 408154 282338 408186 282574
rect 408422 282338 408506 282574
rect 408742 282338 408774 282574
rect 408154 264894 408774 282338
rect 408154 264658 408186 264894
rect 408422 264658 408506 264894
rect 408742 264658 408774 264894
rect 408154 264574 408774 264658
rect 408154 264338 408186 264574
rect 408422 264338 408506 264574
rect 408742 264338 408774 264574
rect 408154 246894 408774 264338
rect 408154 246658 408186 246894
rect 408422 246658 408506 246894
rect 408742 246658 408774 246894
rect 408154 246574 408774 246658
rect 408154 246338 408186 246574
rect 408422 246338 408506 246574
rect 408742 246338 408774 246574
rect 408154 228894 408774 246338
rect 408154 228658 408186 228894
rect 408422 228658 408506 228894
rect 408742 228658 408774 228894
rect 408154 228574 408774 228658
rect 408154 228338 408186 228574
rect 408422 228338 408506 228574
rect 408742 228338 408774 228574
rect 408154 210894 408774 228338
rect 408154 210658 408186 210894
rect 408422 210658 408506 210894
rect 408742 210658 408774 210894
rect 408154 210574 408774 210658
rect 408154 210338 408186 210574
rect 408422 210338 408506 210574
rect 408742 210338 408774 210574
rect 408154 192894 408774 210338
rect 408154 192658 408186 192894
rect 408422 192658 408506 192894
rect 408742 192658 408774 192894
rect 408154 192574 408774 192658
rect 408154 192338 408186 192574
rect 408422 192338 408506 192574
rect 408742 192338 408774 192574
rect 408154 174894 408774 192338
rect 408154 174658 408186 174894
rect 408422 174658 408506 174894
rect 408742 174658 408774 174894
rect 408154 174574 408774 174658
rect 408154 174338 408186 174574
rect 408422 174338 408506 174574
rect 408742 174338 408774 174574
rect 408154 156894 408774 174338
rect 408154 156658 408186 156894
rect 408422 156658 408506 156894
rect 408742 156658 408774 156894
rect 408154 156574 408774 156658
rect 408154 156338 408186 156574
rect 408422 156338 408506 156574
rect 408742 156338 408774 156574
rect 408154 138894 408774 156338
rect 408154 138658 408186 138894
rect 408422 138658 408506 138894
rect 408742 138658 408774 138894
rect 408154 138574 408774 138658
rect 408154 138338 408186 138574
rect 408422 138338 408506 138574
rect 408742 138338 408774 138574
rect 408154 120894 408774 138338
rect 408154 120658 408186 120894
rect 408422 120658 408506 120894
rect 408742 120658 408774 120894
rect 408154 120574 408774 120658
rect 408154 120338 408186 120574
rect 408422 120338 408506 120574
rect 408742 120338 408774 120574
rect 408154 102894 408774 120338
rect 408154 102658 408186 102894
rect 408422 102658 408506 102894
rect 408742 102658 408774 102894
rect 408154 102574 408774 102658
rect 408154 102338 408186 102574
rect 408422 102338 408506 102574
rect 408742 102338 408774 102574
rect 408154 84894 408774 102338
rect 408154 84658 408186 84894
rect 408422 84658 408506 84894
rect 408742 84658 408774 84894
rect 408154 84574 408774 84658
rect 408154 84338 408186 84574
rect 408422 84338 408506 84574
rect 408742 84338 408774 84574
rect 408154 66894 408774 84338
rect 408154 66658 408186 66894
rect 408422 66658 408506 66894
rect 408742 66658 408774 66894
rect 408154 66574 408774 66658
rect 408154 66338 408186 66574
rect 408422 66338 408506 66574
rect 408742 66338 408774 66574
rect 408154 48894 408774 66338
rect 408154 48658 408186 48894
rect 408422 48658 408506 48894
rect 408742 48658 408774 48894
rect 408154 48574 408774 48658
rect 408154 48338 408186 48574
rect 408422 48338 408506 48574
rect 408742 48338 408774 48574
rect 408154 30894 408774 48338
rect 408154 30658 408186 30894
rect 408422 30658 408506 30894
rect 408742 30658 408774 30894
rect 408154 30574 408774 30658
rect 408154 30338 408186 30574
rect 408422 30338 408506 30574
rect 408742 30338 408774 30574
rect 408154 12894 408774 30338
rect 408154 12658 408186 12894
rect 408422 12658 408506 12894
rect 408742 12658 408774 12894
rect 408154 12574 408774 12658
rect 408154 12338 408186 12574
rect 408422 12338 408506 12574
rect 408742 12338 408774 12574
rect 408154 -2776 408774 12338
rect 408154 -3012 408186 -2776
rect 408422 -3012 408506 -2776
rect 408742 -3012 408774 -2776
rect 408154 -3096 408774 -3012
rect 408154 -3332 408186 -3096
rect 408422 -3332 408506 -3096
rect 408742 -3332 408774 -3096
rect 408154 -4324 408774 -3332
rect 411874 463972 412494 464004
rect 411874 463736 411906 463972
rect 412142 463736 412226 463972
rect 412462 463736 412494 463972
rect 411874 463652 412494 463736
rect 411874 463416 411906 463652
rect 412142 463416 412226 463652
rect 412462 463416 412494 463652
rect 411874 448614 412494 463416
rect 411874 448378 411906 448614
rect 412142 448378 412226 448614
rect 412462 448378 412494 448614
rect 411874 448294 412494 448378
rect 411874 448058 411906 448294
rect 412142 448058 412226 448294
rect 412462 448058 412494 448294
rect 411874 430614 412494 448058
rect 411874 430378 411906 430614
rect 412142 430378 412226 430614
rect 412462 430378 412494 430614
rect 411874 430294 412494 430378
rect 411874 430058 411906 430294
rect 412142 430058 412226 430294
rect 412462 430058 412494 430294
rect 411874 412614 412494 430058
rect 411874 412378 411906 412614
rect 412142 412378 412226 412614
rect 412462 412378 412494 412614
rect 411874 412294 412494 412378
rect 411874 412058 411906 412294
rect 412142 412058 412226 412294
rect 412462 412058 412494 412294
rect 411874 394614 412494 412058
rect 411874 394378 411906 394614
rect 412142 394378 412226 394614
rect 412462 394378 412494 394614
rect 411874 394294 412494 394378
rect 411874 394058 411906 394294
rect 412142 394058 412226 394294
rect 412462 394058 412494 394294
rect 411874 376614 412494 394058
rect 411874 376378 411906 376614
rect 412142 376378 412226 376614
rect 412462 376378 412494 376614
rect 411874 376294 412494 376378
rect 411874 376058 411906 376294
rect 412142 376058 412226 376294
rect 412462 376058 412494 376294
rect 411874 358614 412494 376058
rect 411874 358378 411906 358614
rect 412142 358378 412226 358614
rect 412462 358378 412494 358614
rect 411874 358294 412494 358378
rect 411874 358058 411906 358294
rect 412142 358058 412226 358294
rect 412462 358058 412494 358294
rect 411874 340614 412494 358058
rect 411874 340378 411906 340614
rect 412142 340378 412226 340614
rect 412462 340378 412494 340614
rect 411874 340294 412494 340378
rect 411874 340058 411906 340294
rect 412142 340058 412226 340294
rect 412462 340058 412494 340294
rect 411874 322614 412494 340058
rect 411874 322378 411906 322614
rect 412142 322378 412226 322614
rect 412462 322378 412494 322614
rect 411874 322294 412494 322378
rect 411874 322058 411906 322294
rect 412142 322058 412226 322294
rect 412462 322058 412494 322294
rect 411874 304614 412494 322058
rect 411874 304378 411906 304614
rect 412142 304378 412226 304614
rect 412462 304378 412494 304614
rect 411874 304294 412494 304378
rect 411874 304058 411906 304294
rect 412142 304058 412226 304294
rect 412462 304058 412494 304294
rect 411874 286614 412494 304058
rect 411874 286378 411906 286614
rect 412142 286378 412226 286614
rect 412462 286378 412494 286614
rect 411874 286294 412494 286378
rect 411874 286058 411906 286294
rect 412142 286058 412226 286294
rect 412462 286058 412494 286294
rect 411874 268614 412494 286058
rect 411874 268378 411906 268614
rect 412142 268378 412226 268614
rect 412462 268378 412494 268614
rect 411874 268294 412494 268378
rect 411874 268058 411906 268294
rect 412142 268058 412226 268294
rect 412462 268058 412494 268294
rect 411874 250614 412494 268058
rect 411874 250378 411906 250614
rect 412142 250378 412226 250614
rect 412462 250378 412494 250614
rect 411874 250294 412494 250378
rect 411874 250058 411906 250294
rect 412142 250058 412226 250294
rect 412462 250058 412494 250294
rect 411874 232614 412494 250058
rect 411874 232378 411906 232614
rect 412142 232378 412226 232614
rect 412462 232378 412494 232614
rect 411874 232294 412494 232378
rect 411874 232058 411906 232294
rect 412142 232058 412226 232294
rect 412462 232058 412494 232294
rect 411874 214614 412494 232058
rect 411874 214378 411906 214614
rect 412142 214378 412226 214614
rect 412462 214378 412494 214614
rect 411874 214294 412494 214378
rect 411874 214058 411906 214294
rect 412142 214058 412226 214294
rect 412462 214058 412494 214294
rect 411874 196614 412494 214058
rect 411874 196378 411906 196614
rect 412142 196378 412226 196614
rect 412462 196378 412494 196614
rect 411874 196294 412494 196378
rect 411874 196058 411906 196294
rect 412142 196058 412226 196294
rect 412462 196058 412494 196294
rect 411874 178614 412494 196058
rect 411874 178378 411906 178614
rect 412142 178378 412226 178614
rect 412462 178378 412494 178614
rect 411874 178294 412494 178378
rect 411874 178058 411906 178294
rect 412142 178058 412226 178294
rect 412462 178058 412494 178294
rect 411874 160614 412494 178058
rect 411874 160378 411906 160614
rect 412142 160378 412226 160614
rect 412462 160378 412494 160614
rect 411874 160294 412494 160378
rect 411874 160058 411906 160294
rect 412142 160058 412226 160294
rect 412462 160058 412494 160294
rect 411874 142614 412494 160058
rect 411874 142378 411906 142614
rect 412142 142378 412226 142614
rect 412462 142378 412494 142614
rect 411874 142294 412494 142378
rect 411874 142058 411906 142294
rect 412142 142058 412226 142294
rect 412462 142058 412494 142294
rect 411874 124614 412494 142058
rect 411874 124378 411906 124614
rect 412142 124378 412226 124614
rect 412462 124378 412494 124614
rect 411874 124294 412494 124378
rect 411874 124058 411906 124294
rect 412142 124058 412226 124294
rect 412462 124058 412494 124294
rect 411874 106614 412494 124058
rect 411874 106378 411906 106614
rect 412142 106378 412226 106614
rect 412462 106378 412494 106614
rect 411874 106294 412494 106378
rect 411874 106058 411906 106294
rect 412142 106058 412226 106294
rect 412462 106058 412494 106294
rect 411874 88614 412494 106058
rect 411874 88378 411906 88614
rect 412142 88378 412226 88614
rect 412462 88378 412494 88614
rect 411874 88294 412494 88378
rect 411874 88058 411906 88294
rect 412142 88058 412226 88294
rect 412462 88058 412494 88294
rect 411874 70614 412494 88058
rect 411874 70378 411906 70614
rect 412142 70378 412226 70614
rect 412462 70378 412494 70614
rect 411874 70294 412494 70378
rect 411874 70058 411906 70294
rect 412142 70058 412226 70294
rect 412462 70058 412494 70294
rect 411874 52614 412494 70058
rect 411874 52378 411906 52614
rect 412142 52378 412226 52614
rect 412462 52378 412494 52614
rect 411874 52294 412494 52378
rect 411874 52058 411906 52294
rect 412142 52058 412226 52294
rect 412462 52058 412494 52294
rect 411874 34614 412494 52058
rect 411874 34378 411906 34614
rect 412142 34378 412226 34614
rect 412462 34378 412494 34614
rect 411874 34294 412494 34378
rect 411874 34058 411906 34294
rect 412142 34058 412226 34294
rect 412462 34058 412494 34294
rect 411874 16614 412494 34058
rect 411874 16378 411906 16614
rect 412142 16378 412226 16614
rect 412462 16378 412494 16614
rect 411874 16294 412494 16378
rect 411874 16058 411906 16294
rect 412142 16058 412226 16294
rect 412462 16058 412494 16294
rect 411874 -3736 412494 16058
rect 411874 -3972 411906 -3736
rect 412142 -3972 412226 -3736
rect 412462 -3972 412494 -3736
rect 411874 -4056 412494 -3972
rect 411874 -4292 411906 -4056
rect 412142 -4292 412226 -4056
rect 412462 -4292 412494 -4056
rect 411874 -4324 412494 -4292
rect 418714 461092 419334 464004
rect 418714 460856 418746 461092
rect 418982 460856 419066 461092
rect 419302 460856 419334 461092
rect 418714 460772 419334 460856
rect 418714 460536 418746 460772
rect 418982 460536 419066 460772
rect 419302 460536 419334 460772
rect 418714 455454 419334 460536
rect 418714 455218 418746 455454
rect 418982 455218 419066 455454
rect 419302 455218 419334 455454
rect 418714 455134 419334 455218
rect 418714 454898 418746 455134
rect 418982 454898 419066 455134
rect 419302 454898 419334 455134
rect 418714 437454 419334 454898
rect 418714 437218 418746 437454
rect 418982 437218 419066 437454
rect 419302 437218 419334 437454
rect 418714 437134 419334 437218
rect 418714 436898 418746 437134
rect 418982 436898 419066 437134
rect 419302 436898 419334 437134
rect 418714 419454 419334 436898
rect 418714 419218 418746 419454
rect 418982 419218 419066 419454
rect 419302 419218 419334 419454
rect 418714 419134 419334 419218
rect 418714 418898 418746 419134
rect 418982 418898 419066 419134
rect 419302 418898 419334 419134
rect 418714 401454 419334 418898
rect 418714 401218 418746 401454
rect 418982 401218 419066 401454
rect 419302 401218 419334 401454
rect 418714 401134 419334 401218
rect 418714 400898 418746 401134
rect 418982 400898 419066 401134
rect 419302 400898 419334 401134
rect 418714 383454 419334 400898
rect 418714 383218 418746 383454
rect 418982 383218 419066 383454
rect 419302 383218 419334 383454
rect 418714 383134 419334 383218
rect 418714 382898 418746 383134
rect 418982 382898 419066 383134
rect 419302 382898 419334 383134
rect 418714 365454 419334 382898
rect 418714 365218 418746 365454
rect 418982 365218 419066 365454
rect 419302 365218 419334 365454
rect 418714 365134 419334 365218
rect 418714 364898 418746 365134
rect 418982 364898 419066 365134
rect 419302 364898 419334 365134
rect 418714 347454 419334 364898
rect 418714 347218 418746 347454
rect 418982 347218 419066 347454
rect 419302 347218 419334 347454
rect 418714 347134 419334 347218
rect 418714 346898 418746 347134
rect 418982 346898 419066 347134
rect 419302 346898 419334 347134
rect 418714 329454 419334 346898
rect 418714 329218 418746 329454
rect 418982 329218 419066 329454
rect 419302 329218 419334 329454
rect 418714 329134 419334 329218
rect 418714 328898 418746 329134
rect 418982 328898 419066 329134
rect 419302 328898 419334 329134
rect 418714 311454 419334 328898
rect 418714 311218 418746 311454
rect 418982 311218 419066 311454
rect 419302 311218 419334 311454
rect 418714 311134 419334 311218
rect 418714 310898 418746 311134
rect 418982 310898 419066 311134
rect 419302 310898 419334 311134
rect 418714 293454 419334 310898
rect 418714 293218 418746 293454
rect 418982 293218 419066 293454
rect 419302 293218 419334 293454
rect 418714 293134 419334 293218
rect 418714 292898 418746 293134
rect 418982 292898 419066 293134
rect 419302 292898 419334 293134
rect 418714 275454 419334 292898
rect 418714 275218 418746 275454
rect 418982 275218 419066 275454
rect 419302 275218 419334 275454
rect 418714 275134 419334 275218
rect 418714 274898 418746 275134
rect 418982 274898 419066 275134
rect 419302 274898 419334 275134
rect 418714 257454 419334 274898
rect 418714 257218 418746 257454
rect 418982 257218 419066 257454
rect 419302 257218 419334 257454
rect 418714 257134 419334 257218
rect 418714 256898 418746 257134
rect 418982 256898 419066 257134
rect 419302 256898 419334 257134
rect 418714 239454 419334 256898
rect 418714 239218 418746 239454
rect 418982 239218 419066 239454
rect 419302 239218 419334 239454
rect 418714 239134 419334 239218
rect 418714 238898 418746 239134
rect 418982 238898 419066 239134
rect 419302 238898 419334 239134
rect 418714 221454 419334 238898
rect 418714 221218 418746 221454
rect 418982 221218 419066 221454
rect 419302 221218 419334 221454
rect 418714 221134 419334 221218
rect 418714 220898 418746 221134
rect 418982 220898 419066 221134
rect 419302 220898 419334 221134
rect 418714 203454 419334 220898
rect 418714 203218 418746 203454
rect 418982 203218 419066 203454
rect 419302 203218 419334 203454
rect 418714 203134 419334 203218
rect 418714 202898 418746 203134
rect 418982 202898 419066 203134
rect 419302 202898 419334 203134
rect 418714 185454 419334 202898
rect 418714 185218 418746 185454
rect 418982 185218 419066 185454
rect 419302 185218 419334 185454
rect 418714 185134 419334 185218
rect 418714 184898 418746 185134
rect 418982 184898 419066 185134
rect 419302 184898 419334 185134
rect 418714 167454 419334 184898
rect 418714 167218 418746 167454
rect 418982 167218 419066 167454
rect 419302 167218 419334 167454
rect 418714 167134 419334 167218
rect 418714 166898 418746 167134
rect 418982 166898 419066 167134
rect 419302 166898 419334 167134
rect 418714 149454 419334 166898
rect 418714 149218 418746 149454
rect 418982 149218 419066 149454
rect 419302 149218 419334 149454
rect 418714 149134 419334 149218
rect 418714 148898 418746 149134
rect 418982 148898 419066 149134
rect 419302 148898 419334 149134
rect 418714 131454 419334 148898
rect 418714 131218 418746 131454
rect 418982 131218 419066 131454
rect 419302 131218 419334 131454
rect 418714 131134 419334 131218
rect 418714 130898 418746 131134
rect 418982 130898 419066 131134
rect 419302 130898 419334 131134
rect 418714 113454 419334 130898
rect 418714 113218 418746 113454
rect 418982 113218 419066 113454
rect 419302 113218 419334 113454
rect 418714 113134 419334 113218
rect 418714 112898 418746 113134
rect 418982 112898 419066 113134
rect 419302 112898 419334 113134
rect 418714 95454 419334 112898
rect 418714 95218 418746 95454
rect 418982 95218 419066 95454
rect 419302 95218 419334 95454
rect 418714 95134 419334 95218
rect 418714 94898 418746 95134
rect 418982 94898 419066 95134
rect 419302 94898 419334 95134
rect 418714 77454 419334 94898
rect 418714 77218 418746 77454
rect 418982 77218 419066 77454
rect 419302 77218 419334 77454
rect 418714 77134 419334 77218
rect 418714 76898 418746 77134
rect 418982 76898 419066 77134
rect 419302 76898 419334 77134
rect 418714 59454 419334 76898
rect 418714 59218 418746 59454
rect 418982 59218 419066 59454
rect 419302 59218 419334 59454
rect 418714 59134 419334 59218
rect 418714 58898 418746 59134
rect 418982 58898 419066 59134
rect 419302 58898 419334 59134
rect 418714 41454 419334 58898
rect 418714 41218 418746 41454
rect 418982 41218 419066 41454
rect 419302 41218 419334 41454
rect 418714 41134 419334 41218
rect 418714 40898 418746 41134
rect 418982 40898 419066 41134
rect 419302 40898 419334 41134
rect 418714 23454 419334 40898
rect 418714 23218 418746 23454
rect 418982 23218 419066 23454
rect 419302 23218 419334 23454
rect 418714 23134 419334 23218
rect 418714 22898 418746 23134
rect 418982 22898 419066 23134
rect 419302 22898 419334 23134
rect 418714 5454 419334 22898
rect 418714 5218 418746 5454
rect 418982 5218 419066 5454
rect 419302 5218 419334 5454
rect 418714 5134 419334 5218
rect 418714 4898 418746 5134
rect 418982 4898 419066 5134
rect 419302 4898 419334 5134
rect 418714 -856 419334 4898
rect 418714 -1092 418746 -856
rect 418982 -1092 419066 -856
rect 419302 -1092 419334 -856
rect 418714 -1176 419334 -1092
rect 418714 -1412 418746 -1176
rect 418982 -1412 419066 -1176
rect 419302 -1412 419334 -1176
rect 418714 -4324 419334 -1412
rect 422434 462052 423054 464004
rect 422434 461816 422466 462052
rect 422702 461816 422786 462052
rect 423022 461816 423054 462052
rect 422434 461732 423054 461816
rect 422434 461496 422466 461732
rect 422702 461496 422786 461732
rect 423022 461496 423054 461732
rect 422434 441174 423054 461496
rect 422434 440938 422466 441174
rect 422702 440938 422786 441174
rect 423022 440938 423054 441174
rect 422434 440854 423054 440938
rect 422434 440618 422466 440854
rect 422702 440618 422786 440854
rect 423022 440618 423054 440854
rect 422434 423174 423054 440618
rect 422434 422938 422466 423174
rect 422702 422938 422786 423174
rect 423022 422938 423054 423174
rect 422434 422854 423054 422938
rect 422434 422618 422466 422854
rect 422702 422618 422786 422854
rect 423022 422618 423054 422854
rect 422434 405174 423054 422618
rect 422434 404938 422466 405174
rect 422702 404938 422786 405174
rect 423022 404938 423054 405174
rect 422434 404854 423054 404938
rect 422434 404618 422466 404854
rect 422702 404618 422786 404854
rect 423022 404618 423054 404854
rect 422434 387174 423054 404618
rect 422434 386938 422466 387174
rect 422702 386938 422786 387174
rect 423022 386938 423054 387174
rect 422434 386854 423054 386938
rect 422434 386618 422466 386854
rect 422702 386618 422786 386854
rect 423022 386618 423054 386854
rect 422434 369174 423054 386618
rect 422434 368938 422466 369174
rect 422702 368938 422786 369174
rect 423022 368938 423054 369174
rect 422434 368854 423054 368938
rect 422434 368618 422466 368854
rect 422702 368618 422786 368854
rect 423022 368618 423054 368854
rect 422434 351174 423054 368618
rect 422434 350938 422466 351174
rect 422702 350938 422786 351174
rect 423022 350938 423054 351174
rect 422434 350854 423054 350938
rect 422434 350618 422466 350854
rect 422702 350618 422786 350854
rect 423022 350618 423054 350854
rect 422434 333174 423054 350618
rect 422434 332938 422466 333174
rect 422702 332938 422786 333174
rect 423022 332938 423054 333174
rect 422434 332854 423054 332938
rect 422434 332618 422466 332854
rect 422702 332618 422786 332854
rect 423022 332618 423054 332854
rect 422434 315174 423054 332618
rect 422434 314938 422466 315174
rect 422702 314938 422786 315174
rect 423022 314938 423054 315174
rect 422434 314854 423054 314938
rect 422434 314618 422466 314854
rect 422702 314618 422786 314854
rect 423022 314618 423054 314854
rect 422434 297174 423054 314618
rect 422434 296938 422466 297174
rect 422702 296938 422786 297174
rect 423022 296938 423054 297174
rect 422434 296854 423054 296938
rect 422434 296618 422466 296854
rect 422702 296618 422786 296854
rect 423022 296618 423054 296854
rect 422434 279174 423054 296618
rect 422434 278938 422466 279174
rect 422702 278938 422786 279174
rect 423022 278938 423054 279174
rect 422434 278854 423054 278938
rect 422434 278618 422466 278854
rect 422702 278618 422786 278854
rect 423022 278618 423054 278854
rect 422434 261174 423054 278618
rect 422434 260938 422466 261174
rect 422702 260938 422786 261174
rect 423022 260938 423054 261174
rect 422434 260854 423054 260938
rect 422434 260618 422466 260854
rect 422702 260618 422786 260854
rect 423022 260618 423054 260854
rect 422434 243174 423054 260618
rect 422434 242938 422466 243174
rect 422702 242938 422786 243174
rect 423022 242938 423054 243174
rect 422434 242854 423054 242938
rect 422434 242618 422466 242854
rect 422702 242618 422786 242854
rect 423022 242618 423054 242854
rect 422434 225174 423054 242618
rect 422434 224938 422466 225174
rect 422702 224938 422786 225174
rect 423022 224938 423054 225174
rect 422434 224854 423054 224938
rect 422434 224618 422466 224854
rect 422702 224618 422786 224854
rect 423022 224618 423054 224854
rect 422434 207174 423054 224618
rect 422434 206938 422466 207174
rect 422702 206938 422786 207174
rect 423022 206938 423054 207174
rect 422434 206854 423054 206938
rect 422434 206618 422466 206854
rect 422702 206618 422786 206854
rect 423022 206618 423054 206854
rect 422434 189174 423054 206618
rect 422434 188938 422466 189174
rect 422702 188938 422786 189174
rect 423022 188938 423054 189174
rect 422434 188854 423054 188938
rect 422434 188618 422466 188854
rect 422702 188618 422786 188854
rect 423022 188618 423054 188854
rect 422434 171174 423054 188618
rect 422434 170938 422466 171174
rect 422702 170938 422786 171174
rect 423022 170938 423054 171174
rect 422434 170854 423054 170938
rect 422434 170618 422466 170854
rect 422702 170618 422786 170854
rect 423022 170618 423054 170854
rect 422434 153174 423054 170618
rect 422434 152938 422466 153174
rect 422702 152938 422786 153174
rect 423022 152938 423054 153174
rect 422434 152854 423054 152938
rect 422434 152618 422466 152854
rect 422702 152618 422786 152854
rect 423022 152618 423054 152854
rect 422434 135174 423054 152618
rect 422434 134938 422466 135174
rect 422702 134938 422786 135174
rect 423022 134938 423054 135174
rect 422434 134854 423054 134938
rect 422434 134618 422466 134854
rect 422702 134618 422786 134854
rect 423022 134618 423054 134854
rect 422434 117174 423054 134618
rect 422434 116938 422466 117174
rect 422702 116938 422786 117174
rect 423022 116938 423054 117174
rect 422434 116854 423054 116938
rect 422434 116618 422466 116854
rect 422702 116618 422786 116854
rect 423022 116618 423054 116854
rect 422434 99174 423054 116618
rect 422434 98938 422466 99174
rect 422702 98938 422786 99174
rect 423022 98938 423054 99174
rect 422434 98854 423054 98938
rect 422434 98618 422466 98854
rect 422702 98618 422786 98854
rect 423022 98618 423054 98854
rect 422434 81174 423054 98618
rect 422434 80938 422466 81174
rect 422702 80938 422786 81174
rect 423022 80938 423054 81174
rect 422434 80854 423054 80938
rect 422434 80618 422466 80854
rect 422702 80618 422786 80854
rect 423022 80618 423054 80854
rect 422434 63174 423054 80618
rect 422434 62938 422466 63174
rect 422702 62938 422786 63174
rect 423022 62938 423054 63174
rect 422434 62854 423054 62938
rect 422434 62618 422466 62854
rect 422702 62618 422786 62854
rect 423022 62618 423054 62854
rect 422434 45174 423054 62618
rect 422434 44938 422466 45174
rect 422702 44938 422786 45174
rect 423022 44938 423054 45174
rect 422434 44854 423054 44938
rect 422434 44618 422466 44854
rect 422702 44618 422786 44854
rect 423022 44618 423054 44854
rect 422434 27174 423054 44618
rect 422434 26938 422466 27174
rect 422702 26938 422786 27174
rect 423022 26938 423054 27174
rect 422434 26854 423054 26938
rect 422434 26618 422466 26854
rect 422702 26618 422786 26854
rect 423022 26618 423054 26854
rect 422434 9174 423054 26618
rect 422434 8938 422466 9174
rect 422702 8938 422786 9174
rect 423022 8938 423054 9174
rect 422434 8854 423054 8938
rect 422434 8618 422466 8854
rect 422702 8618 422786 8854
rect 423022 8618 423054 8854
rect 422434 -1816 423054 8618
rect 422434 -2052 422466 -1816
rect 422702 -2052 422786 -1816
rect 423022 -2052 423054 -1816
rect 422434 -2136 423054 -2052
rect 422434 -2372 422466 -2136
rect 422702 -2372 422786 -2136
rect 423022 -2372 423054 -2136
rect 422434 -4324 423054 -2372
rect 426154 463012 426774 464004
rect 426154 462776 426186 463012
rect 426422 462776 426506 463012
rect 426742 462776 426774 463012
rect 426154 462692 426774 462776
rect 426154 462456 426186 462692
rect 426422 462456 426506 462692
rect 426742 462456 426774 462692
rect 426154 444894 426774 462456
rect 426154 444658 426186 444894
rect 426422 444658 426506 444894
rect 426742 444658 426774 444894
rect 426154 444574 426774 444658
rect 426154 444338 426186 444574
rect 426422 444338 426506 444574
rect 426742 444338 426774 444574
rect 426154 426894 426774 444338
rect 426154 426658 426186 426894
rect 426422 426658 426506 426894
rect 426742 426658 426774 426894
rect 426154 426574 426774 426658
rect 426154 426338 426186 426574
rect 426422 426338 426506 426574
rect 426742 426338 426774 426574
rect 426154 408894 426774 426338
rect 426154 408658 426186 408894
rect 426422 408658 426506 408894
rect 426742 408658 426774 408894
rect 426154 408574 426774 408658
rect 426154 408338 426186 408574
rect 426422 408338 426506 408574
rect 426742 408338 426774 408574
rect 426154 390894 426774 408338
rect 426154 390658 426186 390894
rect 426422 390658 426506 390894
rect 426742 390658 426774 390894
rect 426154 390574 426774 390658
rect 426154 390338 426186 390574
rect 426422 390338 426506 390574
rect 426742 390338 426774 390574
rect 426154 372894 426774 390338
rect 426154 372658 426186 372894
rect 426422 372658 426506 372894
rect 426742 372658 426774 372894
rect 426154 372574 426774 372658
rect 426154 372338 426186 372574
rect 426422 372338 426506 372574
rect 426742 372338 426774 372574
rect 426154 354894 426774 372338
rect 426154 354658 426186 354894
rect 426422 354658 426506 354894
rect 426742 354658 426774 354894
rect 426154 354574 426774 354658
rect 426154 354338 426186 354574
rect 426422 354338 426506 354574
rect 426742 354338 426774 354574
rect 426154 336894 426774 354338
rect 426154 336658 426186 336894
rect 426422 336658 426506 336894
rect 426742 336658 426774 336894
rect 426154 336574 426774 336658
rect 426154 336338 426186 336574
rect 426422 336338 426506 336574
rect 426742 336338 426774 336574
rect 426154 318894 426774 336338
rect 426154 318658 426186 318894
rect 426422 318658 426506 318894
rect 426742 318658 426774 318894
rect 426154 318574 426774 318658
rect 426154 318338 426186 318574
rect 426422 318338 426506 318574
rect 426742 318338 426774 318574
rect 426154 300894 426774 318338
rect 426154 300658 426186 300894
rect 426422 300658 426506 300894
rect 426742 300658 426774 300894
rect 426154 300574 426774 300658
rect 426154 300338 426186 300574
rect 426422 300338 426506 300574
rect 426742 300338 426774 300574
rect 426154 282894 426774 300338
rect 426154 282658 426186 282894
rect 426422 282658 426506 282894
rect 426742 282658 426774 282894
rect 426154 282574 426774 282658
rect 426154 282338 426186 282574
rect 426422 282338 426506 282574
rect 426742 282338 426774 282574
rect 426154 264894 426774 282338
rect 426154 264658 426186 264894
rect 426422 264658 426506 264894
rect 426742 264658 426774 264894
rect 426154 264574 426774 264658
rect 426154 264338 426186 264574
rect 426422 264338 426506 264574
rect 426742 264338 426774 264574
rect 426154 246894 426774 264338
rect 426154 246658 426186 246894
rect 426422 246658 426506 246894
rect 426742 246658 426774 246894
rect 426154 246574 426774 246658
rect 426154 246338 426186 246574
rect 426422 246338 426506 246574
rect 426742 246338 426774 246574
rect 426154 228894 426774 246338
rect 426154 228658 426186 228894
rect 426422 228658 426506 228894
rect 426742 228658 426774 228894
rect 426154 228574 426774 228658
rect 426154 228338 426186 228574
rect 426422 228338 426506 228574
rect 426742 228338 426774 228574
rect 426154 210894 426774 228338
rect 426154 210658 426186 210894
rect 426422 210658 426506 210894
rect 426742 210658 426774 210894
rect 426154 210574 426774 210658
rect 426154 210338 426186 210574
rect 426422 210338 426506 210574
rect 426742 210338 426774 210574
rect 426154 192894 426774 210338
rect 426154 192658 426186 192894
rect 426422 192658 426506 192894
rect 426742 192658 426774 192894
rect 426154 192574 426774 192658
rect 426154 192338 426186 192574
rect 426422 192338 426506 192574
rect 426742 192338 426774 192574
rect 426154 174894 426774 192338
rect 426154 174658 426186 174894
rect 426422 174658 426506 174894
rect 426742 174658 426774 174894
rect 426154 174574 426774 174658
rect 426154 174338 426186 174574
rect 426422 174338 426506 174574
rect 426742 174338 426774 174574
rect 426154 156894 426774 174338
rect 426154 156658 426186 156894
rect 426422 156658 426506 156894
rect 426742 156658 426774 156894
rect 426154 156574 426774 156658
rect 426154 156338 426186 156574
rect 426422 156338 426506 156574
rect 426742 156338 426774 156574
rect 426154 138894 426774 156338
rect 426154 138658 426186 138894
rect 426422 138658 426506 138894
rect 426742 138658 426774 138894
rect 426154 138574 426774 138658
rect 426154 138338 426186 138574
rect 426422 138338 426506 138574
rect 426742 138338 426774 138574
rect 426154 120894 426774 138338
rect 426154 120658 426186 120894
rect 426422 120658 426506 120894
rect 426742 120658 426774 120894
rect 426154 120574 426774 120658
rect 426154 120338 426186 120574
rect 426422 120338 426506 120574
rect 426742 120338 426774 120574
rect 426154 102894 426774 120338
rect 426154 102658 426186 102894
rect 426422 102658 426506 102894
rect 426742 102658 426774 102894
rect 426154 102574 426774 102658
rect 426154 102338 426186 102574
rect 426422 102338 426506 102574
rect 426742 102338 426774 102574
rect 426154 84894 426774 102338
rect 426154 84658 426186 84894
rect 426422 84658 426506 84894
rect 426742 84658 426774 84894
rect 426154 84574 426774 84658
rect 426154 84338 426186 84574
rect 426422 84338 426506 84574
rect 426742 84338 426774 84574
rect 426154 66894 426774 84338
rect 426154 66658 426186 66894
rect 426422 66658 426506 66894
rect 426742 66658 426774 66894
rect 426154 66574 426774 66658
rect 426154 66338 426186 66574
rect 426422 66338 426506 66574
rect 426742 66338 426774 66574
rect 426154 48894 426774 66338
rect 426154 48658 426186 48894
rect 426422 48658 426506 48894
rect 426742 48658 426774 48894
rect 426154 48574 426774 48658
rect 426154 48338 426186 48574
rect 426422 48338 426506 48574
rect 426742 48338 426774 48574
rect 426154 30894 426774 48338
rect 426154 30658 426186 30894
rect 426422 30658 426506 30894
rect 426742 30658 426774 30894
rect 426154 30574 426774 30658
rect 426154 30338 426186 30574
rect 426422 30338 426506 30574
rect 426742 30338 426774 30574
rect 426154 12894 426774 30338
rect 426154 12658 426186 12894
rect 426422 12658 426506 12894
rect 426742 12658 426774 12894
rect 426154 12574 426774 12658
rect 426154 12338 426186 12574
rect 426422 12338 426506 12574
rect 426742 12338 426774 12574
rect 426154 -2776 426774 12338
rect 426154 -3012 426186 -2776
rect 426422 -3012 426506 -2776
rect 426742 -3012 426774 -2776
rect 426154 -3096 426774 -3012
rect 426154 -3332 426186 -3096
rect 426422 -3332 426506 -3096
rect 426742 -3332 426774 -3096
rect 426154 -4324 426774 -3332
rect 429874 463972 430494 464004
rect 429874 463736 429906 463972
rect 430142 463736 430226 463972
rect 430462 463736 430494 463972
rect 429874 463652 430494 463736
rect 429874 463416 429906 463652
rect 430142 463416 430226 463652
rect 430462 463416 430494 463652
rect 429874 448614 430494 463416
rect 429874 448378 429906 448614
rect 430142 448378 430226 448614
rect 430462 448378 430494 448614
rect 429874 448294 430494 448378
rect 429874 448058 429906 448294
rect 430142 448058 430226 448294
rect 430462 448058 430494 448294
rect 429874 430614 430494 448058
rect 429874 430378 429906 430614
rect 430142 430378 430226 430614
rect 430462 430378 430494 430614
rect 429874 430294 430494 430378
rect 429874 430058 429906 430294
rect 430142 430058 430226 430294
rect 430462 430058 430494 430294
rect 429874 412614 430494 430058
rect 429874 412378 429906 412614
rect 430142 412378 430226 412614
rect 430462 412378 430494 412614
rect 429874 412294 430494 412378
rect 429874 412058 429906 412294
rect 430142 412058 430226 412294
rect 430462 412058 430494 412294
rect 429874 394614 430494 412058
rect 429874 394378 429906 394614
rect 430142 394378 430226 394614
rect 430462 394378 430494 394614
rect 429874 394294 430494 394378
rect 429874 394058 429906 394294
rect 430142 394058 430226 394294
rect 430462 394058 430494 394294
rect 429874 376614 430494 394058
rect 429874 376378 429906 376614
rect 430142 376378 430226 376614
rect 430462 376378 430494 376614
rect 429874 376294 430494 376378
rect 429874 376058 429906 376294
rect 430142 376058 430226 376294
rect 430462 376058 430494 376294
rect 429874 358614 430494 376058
rect 429874 358378 429906 358614
rect 430142 358378 430226 358614
rect 430462 358378 430494 358614
rect 429874 358294 430494 358378
rect 429874 358058 429906 358294
rect 430142 358058 430226 358294
rect 430462 358058 430494 358294
rect 429874 340614 430494 358058
rect 429874 340378 429906 340614
rect 430142 340378 430226 340614
rect 430462 340378 430494 340614
rect 429874 340294 430494 340378
rect 429874 340058 429906 340294
rect 430142 340058 430226 340294
rect 430462 340058 430494 340294
rect 429874 322614 430494 340058
rect 429874 322378 429906 322614
rect 430142 322378 430226 322614
rect 430462 322378 430494 322614
rect 429874 322294 430494 322378
rect 429874 322058 429906 322294
rect 430142 322058 430226 322294
rect 430462 322058 430494 322294
rect 429874 304614 430494 322058
rect 429874 304378 429906 304614
rect 430142 304378 430226 304614
rect 430462 304378 430494 304614
rect 429874 304294 430494 304378
rect 429874 304058 429906 304294
rect 430142 304058 430226 304294
rect 430462 304058 430494 304294
rect 429874 286614 430494 304058
rect 429874 286378 429906 286614
rect 430142 286378 430226 286614
rect 430462 286378 430494 286614
rect 429874 286294 430494 286378
rect 429874 286058 429906 286294
rect 430142 286058 430226 286294
rect 430462 286058 430494 286294
rect 429874 268614 430494 286058
rect 429874 268378 429906 268614
rect 430142 268378 430226 268614
rect 430462 268378 430494 268614
rect 429874 268294 430494 268378
rect 429874 268058 429906 268294
rect 430142 268058 430226 268294
rect 430462 268058 430494 268294
rect 429874 250614 430494 268058
rect 429874 250378 429906 250614
rect 430142 250378 430226 250614
rect 430462 250378 430494 250614
rect 429874 250294 430494 250378
rect 429874 250058 429906 250294
rect 430142 250058 430226 250294
rect 430462 250058 430494 250294
rect 429874 232614 430494 250058
rect 429874 232378 429906 232614
rect 430142 232378 430226 232614
rect 430462 232378 430494 232614
rect 429874 232294 430494 232378
rect 429874 232058 429906 232294
rect 430142 232058 430226 232294
rect 430462 232058 430494 232294
rect 429874 214614 430494 232058
rect 429874 214378 429906 214614
rect 430142 214378 430226 214614
rect 430462 214378 430494 214614
rect 429874 214294 430494 214378
rect 429874 214058 429906 214294
rect 430142 214058 430226 214294
rect 430462 214058 430494 214294
rect 429874 196614 430494 214058
rect 429874 196378 429906 196614
rect 430142 196378 430226 196614
rect 430462 196378 430494 196614
rect 429874 196294 430494 196378
rect 429874 196058 429906 196294
rect 430142 196058 430226 196294
rect 430462 196058 430494 196294
rect 429874 178614 430494 196058
rect 429874 178378 429906 178614
rect 430142 178378 430226 178614
rect 430462 178378 430494 178614
rect 429874 178294 430494 178378
rect 429874 178058 429906 178294
rect 430142 178058 430226 178294
rect 430462 178058 430494 178294
rect 429874 160614 430494 178058
rect 429874 160378 429906 160614
rect 430142 160378 430226 160614
rect 430462 160378 430494 160614
rect 429874 160294 430494 160378
rect 429874 160058 429906 160294
rect 430142 160058 430226 160294
rect 430462 160058 430494 160294
rect 429874 142614 430494 160058
rect 429874 142378 429906 142614
rect 430142 142378 430226 142614
rect 430462 142378 430494 142614
rect 429874 142294 430494 142378
rect 429874 142058 429906 142294
rect 430142 142058 430226 142294
rect 430462 142058 430494 142294
rect 429874 124614 430494 142058
rect 429874 124378 429906 124614
rect 430142 124378 430226 124614
rect 430462 124378 430494 124614
rect 429874 124294 430494 124378
rect 429874 124058 429906 124294
rect 430142 124058 430226 124294
rect 430462 124058 430494 124294
rect 429874 106614 430494 124058
rect 429874 106378 429906 106614
rect 430142 106378 430226 106614
rect 430462 106378 430494 106614
rect 429874 106294 430494 106378
rect 429874 106058 429906 106294
rect 430142 106058 430226 106294
rect 430462 106058 430494 106294
rect 429874 88614 430494 106058
rect 429874 88378 429906 88614
rect 430142 88378 430226 88614
rect 430462 88378 430494 88614
rect 429874 88294 430494 88378
rect 429874 88058 429906 88294
rect 430142 88058 430226 88294
rect 430462 88058 430494 88294
rect 429874 70614 430494 88058
rect 429874 70378 429906 70614
rect 430142 70378 430226 70614
rect 430462 70378 430494 70614
rect 429874 70294 430494 70378
rect 429874 70058 429906 70294
rect 430142 70058 430226 70294
rect 430462 70058 430494 70294
rect 429874 52614 430494 70058
rect 429874 52378 429906 52614
rect 430142 52378 430226 52614
rect 430462 52378 430494 52614
rect 429874 52294 430494 52378
rect 429874 52058 429906 52294
rect 430142 52058 430226 52294
rect 430462 52058 430494 52294
rect 429874 34614 430494 52058
rect 429874 34378 429906 34614
rect 430142 34378 430226 34614
rect 430462 34378 430494 34614
rect 429874 34294 430494 34378
rect 429874 34058 429906 34294
rect 430142 34058 430226 34294
rect 430462 34058 430494 34294
rect 429874 16614 430494 34058
rect 429874 16378 429906 16614
rect 430142 16378 430226 16614
rect 430462 16378 430494 16614
rect 429874 16294 430494 16378
rect 429874 16058 429906 16294
rect 430142 16058 430226 16294
rect 430462 16058 430494 16294
rect 429874 -3736 430494 16058
rect 429874 -3972 429906 -3736
rect 430142 -3972 430226 -3736
rect 430462 -3972 430494 -3736
rect 429874 -4056 430494 -3972
rect 429874 -4292 429906 -4056
rect 430142 -4292 430226 -4056
rect 430462 -4292 430494 -4056
rect 429874 -4324 430494 -4292
rect 436714 461092 437334 464004
rect 436714 460856 436746 461092
rect 436982 460856 437066 461092
rect 437302 460856 437334 461092
rect 436714 460772 437334 460856
rect 436714 460536 436746 460772
rect 436982 460536 437066 460772
rect 437302 460536 437334 460772
rect 436714 455454 437334 460536
rect 436714 455218 436746 455454
rect 436982 455218 437066 455454
rect 437302 455218 437334 455454
rect 436714 455134 437334 455218
rect 436714 454898 436746 455134
rect 436982 454898 437066 455134
rect 437302 454898 437334 455134
rect 436714 437454 437334 454898
rect 436714 437218 436746 437454
rect 436982 437218 437066 437454
rect 437302 437218 437334 437454
rect 436714 437134 437334 437218
rect 436714 436898 436746 437134
rect 436982 436898 437066 437134
rect 437302 436898 437334 437134
rect 436714 419454 437334 436898
rect 436714 419218 436746 419454
rect 436982 419218 437066 419454
rect 437302 419218 437334 419454
rect 436714 419134 437334 419218
rect 436714 418898 436746 419134
rect 436982 418898 437066 419134
rect 437302 418898 437334 419134
rect 436714 401454 437334 418898
rect 436714 401218 436746 401454
rect 436982 401218 437066 401454
rect 437302 401218 437334 401454
rect 436714 401134 437334 401218
rect 436714 400898 436746 401134
rect 436982 400898 437066 401134
rect 437302 400898 437334 401134
rect 436714 383454 437334 400898
rect 436714 383218 436746 383454
rect 436982 383218 437066 383454
rect 437302 383218 437334 383454
rect 436714 383134 437334 383218
rect 436714 382898 436746 383134
rect 436982 382898 437066 383134
rect 437302 382898 437334 383134
rect 436714 365454 437334 382898
rect 436714 365218 436746 365454
rect 436982 365218 437066 365454
rect 437302 365218 437334 365454
rect 436714 365134 437334 365218
rect 436714 364898 436746 365134
rect 436982 364898 437066 365134
rect 437302 364898 437334 365134
rect 436714 347454 437334 364898
rect 436714 347218 436746 347454
rect 436982 347218 437066 347454
rect 437302 347218 437334 347454
rect 436714 347134 437334 347218
rect 436714 346898 436746 347134
rect 436982 346898 437066 347134
rect 437302 346898 437334 347134
rect 436714 329454 437334 346898
rect 436714 329218 436746 329454
rect 436982 329218 437066 329454
rect 437302 329218 437334 329454
rect 436714 329134 437334 329218
rect 436714 328898 436746 329134
rect 436982 328898 437066 329134
rect 437302 328898 437334 329134
rect 436714 311454 437334 328898
rect 436714 311218 436746 311454
rect 436982 311218 437066 311454
rect 437302 311218 437334 311454
rect 436714 311134 437334 311218
rect 436714 310898 436746 311134
rect 436982 310898 437066 311134
rect 437302 310898 437334 311134
rect 436714 293454 437334 310898
rect 436714 293218 436746 293454
rect 436982 293218 437066 293454
rect 437302 293218 437334 293454
rect 436714 293134 437334 293218
rect 436714 292898 436746 293134
rect 436982 292898 437066 293134
rect 437302 292898 437334 293134
rect 436714 275454 437334 292898
rect 436714 275218 436746 275454
rect 436982 275218 437066 275454
rect 437302 275218 437334 275454
rect 436714 275134 437334 275218
rect 436714 274898 436746 275134
rect 436982 274898 437066 275134
rect 437302 274898 437334 275134
rect 436714 257454 437334 274898
rect 436714 257218 436746 257454
rect 436982 257218 437066 257454
rect 437302 257218 437334 257454
rect 436714 257134 437334 257218
rect 436714 256898 436746 257134
rect 436982 256898 437066 257134
rect 437302 256898 437334 257134
rect 436714 239454 437334 256898
rect 436714 239218 436746 239454
rect 436982 239218 437066 239454
rect 437302 239218 437334 239454
rect 436714 239134 437334 239218
rect 436714 238898 436746 239134
rect 436982 238898 437066 239134
rect 437302 238898 437334 239134
rect 436714 221454 437334 238898
rect 436714 221218 436746 221454
rect 436982 221218 437066 221454
rect 437302 221218 437334 221454
rect 436714 221134 437334 221218
rect 436714 220898 436746 221134
rect 436982 220898 437066 221134
rect 437302 220898 437334 221134
rect 436714 203454 437334 220898
rect 436714 203218 436746 203454
rect 436982 203218 437066 203454
rect 437302 203218 437334 203454
rect 436714 203134 437334 203218
rect 436714 202898 436746 203134
rect 436982 202898 437066 203134
rect 437302 202898 437334 203134
rect 436714 185454 437334 202898
rect 436714 185218 436746 185454
rect 436982 185218 437066 185454
rect 437302 185218 437334 185454
rect 436714 185134 437334 185218
rect 436714 184898 436746 185134
rect 436982 184898 437066 185134
rect 437302 184898 437334 185134
rect 436714 167454 437334 184898
rect 436714 167218 436746 167454
rect 436982 167218 437066 167454
rect 437302 167218 437334 167454
rect 436714 167134 437334 167218
rect 436714 166898 436746 167134
rect 436982 166898 437066 167134
rect 437302 166898 437334 167134
rect 436714 149454 437334 166898
rect 436714 149218 436746 149454
rect 436982 149218 437066 149454
rect 437302 149218 437334 149454
rect 436714 149134 437334 149218
rect 436714 148898 436746 149134
rect 436982 148898 437066 149134
rect 437302 148898 437334 149134
rect 436714 131454 437334 148898
rect 436714 131218 436746 131454
rect 436982 131218 437066 131454
rect 437302 131218 437334 131454
rect 436714 131134 437334 131218
rect 436714 130898 436746 131134
rect 436982 130898 437066 131134
rect 437302 130898 437334 131134
rect 436714 113454 437334 130898
rect 436714 113218 436746 113454
rect 436982 113218 437066 113454
rect 437302 113218 437334 113454
rect 436714 113134 437334 113218
rect 436714 112898 436746 113134
rect 436982 112898 437066 113134
rect 437302 112898 437334 113134
rect 436714 95454 437334 112898
rect 436714 95218 436746 95454
rect 436982 95218 437066 95454
rect 437302 95218 437334 95454
rect 436714 95134 437334 95218
rect 436714 94898 436746 95134
rect 436982 94898 437066 95134
rect 437302 94898 437334 95134
rect 436714 77454 437334 94898
rect 436714 77218 436746 77454
rect 436982 77218 437066 77454
rect 437302 77218 437334 77454
rect 436714 77134 437334 77218
rect 436714 76898 436746 77134
rect 436982 76898 437066 77134
rect 437302 76898 437334 77134
rect 436714 59454 437334 76898
rect 436714 59218 436746 59454
rect 436982 59218 437066 59454
rect 437302 59218 437334 59454
rect 436714 59134 437334 59218
rect 436714 58898 436746 59134
rect 436982 58898 437066 59134
rect 437302 58898 437334 59134
rect 436714 41454 437334 58898
rect 436714 41218 436746 41454
rect 436982 41218 437066 41454
rect 437302 41218 437334 41454
rect 436714 41134 437334 41218
rect 436714 40898 436746 41134
rect 436982 40898 437066 41134
rect 437302 40898 437334 41134
rect 436714 23454 437334 40898
rect 436714 23218 436746 23454
rect 436982 23218 437066 23454
rect 437302 23218 437334 23454
rect 436714 23134 437334 23218
rect 436714 22898 436746 23134
rect 436982 22898 437066 23134
rect 437302 22898 437334 23134
rect 436714 5454 437334 22898
rect 436714 5218 436746 5454
rect 436982 5218 437066 5454
rect 437302 5218 437334 5454
rect 436714 5134 437334 5218
rect 436714 4898 436746 5134
rect 436982 4898 437066 5134
rect 437302 4898 437334 5134
rect 436714 -856 437334 4898
rect 436714 -1092 436746 -856
rect 436982 -1092 437066 -856
rect 437302 -1092 437334 -856
rect 436714 -1176 437334 -1092
rect 436714 -1412 436746 -1176
rect 436982 -1412 437066 -1176
rect 437302 -1412 437334 -1176
rect 436714 -4324 437334 -1412
rect 440434 462052 441054 464004
rect 440434 461816 440466 462052
rect 440702 461816 440786 462052
rect 441022 461816 441054 462052
rect 440434 461732 441054 461816
rect 440434 461496 440466 461732
rect 440702 461496 440786 461732
rect 441022 461496 441054 461732
rect 440434 441174 441054 461496
rect 440434 440938 440466 441174
rect 440702 440938 440786 441174
rect 441022 440938 441054 441174
rect 440434 440854 441054 440938
rect 440434 440618 440466 440854
rect 440702 440618 440786 440854
rect 441022 440618 441054 440854
rect 440434 423174 441054 440618
rect 440434 422938 440466 423174
rect 440702 422938 440786 423174
rect 441022 422938 441054 423174
rect 440434 422854 441054 422938
rect 440434 422618 440466 422854
rect 440702 422618 440786 422854
rect 441022 422618 441054 422854
rect 440434 405174 441054 422618
rect 440434 404938 440466 405174
rect 440702 404938 440786 405174
rect 441022 404938 441054 405174
rect 440434 404854 441054 404938
rect 440434 404618 440466 404854
rect 440702 404618 440786 404854
rect 441022 404618 441054 404854
rect 440434 387174 441054 404618
rect 440434 386938 440466 387174
rect 440702 386938 440786 387174
rect 441022 386938 441054 387174
rect 440434 386854 441054 386938
rect 440434 386618 440466 386854
rect 440702 386618 440786 386854
rect 441022 386618 441054 386854
rect 440434 369174 441054 386618
rect 440434 368938 440466 369174
rect 440702 368938 440786 369174
rect 441022 368938 441054 369174
rect 440434 368854 441054 368938
rect 440434 368618 440466 368854
rect 440702 368618 440786 368854
rect 441022 368618 441054 368854
rect 440434 351174 441054 368618
rect 440434 350938 440466 351174
rect 440702 350938 440786 351174
rect 441022 350938 441054 351174
rect 440434 350854 441054 350938
rect 440434 350618 440466 350854
rect 440702 350618 440786 350854
rect 441022 350618 441054 350854
rect 440434 333174 441054 350618
rect 440434 332938 440466 333174
rect 440702 332938 440786 333174
rect 441022 332938 441054 333174
rect 440434 332854 441054 332938
rect 440434 332618 440466 332854
rect 440702 332618 440786 332854
rect 441022 332618 441054 332854
rect 440434 315174 441054 332618
rect 440434 314938 440466 315174
rect 440702 314938 440786 315174
rect 441022 314938 441054 315174
rect 440434 314854 441054 314938
rect 440434 314618 440466 314854
rect 440702 314618 440786 314854
rect 441022 314618 441054 314854
rect 440434 297174 441054 314618
rect 440434 296938 440466 297174
rect 440702 296938 440786 297174
rect 441022 296938 441054 297174
rect 440434 296854 441054 296938
rect 440434 296618 440466 296854
rect 440702 296618 440786 296854
rect 441022 296618 441054 296854
rect 440434 279174 441054 296618
rect 440434 278938 440466 279174
rect 440702 278938 440786 279174
rect 441022 278938 441054 279174
rect 440434 278854 441054 278938
rect 440434 278618 440466 278854
rect 440702 278618 440786 278854
rect 441022 278618 441054 278854
rect 440434 261174 441054 278618
rect 440434 260938 440466 261174
rect 440702 260938 440786 261174
rect 441022 260938 441054 261174
rect 440434 260854 441054 260938
rect 440434 260618 440466 260854
rect 440702 260618 440786 260854
rect 441022 260618 441054 260854
rect 440434 243174 441054 260618
rect 440434 242938 440466 243174
rect 440702 242938 440786 243174
rect 441022 242938 441054 243174
rect 440434 242854 441054 242938
rect 440434 242618 440466 242854
rect 440702 242618 440786 242854
rect 441022 242618 441054 242854
rect 440434 225174 441054 242618
rect 440434 224938 440466 225174
rect 440702 224938 440786 225174
rect 441022 224938 441054 225174
rect 440434 224854 441054 224938
rect 440434 224618 440466 224854
rect 440702 224618 440786 224854
rect 441022 224618 441054 224854
rect 440434 207174 441054 224618
rect 440434 206938 440466 207174
rect 440702 206938 440786 207174
rect 441022 206938 441054 207174
rect 440434 206854 441054 206938
rect 440434 206618 440466 206854
rect 440702 206618 440786 206854
rect 441022 206618 441054 206854
rect 440434 189174 441054 206618
rect 440434 188938 440466 189174
rect 440702 188938 440786 189174
rect 441022 188938 441054 189174
rect 440434 188854 441054 188938
rect 440434 188618 440466 188854
rect 440702 188618 440786 188854
rect 441022 188618 441054 188854
rect 440434 171174 441054 188618
rect 440434 170938 440466 171174
rect 440702 170938 440786 171174
rect 441022 170938 441054 171174
rect 440434 170854 441054 170938
rect 440434 170618 440466 170854
rect 440702 170618 440786 170854
rect 441022 170618 441054 170854
rect 440434 153174 441054 170618
rect 440434 152938 440466 153174
rect 440702 152938 440786 153174
rect 441022 152938 441054 153174
rect 440434 152854 441054 152938
rect 440434 152618 440466 152854
rect 440702 152618 440786 152854
rect 441022 152618 441054 152854
rect 440434 135174 441054 152618
rect 440434 134938 440466 135174
rect 440702 134938 440786 135174
rect 441022 134938 441054 135174
rect 440434 134854 441054 134938
rect 440434 134618 440466 134854
rect 440702 134618 440786 134854
rect 441022 134618 441054 134854
rect 440434 117174 441054 134618
rect 440434 116938 440466 117174
rect 440702 116938 440786 117174
rect 441022 116938 441054 117174
rect 440434 116854 441054 116938
rect 440434 116618 440466 116854
rect 440702 116618 440786 116854
rect 441022 116618 441054 116854
rect 440434 99174 441054 116618
rect 440434 98938 440466 99174
rect 440702 98938 440786 99174
rect 441022 98938 441054 99174
rect 440434 98854 441054 98938
rect 440434 98618 440466 98854
rect 440702 98618 440786 98854
rect 441022 98618 441054 98854
rect 440434 81174 441054 98618
rect 440434 80938 440466 81174
rect 440702 80938 440786 81174
rect 441022 80938 441054 81174
rect 440434 80854 441054 80938
rect 440434 80618 440466 80854
rect 440702 80618 440786 80854
rect 441022 80618 441054 80854
rect 440434 63174 441054 80618
rect 440434 62938 440466 63174
rect 440702 62938 440786 63174
rect 441022 62938 441054 63174
rect 440434 62854 441054 62938
rect 440434 62618 440466 62854
rect 440702 62618 440786 62854
rect 441022 62618 441054 62854
rect 440434 45174 441054 62618
rect 440434 44938 440466 45174
rect 440702 44938 440786 45174
rect 441022 44938 441054 45174
rect 440434 44854 441054 44938
rect 440434 44618 440466 44854
rect 440702 44618 440786 44854
rect 441022 44618 441054 44854
rect 440434 27174 441054 44618
rect 440434 26938 440466 27174
rect 440702 26938 440786 27174
rect 441022 26938 441054 27174
rect 440434 26854 441054 26938
rect 440434 26618 440466 26854
rect 440702 26618 440786 26854
rect 441022 26618 441054 26854
rect 440434 9174 441054 26618
rect 440434 8938 440466 9174
rect 440702 8938 440786 9174
rect 441022 8938 441054 9174
rect 440434 8854 441054 8938
rect 440434 8618 440466 8854
rect 440702 8618 440786 8854
rect 441022 8618 441054 8854
rect 440434 -1816 441054 8618
rect 440434 -2052 440466 -1816
rect 440702 -2052 440786 -1816
rect 441022 -2052 441054 -1816
rect 440434 -2136 441054 -2052
rect 440434 -2372 440466 -2136
rect 440702 -2372 440786 -2136
rect 441022 -2372 441054 -2136
rect 440434 -4324 441054 -2372
rect 444154 463012 444774 464004
rect 444154 462776 444186 463012
rect 444422 462776 444506 463012
rect 444742 462776 444774 463012
rect 444154 462692 444774 462776
rect 444154 462456 444186 462692
rect 444422 462456 444506 462692
rect 444742 462456 444774 462692
rect 444154 444894 444774 462456
rect 444154 444658 444186 444894
rect 444422 444658 444506 444894
rect 444742 444658 444774 444894
rect 444154 444574 444774 444658
rect 444154 444338 444186 444574
rect 444422 444338 444506 444574
rect 444742 444338 444774 444574
rect 444154 426894 444774 444338
rect 444154 426658 444186 426894
rect 444422 426658 444506 426894
rect 444742 426658 444774 426894
rect 444154 426574 444774 426658
rect 444154 426338 444186 426574
rect 444422 426338 444506 426574
rect 444742 426338 444774 426574
rect 444154 408894 444774 426338
rect 444154 408658 444186 408894
rect 444422 408658 444506 408894
rect 444742 408658 444774 408894
rect 444154 408574 444774 408658
rect 444154 408338 444186 408574
rect 444422 408338 444506 408574
rect 444742 408338 444774 408574
rect 444154 390894 444774 408338
rect 444154 390658 444186 390894
rect 444422 390658 444506 390894
rect 444742 390658 444774 390894
rect 444154 390574 444774 390658
rect 444154 390338 444186 390574
rect 444422 390338 444506 390574
rect 444742 390338 444774 390574
rect 444154 372894 444774 390338
rect 444154 372658 444186 372894
rect 444422 372658 444506 372894
rect 444742 372658 444774 372894
rect 444154 372574 444774 372658
rect 444154 372338 444186 372574
rect 444422 372338 444506 372574
rect 444742 372338 444774 372574
rect 444154 354894 444774 372338
rect 444154 354658 444186 354894
rect 444422 354658 444506 354894
rect 444742 354658 444774 354894
rect 444154 354574 444774 354658
rect 444154 354338 444186 354574
rect 444422 354338 444506 354574
rect 444742 354338 444774 354574
rect 444154 336894 444774 354338
rect 444154 336658 444186 336894
rect 444422 336658 444506 336894
rect 444742 336658 444774 336894
rect 444154 336574 444774 336658
rect 444154 336338 444186 336574
rect 444422 336338 444506 336574
rect 444742 336338 444774 336574
rect 444154 318894 444774 336338
rect 444154 318658 444186 318894
rect 444422 318658 444506 318894
rect 444742 318658 444774 318894
rect 444154 318574 444774 318658
rect 444154 318338 444186 318574
rect 444422 318338 444506 318574
rect 444742 318338 444774 318574
rect 444154 300894 444774 318338
rect 444154 300658 444186 300894
rect 444422 300658 444506 300894
rect 444742 300658 444774 300894
rect 444154 300574 444774 300658
rect 444154 300338 444186 300574
rect 444422 300338 444506 300574
rect 444742 300338 444774 300574
rect 444154 282894 444774 300338
rect 444154 282658 444186 282894
rect 444422 282658 444506 282894
rect 444742 282658 444774 282894
rect 444154 282574 444774 282658
rect 444154 282338 444186 282574
rect 444422 282338 444506 282574
rect 444742 282338 444774 282574
rect 444154 264894 444774 282338
rect 444154 264658 444186 264894
rect 444422 264658 444506 264894
rect 444742 264658 444774 264894
rect 444154 264574 444774 264658
rect 444154 264338 444186 264574
rect 444422 264338 444506 264574
rect 444742 264338 444774 264574
rect 444154 246894 444774 264338
rect 444154 246658 444186 246894
rect 444422 246658 444506 246894
rect 444742 246658 444774 246894
rect 444154 246574 444774 246658
rect 444154 246338 444186 246574
rect 444422 246338 444506 246574
rect 444742 246338 444774 246574
rect 444154 228894 444774 246338
rect 444154 228658 444186 228894
rect 444422 228658 444506 228894
rect 444742 228658 444774 228894
rect 444154 228574 444774 228658
rect 444154 228338 444186 228574
rect 444422 228338 444506 228574
rect 444742 228338 444774 228574
rect 444154 210894 444774 228338
rect 444154 210658 444186 210894
rect 444422 210658 444506 210894
rect 444742 210658 444774 210894
rect 444154 210574 444774 210658
rect 444154 210338 444186 210574
rect 444422 210338 444506 210574
rect 444742 210338 444774 210574
rect 444154 192894 444774 210338
rect 444154 192658 444186 192894
rect 444422 192658 444506 192894
rect 444742 192658 444774 192894
rect 444154 192574 444774 192658
rect 444154 192338 444186 192574
rect 444422 192338 444506 192574
rect 444742 192338 444774 192574
rect 444154 174894 444774 192338
rect 444154 174658 444186 174894
rect 444422 174658 444506 174894
rect 444742 174658 444774 174894
rect 444154 174574 444774 174658
rect 444154 174338 444186 174574
rect 444422 174338 444506 174574
rect 444742 174338 444774 174574
rect 444154 156894 444774 174338
rect 444154 156658 444186 156894
rect 444422 156658 444506 156894
rect 444742 156658 444774 156894
rect 444154 156574 444774 156658
rect 444154 156338 444186 156574
rect 444422 156338 444506 156574
rect 444742 156338 444774 156574
rect 444154 138894 444774 156338
rect 444154 138658 444186 138894
rect 444422 138658 444506 138894
rect 444742 138658 444774 138894
rect 444154 138574 444774 138658
rect 444154 138338 444186 138574
rect 444422 138338 444506 138574
rect 444742 138338 444774 138574
rect 444154 120894 444774 138338
rect 444154 120658 444186 120894
rect 444422 120658 444506 120894
rect 444742 120658 444774 120894
rect 444154 120574 444774 120658
rect 444154 120338 444186 120574
rect 444422 120338 444506 120574
rect 444742 120338 444774 120574
rect 444154 102894 444774 120338
rect 444154 102658 444186 102894
rect 444422 102658 444506 102894
rect 444742 102658 444774 102894
rect 444154 102574 444774 102658
rect 444154 102338 444186 102574
rect 444422 102338 444506 102574
rect 444742 102338 444774 102574
rect 444154 84894 444774 102338
rect 444154 84658 444186 84894
rect 444422 84658 444506 84894
rect 444742 84658 444774 84894
rect 444154 84574 444774 84658
rect 444154 84338 444186 84574
rect 444422 84338 444506 84574
rect 444742 84338 444774 84574
rect 444154 66894 444774 84338
rect 444154 66658 444186 66894
rect 444422 66658 444506 66894
rect 444742 66658 444774 66894
rect 444154 66574 444774 66658
rect 444154 66338 444186 66574
rect 444422 66338 444506 66574
rect 444742 66338 444774 66574
rect 444154 48894 444774 66338
rect 444154 48658 444186 48894
rect 444422 48658 444506 48894
rect 444742 48658 444774 48894
rect 444154 48574 444774 48658
rect 444154 48338 444186 48574
rect 444422 48338 444506 48574
rect 444742 48338 444774 48574
rect 444154 30894 444774 48338
rect 444154 30658 444186 30894
rect 444422 30658 444506 30894
rect 444742 30658 444774 30894
rect 444154 30574 444774 30658
rect 444154 30338 444186 30574
rect 444422 30338 444506 30574
rect 444742 30338 444774 30574
rect 444154 12894 444774 30338
rect 444154 12658 444186 12894
rect 444422 12658 444506 12894
rect 444742 12658 444774 12894
rect 444154 12574 444774 12658
rect 444154 12338 444186 12574
rect 444422 12338 444506 12574
rect 444742 12338 444774 12574
rect 444154 -2776 444774 12338
rect 444154 -3012 444186 -2776
rect 444422 -3012 444506 -2776
rect 444742 -3012 444774 -2776
rect 444154 -3096 444774 -3012
rect 444154 -3332 444186 -3096
rect 444422 -3332 444506 -3096
rect 444742 -3332 444774 -3096
rect 444154 -4324 444774 -3332
rect 447874 463972 448494 464004
rect 447874 463736 447906 463972
rect 448142 463736 448226 463972
rect 448462 463736 448494 463972
rect 447874 463652 448494 463736
rect 447874 463416 447906 463652
rect 448142 463416 448226 463652
rect 448462 463416 448494 463652
rect 447874 448614 448494 463416
rect 447874 448378 447906 448614
rect 448142 448378 448226 448614
rect 448462 448378 448494 448614
rect 447874 448294 448494 448378
rect 447874 448058 447906 448294
rect 448142 448058 448226 448294
rect 448462 448058 448494 448294
rect 447874 430614 448494 448058
rect 447874 430378 447906 430614
rect 448142 430378 448226 430614
rect 448462 430378 448494 430614
rect 447874 430294 448494 430378
rect 447874 430058 447906 430294
rect 448142 430058 448226 430294
rect 448462 430058 448494 430294
rect 447874 412614 448494 430058
rect 447874 412378 447906 412614
rect 448142 412378 448226 412614
rect 448462 412378 448494 412614
rect 447874 412294 448494 412378
rect 447874 412058 447906 412294
rect 448142 412058 448226 412294
rect 448462 412058 448494 412294
rect 447874 394614 448494 412058
rect 447874 394378 447906 394614
rect 448142 394378 448226 394614
rect 448462 394378 448494 394614
rect 447874 394294 448494 394378
rect 447874 394058 447906 394294
rect 448142 394058 448226 394294
rect 448462 394058 448494 394294
rect 447874 376614 448494 394058
rect 447874 376378 447906 376614
rect 448142 376378 448226 376614
rect 448462 376378 448494 376614
rect 447874 376294 448494 376378
rect 447874 376058 447906 376294
rect 448142 376058 448226 376294
rect 448462 376058 448494 376294
rect 447874 358614 448494 376058
rect 447874 358378 447906 358614
rect 448142 358378 448226 358614
rect 448462 358378 448494 358614
rect 447874 358294 448494 358378
rect 447874 358058 447906 358294
rect 448142 358058 448226 358294
rect 448462 358058 448494 358294
rect 447874 340614 448494 358058
rect 447874 340378 447906 340614
rect 448142 340378 448226 340614
rect 448462 340378 448494 340614
rect 447874 340294 448494 340378
rect 447874 340058 447906 340294
rect 448142 340058 448226 340294
rect 448462 340058 448494 340294
rect 447874 322614 448494 340058
rect 447874 322378 447906 322614
rect 448142 322378 448226 322614
rect 448462 322378 448494 322614
rect 447874 322294 448494 322378
rect 447874 322058 447906 322294
rect 448142 322058 448226 322294
rect 448462 322058 448494 322294
rect 447874 304614 448494 322058
rect 447874 304378 447906 304614
rect 448142 304378 448226 304614
rect 448462 304378 448494 304614
rect 447874 304294 448494 304378
rect 447874 304058 447906 304294
rect 448142 304058 448226 304294
rect 448462 304058 448494 304294
rect 447874 286614 448494 304058
rect 447874 286378 447906 286614
rect 448142 286378 448226 286614
rect 448462 286378 448494 286614
rect 447874 286294 448494 286378
rect 447874 286058 447906 286294
rect 448142 286058 448226 286294
rect 448462 286058 448494 286294
rect 447874 268614 448494 286058
rect 447874 268378 447906 268614
rect 448142 268378 448226 268614
rect 448462 268378 448494 268614
rect 447874 268294 448494 268378
rect 447874 268058 447906 268294
rect 448142 268058 448226 268294
rect 448462 268058 448494 268294
rect 447874 250614 448494 268058
rect 447874 250378 447906 250614
rect 448142 250378 448226 250614
rect 448462 250378 448494 250614
rect 447874 250294 448494 250378
rect 447874 250058 447906 250294
rect 448142 250058 448226 250294
rect 448462 250058 448494 250294
rect 447874 232614 448494 250058
rect 447874 232378 447906 232614
rect 448142 232378 448226 232614
rect 448462 232378 448494 232614
rect 447874 232294 448494 232378
rect 447874 232058 447906 232294
rect 448142 232058 448226 232294
rect 448462 232058 448494 232294
rect 447874 214614 448494 232058
rect 447874 214378 447906 214614
rect 448142 214378 448226 214614
rect 448462 214378 448494 214614
rect 447874 214294 448494 214378
rect 447874 214058 447906 214294
rect 448142 214058 448226 214294
rect 448462 214058 448494 214294
rect 447874 196614 448494 214058
rect 447874 196378 447906 196614
rect 448142 196378 448226 196614
rect 448462 196378 448494 196614
rect 447874 196294 448494 196378
rect 447874 196058 447906 196294
rect 448142 196058 448226 196294
rect 448462 196058 448494 196294
rect 447874 178614 448494 196058
rect 447874 178378 447906 178614
rect 448142 178378 448226 178614
rect 448462 178378 448494 178614
rect 447874 178294 448494 178378
rect 447874 178058 447906 178294
rect 448142 178058 448226 178294
rect 448462 178058 448494 178294
rect 447874 160614 448494 178058
rect 447874 160378 447906 160614
rect 448142 160378 448226 160614
rect 448462 160378 448494 160614
rect 447874 160294 448494 160378
rect 447874 160058 447906 160294
rect 448142 160058 448226 160294
rect 448462 160058 448494 160294
rect 447874 142614 448494 160058
rect 447874 142378 447906 142614
rect 448142 142378 448226 142614
rect 448462 142378 448494 142614
rect 447874 142294 448494 142378
rect 447874 142058 447906 142294
rect 448142 142058 448226 142294
rect 448462 142058 448494 142294
rect 447874 124614 448494 142058
rect 447874 124378 447906 124614
rect 448142 124378 448226 124614
rect 448462 124378 448494 124614
rect 447874 124294 448494 124378
rect 447874 124058 447906 124294
rect 448142 124058 448226 124294
rect 448462 124058 448494 124294
rect 447874 106614 448494 124058
rect 447874 106378 447906 106614
rect 448142 106378 448226 106614
rect 448462 106378 448494 106614
rect 447874 106294 448494 106378
rect 447874 106058 447906 106294
rect 448142 106058 448226 106294
rect 448462 106058 448494 106294
rect 447874 88614 448494 106058
rect 447874 88378 447906 88614
rect 448142 88378 448226 88614
rect 448462 88378 448494 88614
rect 447874 88294 448494 88378
rect 447874 88058 447906 88294
rect 448142 88058 448226 88294
rect 448462 88058 448494 88294
rect 447874 70614 448494 88058
rect 447874 70378 447906 70614
rect 448142 70378 448226 70614
rect 448462 70378 448494 70614
rect 447874 70294 448494 70378
rect 447874 70058 447906 70294
rect 448142 70058 448226 70294
rect 448462 70058 448494 70294
rect 447874 52614 448494 70058
rect 447874 52378 447906 52614
rect 448142 52378 448226 52614
rect 448462 52378 448494 52614
rect 447874 52294 448494 52378
rect 447874 52058 447906 52294
rect 448142 52058 448226 52294
rect 448462 52058 448494 52294
rect 447874 34614 448494 52058
rect 447874 34378 447906 34614
rect 448142 34378 448226 34614
rect 448462 34378 448494 34614
rect 447874 34294 448494 34378
rect 447874 34058 447906 34294
rect 448142 34058 448226 34294
rect 448462 34058 448494 34294
rect 447874 16614 448494 34058
rect 447874 16378 447906 16614
rect 448142 16378 448226 16614
rect 448462 16378 448494 16614
rect 447874 16294 448494 16378
rect 447874 16058 447906 16294
rect 448142 16058 448226 16294
rect 448462 16058 448494 16294
rect 447874 -3736 448494 16058
rect 447874 -3972 447906 -3736
rect 448142 -3972 448226 -3736
rect 448462 -3972 448494 -3736
rect 447874 -4056 448494 -3972
rect 447874 -4292 447906 -4056
rect 448142 -4292 448226 -4056
rect 448462 -4292 448494 -4056
rect 447874 -4324 448494 -4292
rect 454714 461092 455334 464004
rect 454714 460856 454746 461092
rect 454982 460856 455066 461092
rect 455302 460856 455334 461092
rect 454714 460772 455334 460856
rect 454714 460536 454746 460772
rect 454982 460536 455066 460772
rect 455302 460536 455334 460772
rect 454714 455454 455334 460536
rect 454714 455218 454746 455454
rect 454982 455218 455066 455454
rect 455302 455218 455334 455454
rect 454714 455134 455334 455218
rect 454714 454898 454746 455134
rect 454982 454898 455066 455134
rect 455302 454898 455334 455134
rect 454714 437454 455334 454898
rect 454714 437218 454746 437454
rect 454982 437218 455066 437454
rect 455302 437218 455334 437454
rect 454714 437134 455334 437218
rect 454714 436898 454746 437134
rect 454982 436898 455066 437134
rect 455302 436898 455334 437134
rect 454714 419454 455334 436898
rect 454714 419218 454746 419454
rect 454982 419218 455066 419454
rect 455302 419218 455334 419454
rect 454714 419134 455334 419218
rect 454714 418898 454746 419134
rect 454982 418898 455066 419134
rect 455302 418898 455334 419134
rect 454714 401454 455334 418898
rect 454714 401218 454746 401454
rect 454982 401218 455066 401454
rect 455302 401218 455334 401454
rect 454714 401134 455334 401218
rect 454714 400898 454746 401134
rect 454982 400898 455066 401134
rect 455302 400898 455334 401134
rect 454714 383454 455334 400898
rect 454714 383218 454746 383454
rect 454982 383218 455066 383454
rect 455302 383218 455334 383454
rect 454714 383134 455334 383218
rect 454714 382898 454746 383134
rect 454982 382898 455066 383134
rect 455302 382898 455334 383134
rect 454714 365454 455334 382898
rect 454714 365218 454746 365454
rect 454982 365218 455066 365454
rect 455302 365218 455334 365454
rect 454714 365134 455334 365218
rect 454714 364898 454746 365134
rect 454982 364898 455066 365134
rect 455302 364898 455334 365134
rect 454714 347454 455334 364898
rect 454714 347218 454746 347454
rect 454982 347218 455066 347454
rect 455302 347218 455334 347454
rect 454714 347134 455334 347218
rect 454714 346898 454746 347134
rect 454982 346898 455066 347134
rect 455302 346898 455334 347134
rect 454714 329454 455334 346898
rect 454714 329218 454746 329454
rect 454982 329218 455066 329454
rect 455302 329218 455334 329454
rect 454714 329134 455334 329218
rect 454714 328898 454746 329134
rect 454982 328898 455066 329134
rect 455302 328898 455334 329134
rect 454714 311454 455334 328898
rect 454714 311218 454746 311454
rect 454982 311218 455066 311454
rect 455302 311218 455334 311454
rect 454714 311134 455334 311218
rect 454714 310898 454746 311134
rect 454982 310898 455066 311134
rect 455302 310898 455334 311134
rect 454714 293454 455334 310898
rect 454714 293218 454746 293454
rect 454982 293218 455066 293454
rect 455302 293218 455334 293454
rect 454714 293134 455334 293218
rect 454714 292898 454746 293134
rect 454982 292898 455066 293134
rect 455302 292898 455334 293134
rect 454714 275454 455334 292898
rect 454714 275218 454746 275454
rect 454982 275218 455066 275454
rect 455302 275218 455334 275454
rect 454714 275134 455334 275218
rect 454714 274898 454746 275134
rect 454982 274898 455066 275134
rect 455302 274898 455334 275134
rect 454714 257454 455334 274898
rect 454714 257218 454746 257454
rect 454982 257218 455066 257454
rect 455302 257218 455334 257454
rect 454714 257134 455334 257218
rect 454714 256898 454746 257134
rect 454982 256898 455066 257134
rect 455302 256898 455334 257134
rect 454714 239454 455334 256898
rect 454714 239218 454746 239454
rect 454982 239218 455066 239454
rect 455302 239218 455334 239454
rect 454714 239134 455334 239218
rect 454714 238898 454746 239134
rect 454982 238898 455066 239134
rect 455302 238898 455334 239134
rect 454714 221454 455334 238898
rect 454714 221218 454746 221454
rect 454982 221218 455066 221454
rect 455302 221218 455334 221454
rect 454714 221134 455334 221218
rect 454714 220898 454746 221134
rect 454982 220898 455066 221134
rect 455302 220898 455334 221134
rect 454714 203454 455334 220898
rect 454714 203218 454746 203454
rect 454982 203218 455066 203454
rect 455302 203218 455334 203454
rect 454714 203134 455334 203218
rect 454714 202898 454746 203134
rect 454982 202898 455066 203134
rect 455302 202898 455334 203134
rect 454714 185454 455334 202898
rect 454714 185218 454746 185454
rect 454982 185218 455066 185454
rect 455302 185218 455334 185454
rect 454714 185134 455334 185218
rect 454714 184898 454746 185134
rect 454982 184898 455066 185134
rect 455302 184898 455334 185134
rect 454714 167454 455334 184898
rect 454714 167218 454746 167454
rect 454982 167218 455066 167454
rect 455302 167218 455334 167454
rect 454714 167134 455334 167218
rect 454714 166898 454746 167134
rect 454982 166898 455066 167134
rect 455302 166898 455334 167134
rect 454714 149454 455334 166898
rect 454714 149218 454746 149454
rect 454982 149218 455066 149454
rect 455302 149218 455334 149454
rect 454714 149134 455334 149218
rect 454714 148898 454746 149134
rect 454982 148898 455066 149134
rect 455302 148898 455334 149134
rect 454714 131454 455334 148898
rect 454714 131218 454746 131454
rect 454982 131218 455066 131454
rect 455302 131218 455334 131454
rect 454714 131134 455334 131218
rect 454714 130898 454746 131134
rect 454982 130898 455066 131134
rect 455302 130898 455334 131134
rect 454714 113454 455334 130898
rect 454714 113218 454746 113454
rect 454982 113218 455066 113454
rect 455302 113218 455334 113454
rect 454714 113134 455334 113218
rect 454714 112898 454746 113134
rect 454982 112898 455066 113134
rect 455302 112898 455334 113134
rect 454714 95454 455334 112898
rect 454714 95218 454746 95454
rect 454982 95218 455066 95454
rect 455302 95218 455334 95454
rect 454714 95134 455334 95218
rect 454714 94898 454746 95134
rect 454982 94898 455066 95134
rect 455302 94898 455334 95134
rect 454714 77454 455334 94898
rect 454714 77218 454746 77454
rect 454982 77218 455066 77454
rect 455302 77218 455334 77454
rect 454714 77134 455334 77218
rect 454714 76898 454746 77134
rect 454982 76898 455066 77134
rect 455302 76898 455334 77134
rect 454714 59454 455334 76898
rect 454714 59218 454746 59454
rect 454982 59218 455066 59454
rect 455302 59218 455334 59454
rect 454714 59134 455334 59218
rect 454714 58898 454746 59134
rect 454982 58898 455066 59134
rect 455302 58898 455334 59134
rect 454714 41454 455334 58898
rect 454714 41218 454746 41454
rect 454982 41218 455066 41454
rect 455302 41218 455334 41454
rect 454714 41134 455334 41218
rect 454714 40898 454746 41134
rect 454982 40898 455066 41134
rect 455302 40898 455334 41134
rect 454714 23454 455334 40898
rect 454714 23218 454746 23454
rect 454982 23218 455066 23454
rect 455302 23218 455334 23454
rect 454714 23134 455334 23218
rect 454714 22898 454746 23134
rect 454982 22898 455066 23134
rect 455302 22898 455334 23134
rect 454714 5454 455334 22898
rect 454714 5218 454746 5454
rect 454982 5218 455066 5454
rect 455302 5218 455334 5454
rect 454714 5134 455334 5218
rect 454714 4898 454746 5134
rect 454982 4898 455066 5134
rect 455302 4898 455334 5134
rect 454714 -856 455334 4898
rect 454714 -1092 454746 -856
rect 454982 -1092 455066 -856
rect 455302 -1092 455334 -856
rect 454714 -1176 455334 -1092
rect 454714 -1412 454746 -1176
rect 454982 -1412 455066 -1176
rect 455302 -1412 455334 -1176
rect 454714 -4324 455334 -1412
rect 458434 462052 459054 464004
rect 458434 461816 458466 462052
rect 458702 461816 458786 462052
rect 459022 461816 459054 462052
rect 458434 461732 459054 461816
rect 458434 461496 458466 461732
rect 458702 461496 458786 461732
rect 459022 461496 459054 461732
rect 458434 441174 459054 461496
rect 458434 440938 458466 441174
rect 458702 440938 458786 441174
rect 459022 440938 459054 441174
rect 458434 440854 459054 440938
rect 458434 440618 458466 440854
rect 458702 440618 458786 440854
rect 459022 440618 459054 440854
rect 458434 423174 459054 440618
rect 458434 422938 458466 423174
rect 458702 422938 458786 423174
rect 459022 422938 459054 423174
rect 458434 422854 459054 422938
rect 458434 422618 458466 422854
rect 458702 422618 458786 422854
rect 459022 422618 459054 422854
rect 458434 405174 459054 422618
rect 458434 404938 458466 405174
rect 458702 404938 458786 405174
rect 459022 404938 459054 405174
rect 458434 404854 459054 404938
rect 458434 404618 458466 404854
rect 458702 404618 458786 404854
rect 459022 404618 459054 404854
rect 458434 387174 459054 404618
rect 458434 386938 458466 387174
rect 458702 386938 458786 387174
rect 459022 386938 459054 387174
rect 458434 386854 459054 386938
rect 458434 386618 458466 386854
rect 458702 386618 458786 386854
rect 459022 386618 459054 386854
rect 458434 369174 459054 386618
rect 458434 368938 458466 369174
rect 458702 368938 458786 369174
rect 459022 368938 459054 369174
rect 458434 368854 459054 368938
rect 458434 368618 458466 368854
rect 458702 368618 458786 368854
rect 459022 368618 459054 368854
rect 458434 351174 459054 368618
rect 458434 350938 458466 351174
rect 458702 350938 458786 351174
rect 459022 350938 459054 351174
rect 458434 350854 459054 350938
rect 458434 350618 458466 350854
rect 458702 350618 458786 350854
rect 459022 350618 459054 350854
rect 458434 333174 459054 350618
rect 458434 332938 458466 333174
rect 458702 332938 458786 333174
rect 459022 332938 459054 333174
rect 458434 332854 459054 332938
rect 458434 332618 458466 332854
rect 458702 332618 458786 332854
rect 459022 332618 459054 332854
rect 458434 315174 459054 332618
rect 458434 314938 458466 315174
rect 458702 314938 458786 315174
rect 459022 314938 459054 315174
rect 458434 314854 459054 314938
rect 458434 314618 458466 314854
rect 458702 314618 458786 314854
rect 459022 314618 459054 314854
rect 458434 297174 459054 314618
rect 458434 296938 458466 297174
rect 458702 296938 458786 297174
rect 459022 296938 459054 297174
rect 458434 296854 459054 296938
rect 458434 296618 458466 296854
rect 458702 296618 458786 296854
rect 459022 296618 459054 296854
rect 458434 279174 459054 296618
rect 458434 278938 458466 279174
rect 458702 278938 458786 279174
rect 459022 278938 459054 279174
rect 458434 278854 459054 278938
rect 458434 278618 458466 278854
rect 458702 278618 458786 278854
rect 459022 278618 459054 278854
rect 458434 261174 459054 278618
rect 458434 260938 458466 261174
rect 458702 260938 458786 261174
rect 459022 260938 459054 261174
rect 458434 260854 459054 260938
rect 458434 260618 458466 260854
rect 458702 260618 458786 260854
rect 459022 260618 459054 260854
rect 458434 243174 459054 260618
rect 458434 242938 458466 243174
rect 458702 242938 458786 243174
rect 459022 242938 459054 243174
rect 458434 242854 459054 242938
rect 458434 242618 458466 242854
rect 458702 242618 458786 242854
rect 459022 242618 459054 242854
rect 458434 225174 459054 242618
rect 458434 224938 458466 225174
rect 458702 224938 458786 225174
rect 459022 224938 459054 225174
rect 458434 224854 459054 224938
rect 458434 224618 458466 224854
rect 458702 224618 458786 224854
rect 459022 224618 459054 224854
rect 458434 207174 459054 224618
rect 458434 206938 458466 207174
rect 458702 206938 458786 207174
rect 459022 206938 459054 207174
rect 458434 206854 459054 206938
rect 458434 206618 458466 206854
rect 458702 206618 458786 206854
rect 459022 206618 459054 206854
rect 458434 189174 459054 206618
rect 458434 188938 458466 189174
rect 458702 188938 458786 189174
rect 459022 188938 459054 189174
rect 458434 188854 459054 188938
rect 458434 188618 458466 188854
rect 458702 188618 458786 188854
rect 459022 188618 459054 188854
rect 458434 171174 459054 188618
rect 458434 170938 458466 171174
rect 458702 170938 458786 171174
rect 459022 170938 459054 171174
rect 458434 170854 459054 170938
rect 458434 170618 458466 170854
rect 458702 170618 458786 170854
rect 459022 170618 459054 170854
rect 458434 153174 459054 170618
rect 458434 152938 458466 153174
rect 458702 152938 458786 153174
rect 459022 152938 459054 153174
rect 458434 152854 459054 152938
rect 458434 152618 458466 152854
rect 458702 152618 458786 152854
rect 459022 152618 459054 152854
rect 458434 135174 459054 152618
rect 458434 134938 458466 135174
rect 458702 134938 458786 135174
rect 459022 134938 459054 135174
rect 458434 134854 459054 134938
rect 458434 134618 458466 134854
rect 458702 134618 458786 134854
rect 459022 134618 459054 134854
rect 458434 117174 459054 134618
rect 458434 116938 458466 117174
rect 458702 116938 458786 117174
rect 459022 116938 459054 117174
rect 458434 116854 459054 116938
rect 458434 116618 458466 116854
rect 458702 116618 458786 116854
rect 459022 116618 459054 116854
rect 458434 99174 459054 116618
rect 458434 98938 458466 99174
rect 458702 98938 458786 99174
rect 459022 98938 459054 99174
rect 458434 98854 459054 98938
rect 458434 98618 458466 98854
rect 458702 98618 458786 98854
rect 459022 98618 459054 98854
rect 458434 81174 459054 98618
rect 458434 80938 458466 81174
rect 458702 80938 458786 81174
rect 459022 80938 459054 81174
rect 458434 80854 459054 80938
rect 458434 80618 458466 80854
rect 458702 80618 458786 80854
rect 459022 80618 459054 80854
rect 458434 63174 459054 80618
rect 458434 62938 458466 63174
rect 458702 62938 458786 63174
rect 459022 62938 459054 63174
rect 458434 62854 459054 62938
rect 458434 62618 458466 62854
rect 458702 62618 458786 62854
rect 459022 62618 459054 62854
rect 458434 45174 459054 62618
rect 458434 44938 458466 45174
rect 458702 44938 458786 45174
rect 459022 44938 459054 45174
rect 458434 44854 459054 44938
rect 458434 44618 458466 44854
rect 458702 44618 458786 44854
rect 459022 44618 459054 44854
rect 458434 27174 459054 44618
rect 458434 26938 458466 27174
rect 458702 26938 458786 27174
rect 459022 26938 459054 27174
rect 458434 26854 459054 26938
rect 458434 26618 458466 26854
rect 458702 26618 458786 26854
rect 459022 26618 459054 26854
rect 458434 9174 459054 26618
rect 458434 8938 458466 9174
rect 458702 8938 458786 9174
rect 459022 8938 459054 9174
rect 458434 8854 459054 8938
rect 458434 8618 458466 8854
rect 458702 8618 458786 8854
rect 459022 8618 459054 8854
rect 458434 -1816 459054 8618
rect 458434 -2052 458466 -1816
rect 458702 -2052 458786 -1816
rect 459022 -2052 459054 -1816
rect 458434 -2136 459054 -2052
rect 458434 -2372 458466 -2136
rect 458702 -2372 458786 -2136
rect 459022 -2372 459054 -2136
rect 458434 -4324 459054 -2372
rect 462154 463012 462774 464004
rect 462154 462776 462186 463012
rect 462422 462776 462506 463012
rect 462742 462776 462774 463012
rect 462154 462692 462774 462776
rect 462154 462456 462186 462692
rect 462422 462456 462506 462692
rect 462742 462456 462774 462692
rect 462154 444894 462774 462456
rect 462154 444658 462186 444894
rect 462422 444658 462506 444894
rect 462742 444658 462774 444894
rect 462154 444574 462774 444658
rect 462154 444338 462186 444574
rect 462422 444338 462506 444574
rect 462742 444338 462774 444574
rect 462154 426894 462774 444338
rect 462154 426658 462186 426894
rect 462422 426658 462506 426894
rect 462742 426658 462774 426894
rect 462154 426574 462774 426658
rect 462154 426338 462186 426574
rect 462422 426338 462506 426574
rect 462742 426338 462774 426574
rect 462154 408894 462774 426338
rect 462154 408658 462186 408894
rect 462422 408658 462506 408894
rect 462742 408658 462774 408894
rect 462154 408574 462774 408658
rect 462154 408338 462186 408574
rect 462422 408338 462506 408574
rect 462742 408338 462774 408574
rect 462154 390894 462774 408338
rect 462154 390658 462186 390894
rect 462422 390658 462506 390894
rect 462742 390658 462774 390894
rect 462154 390574 462774 390658
rect 462154 390338 462186 390574
rect 462422 390338 462506 390574
rect 462742 390338 462774 390574
rect 462154 372894 462774 390338
rect 462154 372658 462186 372894
rect 462422 372658 462506 372894
rect 462742 372658 462774 372894
rect 462154 372574 462774 372658
rect 462154 372338 462186 372574
rect 462422 372338 462506 372574
rect 462742 372338 462774 372574
rect 462154 354894 462774 372338
rect 462154 354658 462186 354894
rect 462422 354658 462506 354894
rect 462742 354658 462774 354894
rect 462154 354574 462774 354658
rect 462154 354338 462186 354574
rect 462422 354338 462506 354574
rect 462742 354338 462774 354574
rect 462154 336894 462774 354338
rect 462154 336658 462186 336894
rect 462422 336658 462506 336894
rect 462742 336658 462774 336894
rect 462154 336574 462774 336658
rect 462154 336338 462186 336574
rect 462422 336338 462506 336574
rect 462742 336338 462774 336574
rect 462154 318894 462774 336338
rect 462154 318658 462186 318894
rect 462422 318658 462506 318894
rect 462742 318658 462774 318894
rect 462154 318574 462774 318658
rect 462154 318338 462186 318574
rect 462422 318338 462506 318574
rect 462742 318338 462774 318574
rect 462154 300894 462774 318338
rect 462154 300658 462186 300894
rect 462422 300658 462506 300894
rect 462742 300658 462774 300894
rect 462154 300574 462774 300658
rect 462154 300338 462186 300574
rect 462422 300338 462506 300574
rect 462742 300338 462774 300574
rect 462154 282894 462774 300338
rect 462154 282658 462186 282894
rect 462422 282658 462506 282894
rect 462742 282658 462774 282894
rect 462154 282574 462774 282658
rect 462154 282338 462186 282574
rect 462422 282338 462506 282574
rect 462742 282338 462774 282574
rect 462154 264894 462774 282338
rect 462154 264658 462186 264894
rect 462422 264658 462506 264894
rect 462742 264658 462774 264894
rect 462154 264574 462774 264658
rect 462154 264338 462186 264574
rect 462422 264338 462506 264574
rect 462742 264338 462774 264574
rect 462154 246894 462774 264338
rect 462154 246658 462186 246894
rect 462422 246658 462506 246894
rect 462742 246658 462774 246894
rect 462154 246574 462774 246658
rect 462154 246338 462186 246574
rect 462422 246338 462506 246574
rect 462742 246338 462774 246574
rect 462154 228894 462774 246338
rect 462154 228658 462186 228894
rect 462422 228658 462506 228894
rect 462742 228658 462774 228894
rect 462154 228574 462774 228658
rect 462154 228338 462186 228574
rect 462422 228338 462506 228574
rect 462742 228338 462774 228574
rect 462154 210894 462774 228338
rect 462154 210658 462186 210894
rect 462422 210658 462506 210894
rect 462742 210658 462774 210894
rect 462154 210574 462774 210658
rect 462154 210338 462186 210574
rect 462422 210338 462506 210574
rect 462742 210338 462774 210574
rect 462154 192894 462774 210338
rect 462154 192658 462186 192894
rect 462422 192658 462506 192894
rect 462742 192658 462774 192894
rect 462154 192574 462774 192658
rect 462154 192338 462186 192574
rect 462422 192338 462506 192574
rect 462742 192338 462774 192574
rect 462154 174894 462774 192338
rect 462154 174658 462186 174894
rect 462422 174658 462506 174894
rect 462742 174658 462774 174894
rect 462154 174574 462774 174658
rect 462154 174338 462186 174574
rect 462422 174338 462506 174574
rect 462742 174338 462774 174574
rect 462154 156894 462774 174338
rect 462154 156658 462186 156894
rect 462422 156658 462506 156894
rect 462742 156658 462774 156894
rect 462154 156574 462774 156658
rect 462154 156338 462186 156574
rect 462422 156338 462506 156574
rect 462742 156338 462774 156574
rect 462154 138894 462774 156338
rect 462154 138658 462186 138894
rect 462422 138658 462506 138894
rect 462742 138658 462774 138894
rect 462154 138574 462774 138658
rect 462154 138338 462186 138574
rect 462422 138338 462506 138574
rect 462742 138338 462774 138574
rect 462154 120894 462774 138338
rect 462154 120658 462186 120894
rect 462422 120658 462506 120894
rect 462742 120658 462774 120894
rect 462154 120574 462774 120658
rect 462154 120338 462186 120574
rect 462422 120338 462506 120574
rect 462742 120338 462774 120574
rect 462154 102894 462774 120338
rect 462154 102658 462186 102894
rect 462422 102658 462506 102894
rect 462742 102658 462774 102894
rect 462154 102574 462774 102658
rect 462154 102338 462186 102574
rect 462422 102338 462506 102574
rect 462742 102338 462774 102574
rect 462154 84894 462774 102338
rect 462154 84658 462186 84894
rect 462422 84658 462506 84894
rect 462742 84658 462774 84894
rect 462154 84574 462774 84658
rect 462154 84338 462186 84574
rect 462422 84338 462506 84574
rect 462742 84338 462774 84574
rect 462154 66894 462774 84338
rect 462154 66658 462186 66894
rect 462422 66658 462506 66894
rect 462742 66658 462774 66894
rect 462154 66574 462774 66658
rect 462154 66338 462186 66574
rect 462422 66338 462506 66574
rect 462742 66338 462774 66574
rect 462154 48894 462774 66338
rect 462154 48658 462186 48894
rect 462422 48658 462506 48894
rect 462742 48658 462774 48894
rect 462154 48574 462774 48658
rect 462154 48338 462186 48574
rect 462422 48338 462506 48574
rect 462742 48338 462774 48574
rect 462154 30894 462774 48338
rect 462154 30658 462186 30894
rect 462422 30658 462506 30894
rect 462742 30658 462774 30894
rect 462154 30574 462774 30658
rect 462154 30338 462186 30574
rect 462422 30338 462506 30574
rect 462742 30338 462774 30574
rect 462154 12894 462774 30338
rect 462154 12658 462186 12894
rect 462422 12658 462506 12894
rect 462742 12658 462774 12894
rect 462154 12574 462774 12658
rect 462154 12338 462186 12574
rect 462422 12338 462506 12574
rect 462742 12338 462774 12574
rect 462154 -2776 462774 12338
rect 462154 -3012 462186 -2776
rect 462422 -3012 462506 -2776
rect 462742 -3012 462774 -2776
rect 462154 -3096 462774 -3012
rect 462154 -3332 462186 -3096
rect 462422 -3332 462506 -3096
rect 462742 -3332 462774 -3096
rect 462154 -4324 462774 -3332
rect 465874 463972 466494 464004
rect 465874 463736 465906 463972
rect 466142 463736 466226 463972
rect 466462 463736 466494 463972
rect 465874 463652 466494 463736
rect 465874 463416 465906 463652
rect 466142 463416 466226 463652
rect 466462 463416 466494 463652
rect 465874 448614 466494 463416
rect 465874 448378 465906 448614
rect 466142 448378 466226 448614
rect 466462 448378 466494 448614
rect 465874 448294 466494 448378
rect 465874 448058 465906 448294
rect 466142 448058 466226 448294
rect 466462 448058 466494 448294
rect 465874 430614 466494 448058
rect 465874 430378 465906 430614
rect 466142 430378 466226 430614
rect 466462 430378 466494 430614
rect 465874 430294 466494 430378
rect 465874 430058 465906 430294
rect 466142 430058 466226 430294
rect 466462 430058 466494 430294
rect 465874 412614 466494 430058
rect 465874 412378 465906 412614
rect 466142 412378 466226 412614
rect 466462 412378 466494 412614
rect 465874 412294 466494 412378
rect 465874 412058 465906 412294
rect 466142 412058 466226 412294
rect 466462 412058 466494 412294
rect 465874 394614 466494 412058
rect 465874 394378 465906 394614
rect 466142 394378 466226 394614
rect 466462 394378 466494 394614
rect 465874 394294 466494 394378
rect 465874 394058 465906 394294
rect 466142 394058 466226 394294
rect 466462 394058 466494 394294
rect 465874 376614 466494 394058
rect 465874 376378 465906 376614
rect 466142 376378 466226 376614
rect 466462 376378 466494 376614
rect 465874 376294 466494 376378
rect 465874 376058 465906 376294
rect 466142 376058 466226 376294
rect 466462 376058 466494 376294
rect 465874 358614 466494 376058
rect 465874 358378 465906 358614
rect 466142 358378 466226 358614
rect 466462 358378 466494 358614
rect 465874 358294 466494 358378
rect 465874 358058 465906 358294
rect 466142 358058 466226 358294
rect 466462 358058 466494 358294
rect 465874 340614 466494 358058
rect 465874 340378 465906 340614
rect 466142 340378 466226 340614
rect 466462 340378 466494 340614
rect 465874 340294 466494 340378
rect 465874 340058 465906 340294
rect 466142 340058 466226 340294
rect 466462 340058 466494 340294
rect 465874 322614 466494 340058
rect 465874 322378 465906 322614
rect 466142 322378 466226 322614
rect 466462 322378 466494 322614
rect 465874 322294 466494 322378
rect 465874 322058 465906 322294
rect 466142 322058 466226 322294
rect 466462 322058 466494 322294
rect 465874 304614 466494 322058
rect 465874 304378 465906 304614
rect 466142 304378 466226 304614
rect 466462 304378 466494 304614
rect 465874 304294 466494 304378
rect 465874 304058 465906 304294
rect 466142 304058 466226 304294
rect 466462 304058 466494 304294
rect 465874 286614 466494 304058
rect 465874 286378 465906 286614
rect 466142 286378 466226 286614
rect 466462 286378 466494 286614
rect 465874 286294 466494 286378
rect 465874 286058 465906 286294
rect 466142 286058 466226 286294
rect 466462 286058 466494 286294
rect 465874 268614 466494 286058
rect 465874 268378 465906 268614
rect 466142 268378 466226 268614
rect 466462 268378 466494 268614
rect 465874 268294 466494 268378
rect 465874 268058 465906 268294
rect 466142 268058 466226 268294
rect 466462 268058 466494 268294
rect 465874 250614 466494 268058
rect 465874 250378 465906 250614
rect 466142 250378 466226 250614
rect 466462 250378 466494 250614
rect 465874 250294 466494 250378
rect 465874 250058 465906 250294
rect 466142 250058 466226 250294
rect 466462 250058 466494 250294
rect 465874 232614 466494 250058
rect 465874 232378 465906 232614
rect 466142 232378 466226 232614
rect 466462 232378 466494 232614
rect 465874 232294 466494 232378
rect 465874 232058 465906 232294
rect 466142 232058 466226 232294
rect 466462 232058 466494 232294
rect 465874 214614 466494 232058
rect 465874 214378 465906 214614
rect 466142 214378 466226 214614
rect 466462 214378 466494 214614
rect 465874 214294 466494 214378
rect 465874 214058 465906 214294
rect 466142 214058 466226 214294
rect 466462 214058 466494 214294
rect 465874 196614 466494 214058
rect 465874 196378 465906 196614
rect 466142 196378 466226 196614
rect 466462 196378 466494 196614
rect 465874 196294 466494 196378
rect 465874 196058 465906 196294
rect 466142 196058 466226 196294
rect 466462 196058 466494 196294
rect 465874 178614 466494 196058
rect 465874 178378 465906 178614
rect 466142 178378 466226 178614
rect 466462 178378 466494 178614
rect 465874 178294 466494 178378
rect 465874 178058 465906 178294
rect 466142 178058 466226 178294
rect 466462 178058 466494 178294
rect 465874 160614 466494 178058
rect 465874 160378 465906 160614
rect 466142 160378 466226 160614
rect 466462 160378 466494 160614
rect 465874 160294 466494 160378
rect 465874 160058 465906 160294
rect 466142 160058 466226 160294
rect 466462 160058 466494 160294
rect 465874 142614 466494 160058
rect 465874 142378 465906 142614
rect 466142 142378 466226 142614
rect 466462 142378 466494 142614
rect 465874 142294 466494 142378
rect 465874 142058 465906 142294
rect 466142 142058 466226 142294
rect 466462 142058 466494 142294
rect 465874 124614 466494 142058
rect 465874 124378 465906 124614
rect 466142 124378 466226 124614
rect 466462 124378 466494 124614
rect 465874 124294 466494 124378
rect 465874 124058 465906 124294
rect 466142 124058 466226 124294
rect 466462 124058 466494 124294
rect 465874 106614 466494 124058
rect 465874 106378 465906 106614
rect 466142 106378 466226 106614
rect 466462 106378 466494 106614
rect 465874 106294 466494 106378
rect 465874 106058 465906 106294
rect 466142 106058 466226 106294
rect 466462 106058 466494 106294
rect 465874 88614 466494 106058
rect 465874 88378 465906 88614
rect 466142 88378 466226 88614
rect 466462 88378 466494 88614
rect 465874 88294 466494 88378
rect 465874 88058 465906 88294
rect 466142 88058 466226 88294
rect 466462 88058 466494 88294
rect 465874 70614 466494 88058
rect 465874 70378 465906 70614
rect 466142 70378 466226 70614
rect 466462 70378 466494 70614
rect 465874 70294 466494 70378
rect 465874 70058 465906 70294
rect 466142 70058 466226 70294
rect 466462 70058 466494 70294
rect 465874 52614 466494 70058
rect 465874 52378 465906 52614
rect 466142 52378 466226 52614
rect 466462 52378 466494 52614
rect 465874 52294 466494 52378
rect 465874 52058 465906 52294
rect 466142 52058 466226 52294
rect 466462 52058 466494 52294
rect 465874 34614 466494 52058
rect 465874 34378 465906 34614
rect 466142 34378 466226 34614
rect 466462 34378 466494 34614
rect 465874 34294 466494 34378
rect 465874 34058 465906 34294
rect 466142 34058 466226 34294
rect 466462 34058 466494 34294
rect 465874 16614 466494 34058
rect 465874 16378 465906 16614
rect 466142 16378 466226 16614
rect 466462 16378 466494 16614
rect 465874 16294 466494 16378
rect 465874 16058 465906 16294
rect 466142 16058 466226 16294
rect 466462 16058 466494 16294
rect 465874 -3736 466494 16058
rect 465874 -3972 465906 -3736
rect 466142 -3972 466226 -3736
rect 466462 -3972 466494 -3736
rect 465874 -4056 466494 -3972
rect 465874 -4292 465906 -4056
rect 466142 -4292 466226 -4056
rect 466462 -4292 466494 -4056
rect 465874 -4324 466494 -4292
rect 472714 461092 473334 464004
rect 472714 460856 472746 461092
rect 472982 460856 473066 461092
rect 473302 460856 473334 461092
rect 472714 460772 473334 460856
rect 472714 460536 472746 460772
rect 472982 460536 473066 460772
rect 473302 460536 473334 460772
rect 472714 455454 473334 460536
rect 472714 455218 472746 455454
rect 472982 455218 473066 455454
rect 473302 455218 473334 455454
rect 472714 455134 473334 455218
rect 472714 454898 472746 455134
rect 472982 454898 473066 455134
rect 473302 454898 473334 455134
rect 472714 437454 473334 454898
rect 472714 437218 472746 437454
rect 472982 437218 473066 437454
rect 473302 437218 473334 437454
rect 472714 437134 473334 437218
rect 472714 436898 472746 437134
rect 472982 436898 473066 437134
rect 473302 436898 473334 437134
rect 472714 419454 473334 436898
rect 472714 419218 472746 419454
rect 472982 419218 473066 419454
rect 473302 419218 473334 419454
rect 472714 419134 473334 419218
rect 472714 418898 472746 419134
rect 472982 418898 473066 419134
rect 473302 418898 473334 419134
rect 472714 401454 473334 418898
rect 472714 401218 472746 401454
rect 472982 401218 473066 401454
rect 473302 401218 473334 401454
rect 472714 401134 473334 401218
rect 472714 400898 472746 401134
rect 472982 400898 473066 401134
rect 473302 400898 473334 401134
rect 472714 383454 473334 400898
rect 472714 383218 472746 383454
rect 472982 383218 473066 383454
rect 473302 383218 473334 383454
rect 472714 383134 473334 383218
rect 472714 382898 472746 383134
rect 472982 382898 473066 383134
rect 473302 382898 473334 383134
rect 472714 365454 473334 382898
rect 472714 365218 472746 365454
rect 472982 365218 473066 365454
rect 473302 365218 473334 365454
rect 472714 365134 473334 365218
rect 472714 364898 472746 365134
rect 472982 364898 473066 365134
rect 473302 364898 473334 365134
rect 472714 347454 473334 364898
rect 472714 347218 472746 347454
rect 472982 347218 473066 347454
rect 473302 347218 473334 347454
rect 472714 347134 473334 347218
rect 472714 346898 472746 347134
rect 472982 346898 473066 347134
rect 473302 346898 473334 347134
rect 472714 329454 473334 346898
rect 472714 329218 472746 329454
rect 472982 329218 473066 329454
rect 473302 329218 473334 329454
rect 472714 329134 473334 329218
rect 472714 328898 472746 329134
rect 472982 328898 473066 329134
rect 473302 328898 473334 329134
rect 472714 311454 473334 328898
rect 472714 311218 472746 311454
rect 472982 311218 473066 311454
rect 473302 311218 473334 311454
rect 472714 311134 473334 311218
rect 472714 310898 472746 311134
rect 472982 310898 473066 311134
rect 473302 310898 473334 311134
rect 472714 293454 473334 310898
rect 472714 293218 472746 293454
rect 472982 293218 473066 293454
rect 473302 293218 473334 293454
rect 472714 293134 473334 293218
rect 472714 292898 472746 293134
rect 472982 292898 473066 293134
rect 473302 292898 473334 293134
rect 472714 275454 473334 292898
rect 472714 275218 472746 275454
rect 472982 275218 473066 275454
rect 473302 275218 473334 275454
rect 472714 275134 473334 275218
rect 472714 274898 472746 275134
rect 472982 274898 473066 275134
rect 473302 274898 473334 275134
rect 472714 257454 473334 274898
rect 472714 257218 472746 257454
rect 472982 257218 473066 257454
rect 473302 257218 473334 257454
rect 472714 257134 473334 257218
rect 472714 256898 472746 257134
rect 472982 256898 473066 257134
rect 473302 256898 473334 257134
rect 472714 239454 473334 256898
rect 472714 239218 472746 239454
rect 472982 239218 473066 239454
rect 473302 239218 473334 239454
rect 472714 239134 473334 239218
rect 472714 238898 472746 239134
rect 472982 238898 473066 239134
rect 473302 238898 473334 239134
rect 472714 221454 473334 238898
rect 472714 221218 472746 221454
rect 472982 221218 473066 221454
rect 473302 221218 473334 221454
rect 472714 221134 473334 221218
rect 472714 220898 472746 221134
rect 472982 220898 473066 221134
rect 473302 220898 473334 221134
rect 472714 203454 473334 220898
rect 472714 203218 472746 203454
rect 472982 203218 473066 203454
rect 473302 203218 473334 203454
rect 472714 203134 473334 203218
rect 472714 202898 472746 203134
rect 472982 202898 473066 203134
rect 473302 202898 473334 203134
rect 472714 185454 473334 202898
rect 472714 185218 472746 185454
rect 472982 185218 473066 185454
rect 473302 185218 473334 185454
rect 472714 185134 473334 185218
rect 472714 184898 472746 185134
rect 472982 184898 473066 185134
rect 473302 184898 473334 185134
rect 472714 167454 473334 184898
rect 472714 167218 472746 167454
rect 472982 167218 473066 167454
rect 473302 167218 473334 167454
rect 472714 167134 473334 167218
rect 472714 166898 472746 167134
rect 472982 166898 473066 167134
rect 473302 166898 473334 167134
rect 472714 149454 473334 166898
rect 472714 149218 472746 149454
rect 472982 149218 473066 149454
rect 473302 149218 473334 149454
rect 472714 149134 473334 149218
rect 472714 148898 472746 149134
rect 472982 148898 473066 149134
rect 473302 148898 473334 149134
rect 472714 131454 473334 148898
rect 472714 131218 472746 131454
rect 472982 131218 473066 131454
rect 473302 131218 473334 131454
rect 472714 131134 473334 131218
rect 472714 130898 472746 131134
rect 472982 130898 473066 131134
rect 473302 130898 473334 131134
rect 472714 113454 473334 130898
rect 472714 113218 472746 113454
rect 472982 113218 473066 113454
rect 473302 113218 473334 113454
rect 472714 113134 473334 113218
rect 472714 112898 472746 113134
rect 472982 112898 473066 113134
rect 473302 112898 473334 113134
rect 472714 95454 473334 112898
rect 472714 95218 472746 95454
rect 472982 95218 473066 95454
rect 473302 95218 473334 95454
rect 472714 95134 473334 95218
rect 472714 94898 472746 95134
rect 472982 94898 473066 95134
rect 473302 94898 473334 95134
rect 472714 77454 473334 94898
rect 472714 77218 472746 77454
rect 472982 77218 473066 77454
rect 473302 77218 473334 77454
rect 472714 77134 473334 77218
rect 472714 76898 472746 77134
rect 472982 76898 473066 77134
rect 473302 76898 473334 77134
rect 472714 59454 473334 76898
rect 472714 59218 472746 59454
rect 472982 59218 473066 59454
rect 473302 59218 473334 59454
rect 472714 59134 473334 59218
rect 472714 58898 472746 59134
rect 472982 58898 473066 59134
rect 473302 58898 473334 59134
rect 472714 41454 473334 58898
rect 472714 41218 472746 41454
rect 472982 41218 473066 41454
rect 473302 41218 473334 41454
rect 472714 41134 473334 41218
rect 472714 40898 472746 41134
rect 472982 40898 473066 41134
rect 473302 40898 473334 41134
rect 472714 23454 473334 40898
rect 472714 23218 472746 23454
rect 472982 23218 473066 23454
rect 473302 23218 473334 23454
rect 472714 23134 473334 23218
rect 472714 22898 472746 23134
rect 472982 22898 473066 23134
rect 473302 22898 473334 23134
rect 472714 5454 473334 22898
rect 472714 5218 472746 5454
rect 472982 5218 473066 5454
rect 473302 5218 473334 5454
rect 472714 5134 473334 5218
rect 472714 4898 472746 5134
rect 472982 4898 473066 5134
rect 473302 4898 473334 5134
rect 472714 -856 473334 4898
rect 472714 -1092 472746 -856
rect 472982 -1092 473066 -856
rect 473302 -1092 473334 -856
rect 472714 -1176 473334 -1092
rect 472714 -1412 472746 -1176
rect 472982 -1412 473066 -1176
rect 473302 -1412 473334 -1176
rect 472714 -4324 473334 -1412
rect 476434 462052 477054 464004
rect 476434 461816 476466 462052
rect 476702 461816 476786 462052
rect 477022 461816 477054 462052
rect 476434 461732 477054 461816
rect 476434 461496 476466 461732
rect 476702 461496 476786 461732
rect 477022 461496 477054 461732
rect 476434 441174 477054 461496
rect 476434 440938 476466 441174
rect 476702 440938 476786 441174
rect 477022 440938 477054 441174
rect 476434 440854 477054 440938
rect 476434 440618 476466 440854
rect 476702 440618 476786 440854
rect 477022 440618 477054 440854
rect 476434 423174 477054 440618
rect 476434 422938 476466 423174
rect 476702 422938 476786 423174
rect 477022 422938 477054 423174
rect 476434 422854 477054 422938
rect 476434 422618 476466 422854
rect 476702 422618 476786 422854
rect 477022 422618 477054 422854
rect 476434 405174 477054 422618
rect 476434 404938 476466 405174
rect 476702 404938 476786 405174
rect 477022 404938 477054 405174
rect 476434 404854 477054 404938
rect 476434 404618 476466 404854
rect 476702 404618 476786 404854
rect 477022 404618 477054 404854
rect 476434 387174 477054 404618
rect 476434 386938 476466 387174
rect 476702 386938 476786 387174
rect 477022 386938 477054 387174
rect 476434 386854 477054 386938
rect 476434 386618 476466 386854
rect 476702 386618 476786 386854
rect 477022 386618 477054 386854
rect 476434 369174 477054 386618
rect 476434 368938 476466 369174
rect 476702 368938 476786 369174
rect 477022 368938 477054 369174
rect 476434 368854 477054 368938
rect 476434 368618 476466 368854
rect 476702 368618 476786 368854
rect 477022 368618 477054 368854
rect 476434 351174 477054 368618
rect 476434 350938 476466 351174
rect 476702 350938 476786 351174
rect 477022 350938 477054 351174
rect 476434 350854 477054 350938
rect 476434 350618 476466 350854
rect 476702 350618 476786 350854
rect 477022 350618 477054 350854
rect 476434 333174 477054 350618
rect 476434 332938 476466 333174
rect 476702 332938 476786 333174
rect 477022 332938 477054 333174
rect 476434 332854 477054 332938
rect 476434 332618 476466 332854
rect 476702 332618 476786 332854
rect 477022 332618 477054 332854
rect 476434 315174 477054 332618
rect 476434 314938 476466 315174
rect 476702 314938 476786 315174
rect 477022 314938 477054 315174
rect 476434 314854 477054 314938
rect 476434 314618 476466 314854
rect 476702 314618 476786 314854
rect 477022 314618 477054 314854
rect 476434 297174 477054 314618
rect 476434 296938 476466 297174
rect 476702 296938 476786 297174
rect 477022 296938 477054 297174
rect 476434 296854 477054 296938
rect 476434 296618 476466 296854
rect 476702 296618 476786 296854
rect 477022 296618 477054 296854
rect 476434 279174 477054 296618
rect 476434 278938 476466 279174
rect 476702 278938 476786 279174
rect 477022 278938 477054 279174
rect 476434 278854 477054 278938
rect 476434 278618 476466 278854
rect 476702 278618 476786 278854
rect 477022 278618 477054 278854
rect 476434 261174 477054 278618
rect 476434 260938 476466 261174
rect 476702 260938 476786 261174
rect 477022 260938 477054 261174
rect 476434 260854 477054 260938
rect 476434 260618 476466 260854
rect 476702 260618 476786 260854
rect 477022 260618 477054 260854
rect 476434 243174 477054 260618
rect 476434 242938 476466 243174
rect 476702 242938 476786 243174
rect 477022 242938 477054 243174
rect 476434 242854 477054 242938
rect 476434 242618 476466 242854
rect 476702 242618 476786 242854
rect 477022 242618 477054 242854
rect 476434 225174 477054 242618
rect 476434 224938 476466 225174
rect 476702 224938 476786 225174
rect 477022 224938 477054 225174
rect 476434 224854 477054 224938
rect 476434 224618 476466 224854
rect 476702 224618 476786 224854
rect 477022 224618 477054 224854
rect 476434 207174 477054 224618
rect 476434 206938 476466 207174
rect 476702 206938 476786 207174
rect 477022 206938 477054 207174
rect 476434 206854 477054 206938
rect 476434 206618 476466 206854
rect 476702 206618 476786 206854
rect 477022 206618 477054 206854
rect 476434 189174 477054 206618
rect 476434 188938 476466 189174
rect 476702 188938 476786 189174
rect 477022 188938 477054 189174
rect 476434 188854 477054 188938
rect 476434 188618 476466 188854
rect 476702 188618 476786 188854
rect 477022 188618 477054 188854
rect 476434 171174 477054 188618
rect 476434 170938 476466 171174
rect 476702 170938 476786 171174
rect 477022 170938 477054 171174
rect 476434 170854 477054 170938
rect 476434 170618 476466 170854
rect 476702 170618 476786 170854
rect 477022 170618 477054 170854
rect 476434 153174 477054 170618
rect 476434 152938 476466 153174
rect 476702 152938 476786 153174
rect 477022 152938 477054 153174
rect 476434 152854 477054 152938
rect 476434 152618 476466 152854
rect 476702 152618 476786 152854
rect 477022 152618 477054 152854
rect 476434 135174 477054 152618
rect 476434 134938 476466 135174
rect 476702 134938 476786 135174
rect 477022 134938 477054 135174
rect 476434 134854 477054 134938
rect 476434 134618 476466 134854
rect 476702 134618 476786 134854
rect 477022 134618 477054 134854
rect 476434 117174 477054 134618
rect 476434 116938 476466 117174
rect 476702 116938 476786 117174
rect 477022 116938 477054 117174
rect 476434 116854 477054 116938
rect 476434 116618 476466 116854
rect 476702 116618 476786 116854
rect 477022 116618 477054 116854
rect 476434 99174 477054 116618
rect 476434 98938 476466 99174
rect 476702 98938 476786 99174
rect 477022 98938 477054 99174
rect 476434 98854 477054 98938
rect 476434 98618 476466 98854
rect 476702 98618 476786 98854
rect 477022 98618 477054 98854
rect 476434 81174 477054 98618
rect 476434 80938 476466 81174
rect 476702 80938 476786 81174
rect 477022 80938 477054 81174
rect 476434 80854 477054 80938
rect 476434 80618 476466 80854
rect 476702 80618 476786 80854
rect 477022 80618 477054 80854
rect 476434 63174 477054 80618
rect 476434 62938 476466 63174
rect 476702 62938 476786 63174
rect 477022 62938 477054 63174
rect 476434 62854 477054 62938
rect 476434 62618 476466 62854
rect 476702 62618 476786 62854
rect 477022 62618 477054 62854
rect 476434 45174 477054 62618
rect 476434 44938 476466 45174
rect 476702 44938 476786 45174
rect 477022 44938 477054 45174
rect 476434 44854 477054 44938
rect 476434 44618 476466 44854
rect 476702 44618 476786 44854
rect 477022 44618 477054 44854
rect 476434 27174 477054 44618
rect 476434 26938 476466 27174
rect 476702 26938 476786 27174
rect 477022 26938 477054 27174
rect 476434 26854 477054 26938
rect 476434 26618 476466 26854
rect 476702 26618 476786 26854
rect 477022 26618 477054 26854
rect 476434 9174 477054 26618
rect 476434 8938 476466 9174
rect 476702 8938 476786 9174
rect 477022 8938 477054 9174
rect 476434 8854 477054 8938
rect 476434 8618 476466 8854
rect 476702 8618 476786 8854
rect 477022 8618 477054 8854
rect 476434 -1816 477054 8618
rect 476434 -2052 476466 -1816
rect 476702 -2052 476786 -1816
rect 477022 -2052 477054 -1816
rect 476434 -2136 477054 -2052
rect 476434 -2372 476466 -2136
rect 476702 -2372 476786 -2136
rect 477022 -2372 477054 -2136
rect 476434 -4324 477054 -2372
rect 480154 463012 480774 464004
rect 480154 462776 480186 463012
rect 480422 462776 480506 463012
rect 480742 462776 480774 463012
rect 480154 462692 480774 462776
rect 480154 462456 480186 462692
rect 480422 462456 480506 462692
rect 480742 462456 480774 462692
rect 480154 444894 480774 462456
rect 480154 444658 480186 444894
rect 480422 444658 480506 444894
rect 480742 444658 480774 444894
rect 480154 444574 480774 444658
rect 480154 444338 480186 444574
rect 480422 444338 480506 444574
rect 480742 444338 480774 444574
rect 480154 426894 480774 444338
rect 480154 426658 480186 426894
rect 480422 426658 480506 426894
rect 480742 426658 480774 426894
rect 480154 426574 480774 426658
rect 480154 426338 480186 426574
rect 480422 426338 480506 426574
rect 480742 426338 480774 426574
rect 480154 408894 480774 426338
rect 480154 408658 480186 408894
rect 480422 408658 480506 408894
rect 480742 408658 480774 408894
rect 480154 408574 480774 408658
rect 480154 408338 480186 408574
rect 480422 408338 480506 408574
rect 480742 408338 480774 408574
rect 480154 390894 480774 408338
rect 480154 390658 480186 390894
rect 480422 390658 480506 390894
rect 480742 390658 480774 390894
rect 480154 390574 480774 390658
rect 480154 390338 480186 390574
rect 480422 390338 480506 390574
rect 480742 390338 480774 390574
rect 480154 372894 480774 390338
rect 480154 372658 480186 372894
rect 480422 372658 480506 372894
rect 480742 372658 480774 372894
rect 480154 372574 480774 372658
rect 480154 372338 480186 372574
rect 480422 372338 480506 372574
rect 480742 372338 480774 372574
rect 480154 354894 480774 372338
rect 480154 354658 480186 354894
rect 480422 354658 480506 354894
rect 480742 354658 480774 354894
rect 480154 354574 480774 354658
rect 480154 354338 480186 354574
rect 480422 354338 480506 354574
rect 480742 354338 480774 354574
rect 480154 336894 480774 354338
rect 480154 336658 480186 336894
rect 480422 336658 480506 336894
rect 480742 336658 480774 336894
rect 480154 336574 480774 336658
rect 480154 336338 480186 336574
rect 480422 336338 480506 336574
rect 480742 336338 480774 336574
rect 480154 318894 480774 336338
rect 480154 318658 480186 318894
rect 480422 318658 480506 318894
rect 480742 318658 480774 318894
rect 480154 318574 480774 318658
rect 480154 318338 480186 318574
rect 480422 318338 480506 318574
rect 480742 318338 480774 318574
rect 480154 300894 480774 318338
rect 480154 300658 480186 300894
rect 480422 300658 480506 300894
rect 480742 300658 480774 300894
rect 480154 300574 480774 300658
rect 480154 300338 480186 300574
rect 480422 300338 480506 300574
rect 480742 300338 480774 300574
rect 480154 282894 480774 300338
rect 480154 282658 480186 282894
rect 480422 282658 480506 282894
rect 480742 282658 480774 282894
rect 480154 282574 480774 282658
rect 480154 282338 480186 282574
rect 480422 282338 480506 282574
rect 480742 282338 480774 282574
rect 480154 264894 480774 282338
rect 480154 264658 480186 264894
rect 480422 264658 480506 264894
rect 480742 264658 480774 264894
rect 480154 264574 480774 264658
rect 480154 264338 480186 264574
rect 480422 264338 480506 264574
rect 480742 264338 480774 264574
rect 480154 246894 480774 264338
rect 480154 246658 480186 246894
rect 480422 246658 480506 246894
rect 480742 246658 480774 246894
rect 480154 246574 480774 246658
rect 480154 246338 480186 246574
rect 480422 246338 480506 246574
rect 480742 246338 480774 246574
rect 480154 228894 480774 246338
rect 480154 228658 480186 228894
rect 480422 228658 480506 228894
rect 480742 228658 480774 228894
rect 480154 228574 480774 228658
rect 480154 228338 480186 228574
rect 480422 228338 480506 228574
rect 480742 228338 480774 228574
rect 480154 210894 480774 228338
rect 480154 210658 480186 210894
rect 480422 210658 480506 210894
rect 480742 210658 480774 210894
rect 480154 210574 480774 210658
rect 480154 210338 480186 210574
rect 480422 210338 480506 210574
rect 480742 210338 480774 210574
rect 480154 192894 480774 210338
rect 480154 192658 480186 192894
rect 480422 192658 480506 192894
rect 480742 192658 480774 192894
rect 480154 192574 480774 192658
rect 480154 192338 480186 192574
rect 480422 192338 480506 192574
rect 480742 192338 480774 192574
rect 480154 174894 480774 192338
rect 480154 174658 480186 174894
rect 480422 174658 480506 174894
rect 480742 174658 480774 174894
rect 480154 174574 480774 174658
rect 480154 174338 480186 174574
rect 480422 174338 480506 174574
rect 480742 174338 480774 174574
rect 480154 156894 480774 174338
rect 480154 156658 480186 156894
rect 480422 156658 480506 156894
rect 480742 156658 480774 156894
rect 480154 156574 480774 156658
rect 480154 156338 480186 156574
rect 480422 156338 480506 156574
rect 480742 156338 480774 156574
rect 480154 138894 480774 156338
rect 480154 138658 480186 138894
rect 480422 138658 480506 138894
rect 480742 138658 480774 138894
rect 480154 138574 480774 138658
rect 480154 138338 480186 138574
rect 480422 138338 480506 138574
rect 480742 138338 480774 138574
rect 480154 120894 480774 138338
rect 480154 120658 480186 120894
rect 480422 120658 480506 120894
rect 480742 120658 480774 120894
rect 480154 120574 480774 120658
rect 480154 120338 480186 120574
rect 480422 120338 480506 120574
rect 480742 120338 480774 120574
rect 480154 102894 480774 120338
rect 480154 102658 480186 102894
rect 480422 102658 480506 102894
rect 480742 102658 480774 102894
rect 480154 102574 480774 102658
rect 480154 102338 480186 102574
rect 480422 102338 480506 102574
rect 480742 102338 480774 102574
rect 480154 84894 480774 102338
rect 480154 84658 480186 84894
rect 480422 84658 480506 84894
rect 480742 84658 480774 84894
rect 480154 84574 480774 84658
rect 480154 84338 480186 84574
rect 480422 84338 480506 84574
rect 480742 84338 480774 84574
rect 480154 66894 480774 84338
rect 480154 66658 480186 66894
rect 480422 66658 480506 66894
rect 480742 66658 480774 66894
rect 480154 66574 480774 66658
rect 480154 66338 480186 66574
rect 480422 66338 480506 66574
rect 480742 66338 480774 66574
rect 480154 48894 480774 66338
rect 480154 48658 480186 48894
rect 480422 48658 480506 48894
rect 480742 48658 480774 48894
rect 480154 48574 480774 48658
rect 480154 48338 480186 48574
rect 480422 48338 480506 48574
rect 480742 48338 480774 48574
rect 480154 30894 480774 48338
rect 480154 30658 480186 30894
rect 480422 30658 480506 30894
rect 480742 30658 480774 30894
rect 480154 30574 480774 30658
rect 480154 30338 480186 30574
rect 480422 30338 480506 30574
rect 480742 30338 480774 30574
rect 480154 12894 480774 30338
rect 480154 12658 480186 12894
rect 480422 12658 480506 12894
rect 480742 12658 480774 12894
rect 480154 12574 480774 12658
rect 480154 12338 480186 12574
rect 480422 12338 480506 12574
rect 480742 12338 480774 12574
rect 480154 -2776 480774 12338
rect 480154 -3012 480186 -2776
rect 480422 -3012 480506 -2776
rect 480742 -3012 480774 -2776
rect 480154 -3096 480774 -3012
rect 480154 -3332 480186 -3096
rect 480422 -3332 480506 -3096
rect 480742 -3332 480774 -3096
rect 480154 -4324 480774 -3332
rect 483874 463972 484494 464004
rect 483874 463736 483906 463972
rect 484142 463736 484226 463972
rect 484462 463736 484494 463972
rect 483874 463652 484494 463736
rect 483874 463416 483906 463652
rect 484142 463416 484226 463652
rect 484462 463416 484494 463652
rect 483874 448614 484494 463416
rect 483874 448378 483906 448614
rect 484142 448378 484226 448614
rect 484462 448378 484494 448614
rect 483874 448294 484494 448378
rect 483874 448058 483906 448294
rect 484142 448058 484226 448294
rect 484462 448058 484494 448294
rect 483874 430614 484494 448058
rect 483874 430378 483906 430614
rect 484142 430378 484226 430614
rect 484462 430378 484494 430614
rect 483874 430294 484494 430378
rect 483874 430058 483906 430294
rect 484142 430058 484226 430294
rect 484462 430058 484494 430294
rect 483874 412614 484494 430058
rect 483874 412378 483906 412614
rect 484142 412378 484226 412614
rect 484462 412378 484494 412614
rect 483874 412294 484494 412378
rect 483874 412058 483906 412294
rect 484142 412058 484226 412294
rect 484462 412058 484494 412294
rect 483874 394614 484494 412058
rect 483874 394378 483906 394614
rect 484142 394378 484226 394614
rect 484462 394378 484494 394614
rect 483874 394294 484494 394378
rect 483874 394058 483906 394294
rect 484142 394058 484226 394294
rect 484462 394058 484494 394294
rect 483874 376614 484494 394058
rect 483874 376378 483906 376614
rect 484142 376378 484226 376614
rect 484462 376378 484494 376614
rect 483874 376294 484494 376378
rect 483874 376058 483906 376294
rect 484142 376058 484226 376294
rect 484462 376058 484494 376294
rect 483874 358614 484494 376058
rect 483874 358378 483906 358614
rect 484142 358378 484226 358614
rect 484462 358378 484494 358614
rect 483874 358294 484494 358378
rect 483874 358058 483906 358294
rect 484142 358058 484226 358294
rect 484462 358058 484494 358294
rect 483874 340614 484494 358058
rect 483874 340378 483906 340614
rect 484142 340378 484226 340614
rect 484462 340378 484494 340614
rect 483874 340294 484494 340378
rect 483874 340058 483906 340294
rect 484142 340058 484226 340294
rect 484462 340058 484494 340294
rect 483874 322614 484494 340058
rect 483874 322378 483906 322614
rect 484142 322378 484226 322614
rect 484462 322378 484494 322614
rect 483874 322294 484494 322378
rect 483874 322058 483906 322294
rect 484142 322058 484226 322294
rect 484462 322058 484494 322294
rect 483874 304614 484494 322058
rect 483874 304378 483906 304614
rect 484142 304378 484226 304614
rect 484462 304378 484494 304614
rect 483874 304294 484494 304378
rect 483874 304058 483906 304294
rect 484142 304058 484226 304294
rect 484462 304058 484494 304294
rect 483874 286614 484494 304058
rect 483874 286378 483906 286614
rect 484142 286378 484226 286614
rect 484462 286378 484494 286614
rect 483874 286294 484494 286378
rect 483874 286058 483906 286294
rect 484142 286058 484226 286294
rect 484462 286058 484494 286294
rect 483874 268614 484494 286058
rect 483874 268378 483906 268614
rect 484142 268378 484226 268614
rect 484462 268378 484494 268614
rect 483874 268294 484494 268378
rect 483874 268058 483906 268294
rect 484142 268058 484226 268294
rect 484462 268058 484494 268294
rect 483874 250614 484494 268058
rect 483874 250378 483906 250614
rect 484142 250378 484226 250614
rect 484462 250378 484494 250614
rect 483874 250294 484494 250378
rect 483874 250058 483906 250294
rect 484142 250058 484226 250294
rect 484462 250058 484494 250294
rect 483874 232614 484494 250058
rect 483874 232378 483906 232614
rect 484142 232378 484226 232614
rect 484462 232378 484494 232614
rect 483874 232294 484494 232378
rect 483874 232058 483906 232294
rect 484142 232058 484226 232294
rect 484462 232058 484494 232294
rect 483874 214614 484494 232058
rect 483874 214378 483906 214614
rect 484142 214378 484226 214614
rect 484462 214378 484494 214614
rect 483874 214294 484494 214378
rect 483874 214058 483906 214294
rect 484142 214058 484226 214294
rect 484462 214058 484494 214294
rect 483874 196614 484494 214058
rect 483874 196378 483906 196614
rect 484142 196378 484226 196614
rect 484462 196378 484494 196614
rect 483874 196294 484494 196378
rect 483874 196058 483906 196294
rect 484142 196058 484226 196294
rect 484462 196058 484494 196294
rect 483874 178614 484494 196058
rect 483874 178378 483906 178614
rect 484142 178378 484226 178614
rect 484462 178378 484494 178614
rect 483874 178294 484494 178378
rect 483874 178058 483906 178294
rect 484142 178058 484226 178294
rect 484462 178058 484494 178294
rect 483874 160614 484494 178058
rect 483874 160378 483906 160614
rect 484142 160378 484226 160614
rect 484462 160378 484494 160614
rect 483874 160294 484494 160378
rect 483874 160058 483906 160294
rect 484142 160058 484226 160294
rect 484462 160058 484494 160294
rect 483874 142614 484494 160058
rect 483874 142378 483906 142614
rect 484142 142378 484226 142614
rect 484462 142378 484494 142614
rect 483874 142294 484494 142378
rect 483874 142058 483906 142294
rect 484142 142058 484226 142294
rect 484462 142058 484494 142294
rect 483874 124614 484494 142058
rect 483874 124378 483906 124614
rect 484142 124378 484226 124614
rect 484462 124378 484494 124614
rect 483874 124294 484494 124378
rect 483874 124058 483906 124294
rect 484142 124058 484226 124294
rect 484462 124058 484494 124294
rect 483874 106614 484494 124058
rect 483874 106378 483906 106614
rect 484142 106378 484226 106614
rect 484462 106378 484494 106614
rect 483874 106294 484494 106378
rect 483874 106058 483906 106294
rect 484142 106058 484226 106294
rect 484462 106058 484494 106294
rect 483874 88614 484494 106058
rect 483874 88378 483906 88614
rect 484142 88378 484226 88614
rect 484462 88378 484494 88614
rect 483874 88294 484494 88378
rect 483874 88058 483906 88294
rect 484142 88058 484226 88294
rect 484462 88058 484494 88294
rect 483874 70614 484494 88058
rect 483874 70378 483906 70614
rect 484142 70378 484226 70614
rect 484462 70378 484494 70614
rect 483874 70294 484494 70378
rect 483874 70058 483906 70294
rect 484142 70058 484226 70294
rect 484462 70058 484494 70294
rect 483874 52614 484494 70058
rect 483874 52378 483906 52614
rect 484142 52378 484226 52614
rect 484462 52378 484494 52614
rect 483874 52294 484494 52378
rect 483874 52058 483906 52294
rect 484142 52058 484226 52294
rect 484462 52058 484494 52294
rect 483874 34614 484494 52058
rect 483874 34378 483906 34614
rect 484142 34378 484226 34614
rect 484462 34378 484494 34614
rect 483874 34294 484494 34378
rect 483874 34058 483906 34294
rect 484142 34058 484226 34294
rect 484462 34058 484494 34294
rect 483874 16614 484494 34058
rect 483874 16378 483906 16614
rect 484142 16378 484226 16614
rect 484462 16378 484494 16614
rect 483874 16294 484494 16378
rect 483874 16058 483906 16294
rect 484142 16058 484226 16294
rect 484462 16058 484494 16294
rect 483874 -3736 484494 16058
rect 483874 -3972 483906 -3736
rect 484142 -3972 484226 -3736
rect 484462 -3972 484494 -3736
rect 483874 -4056 484494 -3972
rect 483874 -4292 483906 -4056
rect 484142 -4292 484226 -4056
rect 484462 -4292 484494 -4056
rect 483874 -4324 484494 -4292
rect 490714 461092 491334 464004
rect 490714 460856 490746 461092
rect 490982 460856 491066 461092
rect 491302 460856 491334 461092
rect 490714 460772 491334 460856
rect 490714 460536 490746 460772
rect 490982 460536 491066 460772
rect 491302 460536 491334 460772
rect 490714 455454 491334 460536
rect 490714 455218 490746 455454
rect 490982 455218 491066 455454
rect 491302 455218 491334 455454
rect 490714 455134 491334 455218
rect 490714 454898 490746 455134
rect 490982 454898 491066 455134
rect 491302 454898 491334 455134
rect 490714 437454 491334 454898
rect 490714 437218 490746 437454
rect 490982 437218 491066 437454
rect 491302 437218 491334 437454
rect 490714 437134 491334 437218
rect 490714 436898 490746 437134
rect 490982 436898 491066 437134
rect 491302 436898 491334 437134
rect 490714 419454 491334 436898
rect 490714 419218 490746 419454
rect 490982 419218 491066 419454
rect 491302 419218 491334 419454
rect 490714 419134 491334 419218
rect 490714 418898 490746 419134
rect 490982 418898 491066 419134
rect 491302 418898 491334 419134
rect 490714 401454 491334 418898
rect 490714 401218 490746 401454
rect 490982 401218 491066 401454
rect 491302 401218 491334 401454
rect 490714 401134 491334 401218
rect 490714 400898 490746 401134
rect 490982 400898 491066 401134
rect 491302 400898 491334 401134
rect 490714 383454 491334 400898
rect 490714 383218 490746 383454
rect 490982 383218 491066 383454
rect 491302 383218 491334 383454
rect 490714 383134 491334 383218
rect 490714 382898 490746 383134
rect 490982 382898 491066 383134
rect 491302 382898 491334 383134
rect 490714 365454 491334 382898
rect 490714 365218 490746 365454
rect 490982 365218 491066 365454
rect 491302 365218 491334 365454
rect 490714 365134 491334 365218
rect 490714 364898 490746 365134
rect 490982 364898 491066 365134
rect 491302 364898 491334 365134
rect 490714 347454 491334 364898
rect 490714 347218 490746 347454
rect 490982 347218 491066 347454
rect 491302 347218 491334 347454
rect 490714 347134 491334 347218
rect 490714 346898 490746 347134
rect 490982 346898 491066 347134
rect 491302 346898 491334 347134
rect 490714 329454 491334 346898
rect 490714 329218 490746 329454
rect 490982 329218 491066 329454
rect 491302 329218 491334 329454
rect 490714 329134 491334 329218
rect 490714 328898 490746 329134
rect 490982 328898 491066 329134
rect 491302 328898 491334 329134
rect 490714 311454 491334 328898
rect 490714 311218 490746 311454
rect 490982 311218 491066 311454
rect 491302 311218 491334 311454
rect 490714 311134 491334 311218
rect 490714 310898 490746 311134
rect 490982 310898 491066 311134
rect 491302 310898 491334 311134
rect 490714 293454 491334 310898
rect 490714 293218 490746 293454
rect 490982 293218 491066 293454
rect 491302 293218 491334 293454
rect 490714 293134 491334 293218
rect 490714 292898 490746 293134
rect 490982 292898 491066 293134
rect 491302 292898 491334 293134
rect 490714 275454 491334 292898
rect 490714 275218 490746 275454
rect 490982 275218 491066 275454
rect 491302 275218 491334 275454
rect 490714 275134 491334 275218
rect 490714 274898 490746 275134
rect 490982 274898 491066 275134
rect 491302 274898 491334 275134
rect 490714 257454 491334 274898
rect 490714 257218 490746 257454
rect 490982 257218 491066 257454
rect 491302 257218 491334 257454
rect 490714 257134 491334 257218
rect 490714 256898 490746 257134
rect 490982 256898 491066 257134
rect 491302 256898 491334 257134
rect 490714 239454 491334 256898
rect 490714 239218 490746 239454
rect 490982 239218 491066 239454
rect 491302 239218 491334 239454
rect 490714 239134 491334 239218
rect 490714 238898 490746 239134
rect 490982 238898 491066 239134
rect 491302 238898 491334 239134
rect 490714 221454 491334 238898
rect 490714 221218 490746 221454
rect 490982 221218 491066 221454
rect 491302 221218 491334 221454
rect 490714 221134 491334 221218
rect 490714 220898 490746 221134
rect 490982 220898 491066 221134
rect 491302 220898 491334 221134
rect 490714 203454 491334 220898
rect 490714 203218 490746 203454
rect 490982 203218 491066 203454
rect 491302 203218 491334 203454
rect 490714 203134 491334 203218
rect 490714 202898 490746 203134
rect 490982 202898 491066 203134
rect 491302 202898 491334 203134
rect 490714 185454 491334 202898
rect 490714 185218 490746 185454
rect 490982 185218 491066 185454
rect 491302 185218 491334 185454
rect 490714 185134 491334 185218
rect 490714 184898 490746 185134
rect 490982 184898 491066 185134
rect 491302 184898 491334 185134
rect 490714 167454 491334 184898
rect 490714 167218 490746 167454
rect 490982 167218 491066 167454
rect 491302 167218 491334 167454
rect 490714 167134 491334 167218
rect 490714 166898 490746 167134
rect 490982 166898 491066 167134
rect 491302 166898 491334 167134
rect 490714 149454 491334 166898
rect 490714 149218 490746 149454
rect 490982 149218 491066 149454
rect 491302 149218 491334 149454
rect 490714 149134 491334 149218
rect 490714 148898 490746 149134
rect 490982 148898 491066 149134
rect 491302 148898 491334 149134
rect 490714 131454 491334 148898
rect 490714 131218 490746 131454
rect 490982 131218 491066 131454
rect 491302 131218 491334 131454
rect 490714 131134 491334 131218
rect 490714 130898 490746 131134
rect 490982 130898 491066 131134
rect 491302 130898 491334 131134
rect 490714 113454 491334 130898
rect 490714 113218 490746 113454
rect 490982 113218 491066 113454
rect 491302 113218 491334 113454
rect 490714 113134 491334 113218
rect 490714 112898 490746 113134
rect 490982 112898 491066 113134
rect 491302 112898 491334 113134
rect 490714 95454 491334 112898
rect 490714 95218 490746 95454
rect 490982 95218 491066 95454
rect 491302 95218 491334 95454
rect 490714 95134 491334 95218
rect 490714 94898 490746 95134
rect 490982 94898 491066 95134
rect 491302 94898 491334 95134
rect 490714 77454 491334 94898
rect 490714 77218 490746 77454
rect 490982 77218 491066 77454
rect 491302 77218 491334 77454
rect 490714 77134 491334 77218
rect 490714 76898 490746 77134
rect 490982 76898 491066 77134
rect 491302 76898 491334 77134
rect 490714 59454 491334 76898
rect 490714 59218 490746 59454
rect 490982 59218 491066 59454
rect 491302 59218 491334 59454
rect 490714 59134 491334 59218
rect 490714 58898 490746 59134
rect 490982 58898 491066 59134
rect 491302 58898 491334 59134
rect 490714 41454 491334 58898
rect 490714 41218 490746 41454
rect 490982 41218 491066 41454
rect 491302 41218 491334 41454
rect 490714 41134 491334 41218
rect 490714 40898 490746 41134
rect 490982 40898 491066 41134
rect 491302 40898 491334 41134
rect 490714 23454 491334 40898
rect 490714 23218 490746 23454
rect 490982 23218 491066 23454
rect 491302 23218 491334 23454
rect 490714 23134 491334 23218
rect 490714 22898 490746 23134
rect 490982 22898 491066 23134
rect 491302 22898 491334 23134
rect 490714 5454 491334 22898
rect 490714 5218 490746 5454
rect 490982 5218 491066 5454
rect 491302 5218 491334 5454
rect 490714 5134 491334 5218
rect 490714 4898 490746 5134
rect 490982 4898 491066 5134
rect 491302 4898 491334 5134
rect 490714 -856 491334 4898
rect 490714 -1092 490746 -856
rect 490982 -1092 491066 -856
rect 491302 -1092 491334 -856
rect 490714 -1176 491334 -1092
rect 490714 -1412 490746 -1176
rect 490982 -1412 491066 -1176
rect 491302 -1412 491334 -1176
rect 490714 -4324 491334 -1412
rect 494434 462052 495054 464004
rect 494434 461816 494466 462052
rect 494702 461816 494786 462052
rect 495022 461816 495054 462052
rect 494434 461732 495054 461816
rect 494434 461496 494466 461732
rect 494702 461496 494786 461732
rect 495022 461496 495054 461732
rect 494434 441174 495054 461496
rect 494434 440938 494466 441174
rect 494702 440938 494786 441174
rect 495022 440938 495054 441174
rect 494434 440854 495054 440938
rect 494434 440618 494466 440854
rect 494702 440618 494786 440854
rect 495022 440618 495054 440854
rect 494434 423174 495054 440618
rect 494434 422938 494466 423174
rect 494702 422938 494786 423174
rect 495022 422938 495054 423174
rect 494434 422854 495054 422938
rect 494434 422618 494466 422854
rect 494702 422618 494786 422854
rect 495022 422618 495054 422854
rect 494434 405174 495054 422618
rect 494434 404938 494466 405174
rect 494702 404938 494786 405174
rect 495022 404938 495054 405174
rect 494434 404854 495054 404938
rect 494434 404618 494466 404854
rect 494702 404618 494786 404854
rect 495022 404618 495054 404854
rect 494434 387174 495054 404618
rect 494434 386938 494466 387174
rect 494702 386938 494786 387174
rect 495022 386938 495054 387174
rect 494434 386854 495054 386938
rect 494434 386618 494466 386854
rect 494702 386618 494786 386854
rect 495022 386618 495054 386854
rect 494434 369174 495054 386618
rect 494434 368938 494466 369174
rect 494702 368938 494786 369174
rect 495022 368938 495054 369174
rect 494434 368854 495054 368938
rect 494434 368618 494466 368854
rect 494702 368618 494786 368854
rect 495022 368618 495054 368854
rect 494434 351174 495054 368618
rect 494434 350938 494466 351174
rect 494702 350938 494786 351174
rect 495022 350938 495054 351174
rect 494434 350854 495054 350938
rect 494434 350618 494466 350854
rect 494702 350618 494786 350854
rect 495022 350618 495054 350854
rect 494434 333174 495054 350618
rect 494434 332938 494466 333174
rect 494702 332938 494786 333174
rect 495022 332938 495054 333174
rect 494434 332854 495054 332938
rect 494434 332618 494466 332854
rect 494702 332618 494786 332854
rect 495022 332618 495054 332854
rect 494434 315174 495054 332618
rect 494434 314938 494466 315174
rect 494702 314938 494786 315174
rect 495022 314938 495054 315174
rect 494434 314854 495054 314938
rect 494434 314618 494466 314854
rect 494702 314618 494786 314854
rect 495022 314618 495054 314854
rect 494434 297174 495054 314618
rect 494434 296938 494466 297174
rect 494702 296938 494786 297174
rect 495022 296938 495054 297174
rect 494434 296854 495054 296938
rect 494434 296618 494466 296854
rect 494702 296618 494786 296854
rect 495022 296618 495054 296854
rect 494434 279174 495054 296618
rect 494434 278938 494466 279174
rect 494702 278938 494786 279174
rect 495022 278938 495054 279174
rect 494434 278854 495054 278938
rect 494434 278618 494466 278854
rect 494702 278618 494786 278854
rect 495022 278618 495054 278854
rect 494434 261174 495054 278618
rect 494434 260938 494466 261174
rect 494702 260938 494786 261174
rect 495022 260938 495054 261174
rect 494434 260854 495054 260938
rect 494434 260618 494466 260854
rect 494702 260618 494786 260854
rect 495022 260618 495054 260854
rect 494434 243174 495054 260618
rect 494434 242938 494466 243174
rect 494702 242938 494786 243174
rect 495022 242938 495054 243174
rect 494434 242854 495054 242938
rect 494434 242618 494466 242854
rect 494702 242618 494786 242854
rect 495022 242618 495054 242854
rect 494434 225174 495054 242618
rect 494434 224938 494466 225174
rect 494702 224938 494786 225174
rect 495022 224938 495054 225174
rect 494434 224854 495054 224938
rect 494434 224618 494466 224854
rect 494702 224618 494786 224854
rect 495022 224618 495054 224854
rect 494434 207174 495054 224618
rect 494434 206938 494466 207174
rect 494702 206938 494786 207174
rect 495022 206938 495054 207174
rect 494434 206854 495054 206938
rect 494434 206618 494466 206854
rect 494702 206618 494786 206854
rect 495022 206618 495054 206854
rect 494434 189174 495054 206618
rect 494434 188938 494466 189174
rect 494702 188938 494786 189174
rect 495022 188938 495054 189174
rect 494434 188854 495054 188938
rect 494434 188618 494466 188854
rect 494702 188618 494786 188854
rect 495022 188618 495054 188854
rect 494434 171174 495054 188618
rect 494434 170938 494466 171174
rect 494702 170938 494786 171174
rect 495022 170938 495054 171174
rect 494434 170854 495054 170938
rect 494434 170618 494466 170854
rect 494702 170618 494786 170854
rect 495022 170618 495054 170854
rect 494434 153174 495054 170618
rect 494434 152938 494466 153174
rect 494702 152938 494786 153174
rect 495022 152938 495054 153174
rect 494434 152854 495054 152938
rect 494434 152618 494466 152854
rect 494702 152618 494786 152854
rect 495022 152618 495054 152854
rect 494434 135174 495054 152618
rect 494434 134938 494466 135174
rect 494702 134938 494786 135174
rect 495022 134938 495054 135174
rect 494434 134854 495054 134938
rect 494434 134618 494466 134854
rect 494702 134618 494786 134854
rect 495022 134618 495054 134854
rect 494434 117174 495054 134618
rect 494434 116938 494466 117174
rect 494702 116938 494786 117174
rect 495022 116938 495054 117174
rect 494434 116854 495054 116938
rect 494434 116618 494466 116854
rect 494702 116618 494786 116854
rect 495022 116618 495054 116854
rect 494434 99174 495054 116618
rect 494434 98938 494466 99174
rect 494702 98938 494786 99174
rect 495022 98938 495054 99174
rect 494434 98854 495054 98938
rect 494434 98618 494466 98854
rect 494702 98618 494786 98854
rect 495022 98618 495054 98854
rect 494434 81174 495054 98618
rect 494434 80938 494466 81174
rect 494702 80938 494786 81174
rect 495022 80938 495054 81174
rect 494434 80854 495054 80938
rect 494434 80618 494466 80854
rect 494702 80618 494786 80854
rect 495022 80618 495054 80854
rect 494434 63174 495054 80618
rect 494434 62938 494466 63174
rect 494702 62938 494786 63174
rect 495022 62938 495054 63174
rect 494434 62854 495054 62938
rect 494434 62618 494466 62854
rect 494702 62618 494786 62854
rect 495022 62618 495054 62854
rect 494434 45174 495054 62618
rect 494434 44938 494466 45174
rect 494702 44938 494786 45174
rect 495022 44938 495054 45174
rect 494434 44854 495054 44938
rect 494434 44618 494466 44854
rect 494702 44618 494786 44854
rect 495022 44618 495054 44854
rect 494434 27174 495054 44618
rect 494434 26938 494466 27174
rect 494702 26938 494786 27174
rect 495022 26938 495054 27174
rect 494434 26854 495054 26938
rect 494434 26618 494466 26854
rect 494702 26618 494786 26854
rect 495022 26618 495054 26854
rect 494434 9174 495054 26618
rect 494434 8938 494466 9174
rect 494702 8938 494786 9174
rect 495022 8938 495054 9174
rect 494434 8854 495054 8938
rect 494434 8618 494466 8854
rect 494702 8618 494786 8854
rect 495022 8618 495054 8854
rect 494434 -1816 495054 8618
rect 494434 -2052 494466 -1816
rect 494702 -2052 494786 -1816
rect 495022 -2052 495054 -1816
rect 494434 -2136 495054 -2052
rect 494434 -2372 494466 -2136
rect 494702 -2372 494786 -2136
rect 495022 -2372 495054 -2136
rect 494434 -4324 495054 -2372
rect 498154 463012 498774 464004
rect 498154 462776 498186 463012
rect 498422 462776 498506 463012
rect 498742 462776 498774 463012
rect 498154 462692 498774 462776
rect 498154 462456 498186 462692
rect 498422 462456 498506 462692
rect 498742 462456 498774 462692
rect 498154 444894 498774 462456
rect 498154 444658 498186 444894
rect 498422 444658 498506 444894
rect 498742 444658 498774 444894
rect 498154 444574 498774 444658
rect 498154 444338 498186 444574
rect 498422 444338 498506 444574
rect 498742 444338 498774 444574
rect 498154 426894 498774 444338
rect 498154 426658 498186 426894
rect 498422 426658 498506 426894
rect 498742 426658 498774 426894
rect 498154 426574 498774 426658
rect 498154 426338 498186 426574
rect 498422 426338 498506 426574
rect 498742 426338 498774 426574
rect 498154 408894 498774 426338
rect 498154 408658 498186 408894
rect 498422 408658 498506 408894
rect 498742 408658 498774 408894
rect 498154 408574 498774 408658
rect 498154 408338 498186 408574
rect 498422 408338 498506 408574
rect 498742 408338 498774 408574
rect 498154 390894 498774 408338
rect 498154 390658 498186 390894
rect 498422 390658 498506 390894
rect 498742 390658 498774 390894
rect 498154 390574 498774 390658
rect 498154 390338 498186 390574
rect 498422 390338 498506 390574
rect 498742 390338 498774 390574
rect 498154 372894 498774 390338
rect 498154 372658 498186 372894
rect 498422 372658 498506 372894
rect 498742 372658 498774 372894
rect 498154 372574 498774 372658
rect 498154 372338 498186 372574
rect 498422 372338 498506 372574
rect 498742 372338 498774 372574
rect 498154 354894 498774 372338
rect 498154 354658 498186 354894
rect 498422 354658 498506 354894
rect 498742 354658 498774 354894
rect 498154 354574 498774 354658
rect 498154 354338 498186 354574
rect 498422 354338 498506 354574
rect 498742 354338 498774 354574
rect 498154 336894 498774 354338
rect 498154 336658 498186 336894
rect 498422 336658 498506 336894
rect 498742 336658 498774 336894
rect 498154 336574 498774 336658
rect 498154 336338 498186 336574
rect 498422 336338 498506 336574
rect 498742 336338 498774 336574
rect 498154 318894 498774 336338
rect 498154 318658 498186 318894
rect 498422 318658 498506 318894
rect 498742 318658 498774 318894
rect 498154 318574 498774 318658
rect 498154 318338 498186 318574
rect 498422 318338 498506 318574
rect 498742 318338 498774 318574
rect 498154 300894 498774 318338
rect 498154 300658 498186 300894
rect 498422 300658 498506 300894
rect 498742 300658 498774 300894
rect 498154 300574 498774 300658
rect 498154 300338 498186 300574
rect 498422 300338 498506 300574
rect 498742 300338 498774 300574
rect 498154 282894 498774 300338
rect 498154 282658 498186 282894
rect 498422 282658 498506 282894
rect 498742 282658 498774 282894
rect 498154 282574 498774 282658
rect 498154 282338 498186 282574
rect 498422 282338 498506 282574
rect 498742 282338 498774 282574
rect 498154 264894 498774 282338
rect 498154 264658 498186 264894
rect 498422 264658 498506 264894
rect 498742 264658 498774 264894
rect 498154 264574 498774 264658
rect 498154 264338 498186 264574
rect 498422 264338 498506 264574
rect 498742 264338 498774 264574
rect 498154 246894 498774 264338
rect 498154 246658 498186 246894
rect 498422 246658 498506 246894
rect 498742 246658 498774 246894
rect 498154 246574 498774 246658
rect 498154 246338 498186 246574
rect 498422 246338 498506 246574
rect 498742 246338 498774 246574
rect 498154 228894 498774 246338
rect 498154 228658 498186 228894
rect 498422 228658 498506 228894
rect 498742 228658 498774 228894
rect 498154 228574 498774 228658
rect 498154 228338 498186 228574
rect 498422 228338 498506 228574
rect 498742 228338 498774 228574
rect 498154 210894 498774 228338
rect 498154 210658 498186 210894
rect 498422 210658 498506 210894
rect 498742 210658 498774 210894
rect 498154 210574 498774 210658
rect 498154 210338 498186 210574
rect 498422 210338 498506 210574
rect 498742 210338 498774 210574
rect 498154 192894 498774 210338
rect 498154 192658 498186 192894
rect 498422 192658 498506 192894
rect 498742 192658 498774 192894
rect 498154 192574 498774 192658
rect 498154 192338 498186 192574
rect 498422 192338 498506 192574
rect 498742 192338 498774 192574
rect 498154 174894 498774 192338
rect 498154 174658 498186 174894
rect 498422 174658 498506 174894
rect 498742 174658 498774 174894
rect 498154 174574 498774 174658
rect 498154 174338 498186 174574
rect 498422 174338 498506 174574
rect 498742 174338 498774 174574
rect 498154 156894 498774 174338
rect 498154 156658 498186 156894
rect 498422 156658 498506 156894
rect 498742 156658 498774 156894
rect 498154 156574 498774 156658
rect 498154 156338 498186 156574
rect 498422 156338 498506 156574
rect 498742 156338 498774 156574
rect 498154 138894 498774 156338
rect 498154 138658 498186 138894
rect 498422 138658 498506 138894
rect 498742 138658 498774 138894
rect 498154 138574 498774 138658
rect 498154 138338 498186 138574
rect 498422 138338 498506 138574
rect 498742 138338 498774 138574
rect 498154 120894 498774 138338
rect 498154 120658 498186 120894
rect 498422 120658 498506 120894
rect 498742 120658 498774 120894
rect 498154 120574 498774 120658
rect 498154 120338 498186 120574
rect 498422 120338 498506 120574
rect 498742 120338 498774 120574
rect 498154 102894 498774 120338
rect 498154 102658 498186 102894
rect 498422 102658 498506 102894
rect 498742 102658 498774 102894
rect 498154 102574 498774 102658
rect 498154 102338 498186 102574
rect 498422 102338 498506 102574
rect 498742 102338 498774 102574
rect 498154 84894 498774 102338
rect 498154 84658 498186 84894
rect 498422 84658 498506 84894
rect 498742 84658 498774 84894
rect 498154 84574 498774 84658
rect 498154 84338 498186 84574
rect 498422 84338 498506 84574
rect 498742 84338 498774 84574
rect 498154 66894 498774 84338
rect 498154 66658 498186 66894
rect 498422 66658 498506 66894
rect 498742 66658 498774 66894
rect 498154 66574 498774 66658
rect 498154 66338 498186 66574
rect 498422 66338 498506 66574
rect 498742 66338 498774 66574
rect 498154 48894 498774 66338
rect 498154 48658 498186 48894
rect 498422 48658 498506 48894
rect 498742 48658 498774 48894
rect 498154 48574 498774 48658
rect 498154 48338 498186 48574
rect 498422 48338 498506 48574
rect 498742 48338 498774 48574
rect 498154 30894 498774 48338
rect 498154 30658 498186 30894
rect 498422 30658 498506 30894
rect 498742 30658 498774 30894
rect 498154 30574 498774 30658
rect 498154 30338 498186 30574
rect 498422 30338 498506 30574
rect 498742 30338 498774 30574
rect 498154 12894 498774 30338
rect 498154 12658 498186 12894
rect 498422 12658 498506 12894
rect 498742 12658 498774 12894
rect 498154 12574 498774 12658
rect 498154 12338 498186 12574
rect 498422 12338 498506 12574
rect 498742 12338 498774 12574
rect 498154 -2776 498774 12338
rect 501874 463972 502494 464004
rect 501874 463736 501906 463972
rect 502142 463736 502226 463972
rect 502462 463736 502494 463972
rect 501874 463652 502494 463736
rect 501874 463416 501906 463652
rect 502142 463416 502226 463652
rect 502462 463416 502494 463652
rect 501874 448614 502494 463416
rect 501874 448378 501906 448614
rect 502142 448378 502226 448614
rect 502462 448378 502494 448614
rect 501874 448294 502494 448378
rect 501874 448058 501906 448294
rect 502142 448058 502226 448294
rect 502462 448058 502494 448294
rect 501874 430614 502494 448058
rect 501874 430378 501906 430614
rect 502142 430378 502226 430614
rect 502462 430378 502494 430614
rect 501874 430294 502494 430378
rect 501874 430058 501906 430294
rect 502142 430058 502226 430294
rect 502462 430058 502494 430294
rect 501874 412614 502494 430058
rect 501874 412378 501906 412614
rect 502142 412378 502226 412614
rect 502462 412378 502494 412614
rect 501874 412294 502494 412378
rect 501874 412058 501906 412294
rect 502142 412058 502226 412294
rect 502462 412058 502494 412294
rect 501874 394614 502494 412058
rect 501874 394378 501906 394614
rect 502142 394378 502226 394614
rect 502462 394378 502494 394614
rect 501874 394294 502494 394378
rect 501874 394058 501906 394294
rect 502142 394058 502226 394294
rect 502462 394058 502494 394294
rect 501874 376614 502494 394058
rect 501874 376378 501906 376614
rect 502142 376378 502226 376614
rect 502462 376378 502494 376614
rect 501874 376294 502494 376378
rect 501874 376058 501906 376294
rect 502142 376058 502226 376294
rect 502462 376058 502494 376294
rect 501874 358614 502494 376058
rect 501874 358378 501906 358614
rect 502142 358378 502226 358614
rect 502462 358378 502494 358614
rect 501874 358294 502494 358378
rect 501874 358058 501906 358294
rect 502142 358058 502226 358294
rect 502462 358058 502494 358294
rect 501874 340614 502494 358058
rect 501874 340378 501906 340614
rect 502142 340378 502226 340614
rect 502462 340378 502494 340614
rect 501874 340294 502494 340378
rect 501874 340058 501906 340294
rect 502142 340058 502226 340294
rect 502462 340058 502494 340294
rect 501874 322614 502494 340058
rect 501874 322378 501906 322614
rect 502142 322378 502226 322614
rect 502462 322378 502494 322614
rect 501874 322294 502494 322378
rect 501874 322058 501906 322294
rect 502142 322058 502226 322294
rect 502462 322058 502494 322294
rect 501874 304614 502494 322058
rect 501874 304378 501906 304614
rect 502142 304378 502226 304614
rect 502462 304378 502494 304614
rect 501874 304294 502494 304378
rect 501874 304058 501906 304294
rect 502142 304058 502226 304294
rect 502462 304058 502494 304294
rect 501874 286614 502494 304058
rect 501874 286378 501906 286614
rect 502142 286378 502226 286614
rect 502462 286378 502494 286614
rect 501874 286294 502494 286378
rect 501874 286058 501906 286294
rect 502142 286058 502226 286294
rect 502462 286058 502494 286294
rect 501874 268614 502494 286058
rect 501874 268378 501906 268614
rect 502142 268378 502226 268614
rect 502462 268378 502494 268614
rect 501874 268294 502494 268378
rect 501874 268058 501906 268294
rect 502142 268058 502226 268294
rect 502462 268058 502494 268294
rect 501874 250614 502494 268058
rect 501874 250378 501906 250614
rect 502142 250378 502226 250614
rect 502462 250378 502494 250614
rect 501874 250294 502494 250378
rect 501874 250058 501906 250294
rect 502142 250058 502226 250294
rect 502462 250058 502494 250294
rect 501874 232614 502494 250058
rect 501874 232378 501906 232614
rect 502142 232378 502226 232614
rect 502462 232378 502494 232614
rect 501874 232294 502494 232378
rect 501874 232058 501906 232294
rect 502142 232058 502226 232294
rect 502462 232058 502494 232294
rect 501874 214614 502494 232058
rect 501874 214378 501906 214614
rect 502142 214378 502226 214614
rect 502462 214378 502494 214614
rect 501874 214294 502494 214378
rect 501874 214058 501906 214294
rect 502142 214058 502226 214294
rect 502462 214058 502494 214294
rect 501874 196614 502494 214058
rect 501874 196378 501906 196614
rect 502142 196378 502226 196614
rect 502462 196378 502494 196614
rect 501874 196294 502494 196378
rect 501874 196058 501906 196294
rect 502142 196058 502226 196294
rect 502462 196058 502494 196294
rect 501874 178614 502494 196058
rect 501874 178378 501906 178614
rect 502142 178378 502226 178614
rect 502462 178378 502494 178614
rect 501874 178294 502494 178378
rect 501874 178058 501906 178294
rect 502142 178058 502226 178294
rect 502462 178058 502494 178294
rect 501874 160614 502494 178058
rect 501874 160378 501906 160614
rect 502142 160378 502226 160614
rect 502462 160378 502494 160614
rect 501874 160294 502494 160378
rect 501874 160058 501906 160294
rect 502142 160058 502226 160294
rect 502462 160058 502494 160294
rect 501874 142614 502494 160058
rect 501874 142378 501906 142614
rect 502142 142378 502226 142614
rect 502462 142378 502494 142614
rect 501874 142294 502494 142378
rect 501874 142058 501906 142294
rect 502142 142058 502226 142294
rect 502462 142058 502494 142294
rect 501874 124614 502494 142058
rect 501874 124378 501906 124614
rect 502142 124378 502226 124614
rect 502462 124378 502494 124614
rect 501874 124294 502494 124378
rect 501874 124058 501906 124294
rect 502142 124058 502226 124294
rect 502462 124058 502494 124294
rect 501874 106614 502494 124058
rect 501874 106378 501906 106614
rect 502142 106378 502226 106614
rect 502462 106378 502494 106614
rect 501874 106294 502494 106378
rect 501874 106058 501906 106294
rect 502142 106058 502226 106294
rect 502462 106058 502494 106294
rect 501874 88614 502494 106058
rect 501874 88378 501906 88614
rect 502142 88378 502226 88614
rect 502462 88378 502494 88614
rect 501874 88294 502494 88378
rect 501874 88058 501906 88294
rect 502142 88058 502226 88294
rect 502462 88058 502494 88294
rect 501874 70614 502494 88058
rect 501874 70378 501906 70614
rect 502142 70378 502226 70614
rect 502462 70378 502494 70614
rect 501874 70294 502494 70378
rect 501874 70058 501906 70294
rect 502142 70058 502226 70294
rect 502462 70058 502494 70294
rect 501874 52614 502494 70058
rect 501874 52378 501906 52614
rect 502142 52378 502226 52614
rect 502462 52378 502494 52614
rect 501874 52294 502494 52378
rect 501874 52058 501906 52294
rect 502142 52058 502226 52294
rect 502462 52058 502494 52294
rect 501874 34614 502494 52058
rect 501874 34378 501906 34614
rect 502142 34378 502226 34614
rect 502462 34378 502494 34614
rect 501874 34294 502494 34378
rect 501874 34058 501906 34294
rect 502142 34058 502226 34294
rect 502462 34058 502494 34294
rect 501874 16614 502494 34058
rect 501874 16378 501906 16614
rect 502142 16378 502226 16614
rect 502462 16378 502494 16614
rect 501874 16294 502494 16378
rect 501874 16058 501906 16294
rect 502142 16058 502226 16294
rect 502462 16058 502494 16294
rect 501874 880 502494 16058
rect 508714 461092 509334 464004
rect 508714 460856 508746 461092
rect 508982 460856 509066 461092
rect 509302 460856 509334 461092
rect 508714 460772 509334 460856
rect 508714 460536 508746 460772
rect 508982 460536 509066 460772
rect 509302 460536 509334 460772
rect 508714 455454 509334 460536
rect 508714 455218 508746 455454
rect 508982 455218 509066 455454
rect 509302 455218 509334 455454
rect 508714 455134 509334 455218
rect 508714 454898 508746 455134
rect 508982 454898 509066 455134
rect 509302 454898 509334 455134
rect 508714 437454 509334 454898
rect 508714 437218 508746 437454
rect 508982 437218 509066 437454
rect 509302 437218 509334 437454
rect 508714 437134 509334 437218
rect 508714 436898 508746 437134
rect 508982 436898 509066 437134
rect 509302 436898 509334 437134
rect 508714 419454 509334 436898
rect 508714 419218 508746 419454
rect 508982 419218 509066 419454
rect 509302 419218 509334 419454
rect 508714 419134 509334 419218
rect 508714 418898 508746 419134
rect 508982 418898 509066 419134
rect 509302 418898 509334 419134
rect 508714 401454 509334 418898
rect 508714 401218 508746 401454
rect 508982 401218 509066 401454
rect 509302 401218 509334 401454
rect 508714 401134 509334 401218
rect 508714 400898 508746 401134
rect 508982 400898 509066 401134
rect 509302 400898 509334 401134
rect 508714 383454 509334 400898
rect 508714 383218 508746 383454
rect 508982 383218 509066 383454
rect 509302 383218 509334 383454
rect 508714 383134 509334 383218
rect 508714 382898 508746 383134
rect 508982 382898 509066 383134
rect 509302 382898 509334 383134
rect 508714 365454 509334 382898
rect 508714 365218 508746 365454
rect 508982 365218 509066 365454
rect 509302 365218 509334 365454
rect 508714 365134 509334 365218
rect 508714 364898 508746 365134
rect 508982 364898 509066 365134
rect 509302 364898 509334 365134
rect 508714 347454 509334 364898
rect 508714 347218 508746 347454
rect 508982 347218 509066 347454
rect 509302 347218 509334 347454
rect 508714 347134 509334 347218
rect 508714 346898 508746 347134
rect 508982 346898 509066 347134
rect 509302 346898 509334 347134
rect 508714 329454 509334 346898
rect 508714 329218 508746 329454
rect 508982 329218 509066 329454
rect 509302 329218 509334 329454
rect 508714 329134 509334 329218
rect 508714 328898 508746 329134
rect 508982 328898 509066 329134
rect 509302 328898 509334 329134
rect 508714 311454 509334 328898
rect 508714 311218 508746 311454
rect 508982 311218 509066 311454
rect 509302 311218 509334 311454
rect 508714 311134 509334 311218
rect 508714 310898 508746 311134
rect 508982 310898 509066 311134
rect 509302 310898 509334 311134
rect 508714 293454 509334 310898
rect 508714 293218 508746 293454
rect 508982 293218 509066 293454
rect 509302 293218 509334 293454
rect 508714 293134 509334 293218
rect 508714 292898 508746 293134
rect 508982 292898 509066 293134
rect 509302 292898 509334 293134
rect 508714 275454 509334 292898
rect 508714 275218 508746 275454
rect 508982 275218 509066 275454
rect 509302 275218 509334 275454
rect 508714 275134 509334 275218
rect 508714 274898 508746 275134
rect 508982 274898 509066 275134
rect 509302 274898 509334 275134
rect 508714 257454 509334 274898
rect 508714 257218 508746 257454
rect 508982 257218 509066 257454
rect 509302 257218 509334 257454
rect 508714 257134 509334 257218
rect 508714 256898 508746 257134
rect 508982 256898 509066 257134
rect 509302 256898 509334 257134
rect 508714 239454 509334 256898
rect 508714 239218 508746 239454
rect 508982 239218 509066 239454
rect 509302 239218 509334 239454
rect 508714 239134 509334 239218
rect 508714 238898 508746 239134
rect 508982 238898 509066 239134
rect 509302 238898 509334 239134
rect 508714 221454 509334 238898
rect 508714 221218 508746 221454
rect 508982 221218 509066 221454
rect 509302 221218 509334 221454
rect 508714 221134 509334 221218
rect 508714 220898 508746 221134
rect 508982 220898 509066 221134
rect 509302 220898 509334 221134
rect 508714 203454 509334 220898
rect 508714 203218 508746 203454
rect 508982 203218 509066 203454
rect 509302 203218 509334 203454
rect 508714 203134 509334 203218
rect 508714 202898 508746 203134
rect 508982 202898 509066 203134
rect 509302 202898 509334 203134
rect 508714 185454 509334 202898
rect 508714 185218 508746 185454
rect 508982 185218 509066 185454
rect 509302 185218 509334 185454
rect 508714 185134 509334 185218
rect 508714 184898 508746 185134
rect 508982 184898 509066 185134
rect 509302 184898 509334 185134
rect 508714 167454 509334 184898
rect 508714 167218 508746 167454
rect 508982 167218 509066 167454
rect 509302 167218 509334 167454
rect 508714 167134 509334 167218
rect 508714 166898 508746 167134
rect 508982 166898 509066 167134
rect 509302 166898 509334 167134
rect 508714 149454 509334 166898
rect 508714 149218 508746 149454
rect 508982 149218 509066 149454
rect 509302 149218 509334 149454
rect 508714 149134 509334 149218
rect 508714 148898 508746 149134
rect 508982 148898 509066 149134
rect 509302 148898 509334 149134
rect 508714 131454 509334 148898
rect 508714 131218 508746 131454
rect 508982 131218 509066 131454
rect 509302 131218 509334 131454
rect 508714 131134 509334 131218
rect 508714 130898 508746 131134
rect 508982 130898 509066 131134
rect 509302 130898 509334 131134
rect 508714 113454 509334 130898
rect 508714 113218 508746 113454
rect 508982 113218 509066 113454
rect 509302 113218 509334 113454
rect 508714 113134 509334 113218
rect 508714 112898 508746 113134
rect 508982 112898 509066 113134
rect 509302 112898 509334 113134
rect 508714 95454 509334 112898
rect 508714 95218 508746 95454
rect 508982 95218 509066 95454
rect 509302 95218 509334 95454
rect 508714 95134 509334 95218
rect 508714 94898 508746 95134
rect 508982 94898 509066 95134
rect 509302 94898 509334 95134
rect 508714 77454 509334 94898
rect 508714 77218 508746 77454
rect 508982 77218 509066 77454
rect 509302 77218 509334 77454
rect 508714 77134 509334 77218
rect 508714 76898 508746 77134
rect 508982 76898 509066 77134
rect 509302 76898 509334 77134
rect 508714 59454 509334 76898
rect 508714 59218 508746 59454
rect 508982 59218 509066 59454
rect 509302 59218 509334 59454
rect 508714 59134 509334 59218
rect 508714 58898 508746 59134
rect 508982 58898 509066 59134
rect 509302 58898 509334 59134
rect 508714 41454 509334 58898
rect 508714 41218 508746 41454
rect 508982 41218 509066 41454
rect 509302 41218 509334 41454
rect 508714 41134 509334 41218
rect 508714 40898 508746 41134
rect 508982 40898 509066 41134
rect 509302 40898 509334 41134
rect 508714 23454 509334 40898
rect 508714 23218 508746 23454
rect 508982 23218 509066 23454
rect 509302 23218 509334 23454
rect 508714 23134 509334 23218
rect 508714 22898 508746 23134
rect 508982 22898 509066 23134
rect 509302 22898 509334 23134
rect 508714 5454 509334 22898
rect 508714 5218 508746 5454
rect 508982 5218 509066 5454
rect 509302 5218 509334 5454
rect 508714 5134 509334 5218
rect 508714 4898 508746 5134
rect 508982 4898 509066 5134
rect 509302 4898 509334 5134
rect 508714 880 509334 4898
rect 512434 462052 513054 464004
rect 512434 461816 512466 462052
rect 512702 461816 512786 462052
rect 513022 461816 513054 462052
rect 512434 461732 513054 461816
rect 512434 461496 512466 461732
rect 512702 461496 512786 461732
rect 513022 461496 513054 461732
rect 512434 441174 513054 461496
rect 512434 440938 512466 441174
rect 512702 440938 512786 441174
rect 513022 440938 513054 441174
rect 512434 440854 513054 440938
rect 512434 440618 512466 440854
rect 512702 440618 512786 440854
rect 513022 440618 513054 440854
rect 512434 423174 513054 440618
rect 512434 422938 512466 423174
rect 512702 422938 512786 423174
rect 513022 422938 513054 423174
rect 512434 422854 513054 422938
rect 512434 422618 512466 422854
rect 512702 422618 512786 422854
rect 513022 422618 513054 422854
rect 512434 405174 513054 422618
rect 512434 404938 512466 405174
rect 512702 404938 512786 405174
rect 513022 404938 513054 405174
rect 512434 404854 513054 404938
rect 512434 404618 512466 404854
rect 512702 404618 512786 404854
rect 513022 404618 513054 404854
rect 512434 387174 513054 404618
rect 512434 386938 512466 387174
rect 512702 386938 512786 387174
rect 513022 386938 513054 387174
rect 512434 386854 513054 386938
rect 512434 386618 512466 386854
rect 512702 386618 512786 386854
rect 513022 386618 513054 386854
rect 512434 369174 513054 386618
rect 512434 368938 512466 369174
rect 512702 368938 512786 369174
rect 513022 368938 513054 369174
rect 512434 368854 513054 368938
rect 512434 368618 512466 368854
rect 512702 368618 512786 368854
rect 513022 368618 513054 368854
rect 512434 351174 513054 368618
rect 512434 350938 512466 351174
rect 512702 350938 512786 351174
rect 513022 350938 513054 351174
rect 512434 350854 513054 350938
rect 512434 350618 512466 350854
rect 512702 350618 512786 350854
rect 513022 350618 513054 350854
rect 512434 333174 513054 350618
rect 512434 332938 512466 333174
rect 512702 332938 512786 333174
rect 513022 332938 513054 333174
rect 512434 332854 513054 332938
rect 512434 332618 512466 332854
rect 512702 332618 512786 332854
rect 513022 332618 513054 332854
rect 512434 315174 513054 332618
rect 512434 314938 512466 315174
rect 512702 314938 512786 315174
rect 513022 314938 513054 315174
rect 512434 314854 513054 314938
rect 512434 314618 512466 314854
rect 512702 314618 512786 314854
rect 513022 314618 513054 314854
rect 512434 297174 513054 314618
rect 512434 296938 512466 297174
rect 512702 296938 512786 297174
rect 513022 296938 513054 297174
rect 512434 296854 513054 296938
rect 512434 296618 512466 296854
rect 512702 296618 512786 296854
rect 513022 296618 513054 296854
rect 512434 279174 513054 296618
rect 512434 278938 512466 279174
rect 512702 278938 512786 279174
rect 513022 278938 513054 279174
rect 512434 278854 513054 278938
rect 512434 278618 512466 278854
rect 512702 278618 512786 278854
rect 513022 278618 513054 278854
rect 512434 261174 513054 278618
rect 512434 260938 512466 261174
rect 512702 260938 512786 261174
rect 513022 260938 513054 261174
rect 512434 260854 513054 260938
rect 512434 260618 512466 260854
rect 512702 260618 512786 260854
rect 513022 260618 513054 260854
rect 512434 243174 513054 260618
rect 512434 242938 512466 243174
rect 512702 242938 512786 243174
rect 513022 242938 513054 243174
rect 512434 242854 513054 242938
rect 512434 242618 512466 242854
rect 512702 242618 512786 242854
rect 513022 242618 513054 242854
rect 512434 225174 513054 242618
rect 512434 224938 512466 225174
rect 512702 224938 512786 225174
rect 513022 224938 513054 225174
rect 512434 224854 513054 224938
rect 512434 224618 512466 224854
rect 512702 224618 512786 224854
rect 513022 224618 513054 224854
rect 512434 207174 513054 224618
rect 512434 206938 512466 207174
rect 512702 206938 512786 207174
rect 513022 206938 513054 207174
rect 512434 206854 513054 206938
rect 512434 206618 512466 206854
rect 512702 206618 512786 206854
rect 513022 206618 513054 206854
rect 512434 189174 513054 206618
rect 512434 188938 512466 189174
rect 512702 188938 512786 189174
rect 513022 188938 513054 189174
rect 512434 188854 513054 188938
rect 512434 188618 512466 188854
rect 512702 188618 512786 188854
rect 513022 188618 513054 188854
rect 512434 171174 513054 188618
rect 512434 170938 512466 171174
rect 512702 170938 512786 171174
rect 513022 170938 513054 171174
rect 512434 170854 513054 170938
rect 512434 170618 512466 170854
rect 512702 170618 512786 170854
rect 513022 170618 513054 170854
rect 512434 153174 513054 170618
rect 512434 152938 512466 153174
rect 512702 152938 512786 153174
rect 513022 152938 513054 153174
rect 512434 152854 513054 152938
rect 512434 152618 512466 152854
rect 512702 152618 512786 152854
rect 513022 152618 513054 152854
rect 512434 135174 513054 152618
rect 512434 134938 512466 135174
rect 512702 134938 512786 135174
rect 513022 134938 513054 135174
rect 512434 134854 513054 134938
rect 512434 134618 512466 134854
rect 512702 134618 512786 134854
rect 513022 134618 513054 134854
rect 512434 117174 513054 134618
rect 512434 116938 512466 117174
rect 512702 116938 512786 117174
rect 513022 116938 513054 117174
rect 512434 116854 513054 116938
rect 512434 116618 512466 116854
rect 512702 116618 512786 116854
rect 513022 116618 513054 116854
rect 512434 99174 513054 116618
rect 512434 98938 512466 99174
rect 512702 98938 512786 99174
rect 513022 98938 513054 99174
rect 512434 98854 513054 98938
rect 512434 98618 512466 98854
rect 512702 98618 512786 98854
rect 513022 98618 513054 98854
rect 512434 81174 513054 98618
rect 512434 80938 512466 81174
rect 512702 80938 512786 81174
rect 513022 80938 513054 81174
rect 512434 80854 513054 80938
rect 512434 80618 512466 80854
rect 512702 80618 512786 80854
rect 513022 80618 513054 80854
rect 512434 63174 513054 80618
rect 512434 62938 512466 63174
rect 512702 62938 512786 63174
rect 513022 62938 513054 63174
rect 512434 62854 513054 62938
rect 512434 62618 512466 62854
rect 512702 62618 512786 62854
rect 513022 62618 513054 62854
rect 512434 45174 513054 62618
rect 512434 44938 512466 45174
rect 512702 44938 512786 45174
rect 513022 44938 513054 45174
rect 512434 44854 513054 44938
rect 512434 44618 512466 44854
rect 512702 44618 512786 44854
rect 513022 44618 513054 44854
rect 512434 27174 513054 44618
rect 512434 26938 512466 27174
rect 512702 26938 512786 27174
rect 513022 26938 513054 27174
rect 512434 26854 513054 26938
rect 512434 26618 512466 26854
rect 512702 26618 512786 26854
rect 513022 26618 513054 26854
rect 512434 9174 513054 26618
rect 512434 8938 512466 9174
rect 512702 8938 512786 9174
rect 513022 8938 513054 9174
rect 512434 8854 513054 8938
rect 512434 8618 512466 8854
rect 512702 8618 512786 8854
rect 513022 8618 513054 8854
rect 512434 880 513054 8618
rect 516154 463012 516774 464004
rect 516154 462776 516186 463012
rect 516422 462776 516506 463012
rect 516742 462776 516774 463012
rect 516154 462692 516774 462776
rect 516154 462456 516186 462692
rect 516422 462456 516506 462692
rect 516742 462456 516774 462692
rect 516154 444894 516774 462456
rect 516154 444658 516186 444894
rect 516422 444658 516506 444894
rect 516742 444658 516774 444894
rect 516154 444574 516774 444658
rect 516154 444338 516186 444574
rect 516422 444338 516506 444574
rect 516742 444338 516774 444574
rect 516154 426894 516774 444338
rect 516154 426658 516186 426894
rect 516422 426658 516506 426894
rect 516742 426658 516774 426894
rect 516154 426574 516774 426658
rect 516154 426338 516186 426574
rect 516422 426338 516506 426574
rect 516742 426338 516774 426574
rect 516154 408894 516774 426338
rect 516154 408658 516186 408894
rect 516422 408658 516506 408894
rect 516742 408658 516774 408894
rect 516154 408574 516774 408658
rect 516154 408338 516186 408574
rect 516422 408338 516506 408574
rect 516742 408338 516774 408574
rect 516154 390894 516774 408338
rect 516154 390658 516186 390894
rect 516422 390658 516506 390894
rect 516742 390658 516774 390894
rect 516154 390574 516774 390658
rect 516154 390338 516186 390574
rect 516422 390338 516506 390574
rect 516742 390338 516774 390574
rect 516154 372894 516774 390338
rect 516154 372658 516186 372894
rect 516422 372658 516506 372894
rect 516742 372658 516774 372894
rect 516154 372574 516774 372658
rect 516154 372338 516186 372574
rect 516422 372338 516506 372574
rect 516742 372338 516774 372574
rect 516154 354894 516774 372338
rect 516154 354658 516186 354894
rect 516422 354658 516506 354894
rect 516742 354658 516774 354894
rect 516154 354574 516774 354658
rect 516154 354338 516186 354574
rect 516422 354338 516506 354574
rect 516742 354338 516774 354574
rect 516154 336894 516774 354338
rect 516154 336658 516186 336894
rect 516422 336658 516506 336894
rect 516742 336658 516774 336894
rect 516154 336574 516774 336658
rect 516154 336338 516186 336574
rect 516422 336338 516506 336574
rect 516742 336338 516774 336574
rect 516154 318894 516774 336338
rect 516154 318658 516186 318894
rect 516422 318658 516506 318894
rect 516742 318658 516774 318894
rect 516154 318574 516774 318658
rect 516154 318338 516186 318574
rect 516422 318338 516506 318574
rect 516742 318338 516774 318574
rect 516154 300894 516774 318338
rect 516154 300658 516186 300894
rect 516422 300658 516506 300894
rect 516742 300658 516774 300894
rect 516154 300574 516774 300658
rect 516154 300338 516186 300574
rect 516422 300338 516506 300574
rect 516742 300338 516774 300574
rect 516154 282894 516774 300338
rect 516154 282658 516186 282894
rect 516422 282658 516506 282894
rect 516742 282658 516774 282894
rect 516154 282574 516774 282658
rect 516154 282338 516186 282574
rect 516422 282338 516506 282574
rect 516742 282338 516774 282574
rect 516154 264894 516774 282338
rect 516154 264658 516186 264894
rect 516422 264658 516506 264894
rect 516742 264658 516774 264894
rect 516154 264574 516774 264658
rect 516154 264338 516186 264574
rect 516422 264338 516506 264574
rect 516742 264338 516774 264574
rect 516154 246894 516774 264338
rect 516154 246658 516186 246894
rect 516422 246658 516506 246894
rect 516742 246658 516774 246894
rect 516154 246574 516774 246658
rect 516154 246338 516186 246574
rect 516422 246338 516506 246574
rect 516742 246338 516774 246574
rect 516154 228894 516774 246338
rect 516154 228658 516186 228894
rect 516422 228658 516506 228894
rect 516742 228658 516774 228894
rect 516154 228574 516774 228658
rect 516154 228338 516186 228574
rect 516422 228338 516506 228574
rect 516742 228338 516774 228574
rect 516154 210894 516774 228338
rect 516154 210658 516186 210894
rect 516422 210658 516506 210894
rect 516742 210658 516774 210894
rect 516154 210574 516774 210658
rect 516154 210338 516186 210574
rect 516422 210338 516506 210574
rect 516742 210338 516774 210574
rect 516154 192894 516774 210338
rect 516154 192658 516186 192894
rect 516422 192658 516506 192894
rect 516742 192658 516774 192894
rect 516154 192574 516774 192658
rect 516154 192338 516186 192574
rect 516422 192338 516506 192574
rect 516742 192338 516774 192574
rect 516154 174894 516774 192338
rect 516154 174658 516186 174894
rect 516422 174658 516506 174894
rect 516742 174658 516774 174894
rect 516154 174574 516774 174658
rect 516154 174338 516186 174574
rect 516422 174338 516506 174574
rect 516742 174338 516774 174574
rect 516154 156894 516774 174338
rect 516154 156658 516186 156894
rect 516422 156658 516506 156894
rect 516742 156658 516774 156894
rect 516154 156574 516774 156658
rect 516154 156338 516186 156574
rect 516422 156338 516506 156574
rect 516742 156338 516774 156574
rect 516154 138894 516774 156338
rect 516154 138658 516186 138894
rect 516422 138658 516506 138894
rect 516742 138658 516774 138894
rect 516154 138574 516774 138658
rect 516154 138338 516186 138574
rect 516422 138338 516506 138574
rect 516742 138338 516774 138574
rect 516154 120894 516774 138338
rect 516154 120658 516186 120894
rect 516422 120658 516506 120894
rect 516742 120658 516774 120894
rect 516154 120574 516774 120658
rect 516154 120338 516186 120574
rect 516422 120338 516506 120574
rect 516742 120338 516774 120574
rect 516154 102894 516774 120338
rect 516154 102658 516186 102894
rect 516422 102658 516506 102894
rect 516742 102658 516774 102894
rect 516154 102574 516774 102658
rect 516154 102338 516186 102574
rect 516422 102338 516506 102574
rect 516742 102338 516774 102574
rect 516154 84894 516774 102338
rect 516154 84658 516186 84894
rect 516422 84658 516506 84894
rect 516742 84658 516774 84894
rect 516154 84574 516774 84658
rect 516154 84338 516186 84574
rect 516422 84338 516506 84574
rect 516742 84338 516774 84574
rect 516154 66894 516774 84338
rect 516154 66658 516186 66894
rect 516422 66658 516506 66894
rect 516742 66658 516774 66894
rect 516154 66574 516774 66658
rect 516154 66338 516186 66574
rect 516422 66338 516506 66574
rect 516742 66338 516774 66574
rect 516154 48894 516774 66338
rect 516154 48658 516186 48894
rect 516422 48658 516506 48894
rect 516742 48658 516774 48894
rect 516154 48574 516774 48658
rect 516154 48338 516186 48574
rect 516422 48338 516506 48574
rect 516742 48338 516774 48574
rect 516154 30894 516774 48338
rect 516154 30658 516186 30894
rect 516422 30658 516506 30894
rect 516742 30658 516774 30894
rect 516154 30574 516774 30658
rect 516154 30338 516186 30574
rect 516422 30338 516506 30574
rect 516742 30338 516774 30574
rect 516154 12894 516774 30338
rect 516154 12658 516186 12894
rect 516422 12658 516506 12894
rect 516742 12658 516774 12894
rect 516154 12574 516774 12658
rect 516154 12338 516186 12574
rect 516422 12338 516506 12574
rect 516742 12338 516774 12574
rect 516154 880 516774 12338
rect 519874 463972 520494 464004
rect 519874 463736 519906 463972
rect 520142 463736 520226 463972
rect 520462 463736 520494 463972
rect 519874 463652 520494 463736
rect 519874 463416 519906 463652
rect 520142 463416 520226 463652
rect 520462 463416 520494 463652
rect 519874 448614 520494 463416
rect 519874 448378 519906 448614
rect 520142 448378 520226 448614
rect 520462 448378 520494 448614
rect 519874 448294 520494 448378
rect 519874 448058 519906 448294
rect 520142 448058 520226 448294
rect 520462 448058 520494 448294
rect 519874 430614 520494 448058
rect 519874 430378 519906 430614
rect 520142 430378 520226 430614
rect 520462 430378 520494 430614
rect 519874 430294 520494 430378
rect 519874 430058 519906 430294
rect 520142 430058 520226 430294
rect 520462 430058 520494 430294
rect 519874 412614 520494 430058
rect 519874 412378 519906 412614
rect 520142 412378 520226 412614
rect 520462 412378 520494 412614
rect 519874 412294 520494 412378
rect 519874 412058 519906 412294
rect 520142 412058 520226 412294
rect 520462 412058 520494 412294
rect 519874 394614 520494 412058
rect 519874 394378 519906 394614
rect 520142 394378 520226 394614
rect 520462 394378 520494 394614
rect 519874 394294 520494 394378
rect 519874 394058 519906 394294
rect 520142 394058 520226 394294
rect 520462 394058 520494 394294
rect 519874 376614 520494 394058
rect 519874 376378 519906 376614
rect 520142 376378 520226 376614
rect 520462 376378 520494 376614
rect 519874 376294 520494 376378
rect 519874 376058 519906 376294
rect 520142 376058 520226 376294
rect 520462 376058 520494 376294
rect 519874 358614 520494 376058
rect 519874 358378 519906 358614
rect 520142 358378 520226 358614
rect 520462 358378 520494 358614
rect 519874 358294 520494 358378
rect 519874 358058 519906 358294
rect 520142 358058 520226 358294
rect 520462 358058 520494 358294
rect 519874 340614 520494 358058
rect 519874 340378 519906 340614
rect 520142 340378 520226 340614
rect 520462 340378 520494 340614
rect 519874 340294 520494 340378
rect 519874 340058 519906 340294
rect 520142 340058 520226 340294
rect 520462 340058 520494 340294
rect 519874 322614 520494 340058
rect 519874 322378 519906 322614
rect 520142 322378 520226 322614
rect 520462 322378 520494 322614
rect 519874 322294 520494 322378
rect 519874 322058 519906 322294
rect 520142 322058 520226 322294
rect 520462 322058 520494 322294
rect 519874 304614 520494 322058
rect 519874 304378 519906 304614
rect 520142 304378 520226 304614
rect 520462 304378 520494 304614
rect 519874 304294 520494 304378
rect 519874 304058 519906 304294
rect 520142 304058 520226 304294
rect 520462 304058 520494 304294
rect 519874 286614 520494 304058
rect 519874 286378 519906 286614
rect 520142 286378 520226 286614
rect 520462 286378 520494 286614
rect 519874 286294 520494 286378
rect 519874 286058 519906 286294
rect 520142 286058 520226 286294
rect 520462 286058 520494 286294
rect 519874 268614 520494 286058
rect 519874 268378 519906 268614
rect 520142 268378 520226 268614
rect 520462 268378 520494 268614
rect 519874 268294 520494 268378
rect 519874 268058 519906 268294
rect 520142 268058 520226 268294
rect 520462 268058 520494 268294
rect 519874 250614 520494 268058
rect 519874 250378 519906 250614
rect 520142 250378 520226 250614
rect 520462 250378 520494 250614
rect 519874 250294 520494 250378
rect 519874 250058 519906 250294
rect 520142 250058 520226 250294
rect 520462 250058 520494 250294
rect 519874 232614 520494 250058
rect 519874 232378 519906 232614
rect 520142 232378 520226 232614
rect 520462 232378 520494 232614
rect 519874 232294 520494 232378
rect 519874 232058 519906 232294
rect 520142 232058 520226 232294
rect 520462 232058 520494 232294
rect 519874 214614 520494 232058
rect 519874 214378 519906 214614
rect 520142 214378 520226 214614
rect 520462 214378 520494 214614
rect 519874 214294 520494 214378
rect 519874 214058 519906 214294
rect 520142 214058 520226 214294
rect 520462 214058 520494 214294
rect 519874 196614 520494 214058
rect 519874 196378 519906 196614
rect 520142 196378 520226 196614
rect 520462 196378 520494 196614
rect 519874 196294 520494 196378
rect 519874 196058 519906 196294
rect 520142 196058 520226 196294
rect 520462 196058 520494 196294
rect 519874 178614 520494 196058
rect 519874 178378 519906 178614
rect 520142 178378 520226 178614
rect 520462 178378 520494 178614
rect 519874 178294 520494 178378
rect 519874 178058 519906 178294
rect 520142 178058 520226 178294
rect 520462 178058 520494 178294
rect 519874 160614 520494 178058
rect 519874 160378 519906 160614
rect 520142 160378 520226 160614
rect 520462 160378 520494 160614
rect 519874 160294 520494 160378
rect 519874 160058 519906 160294
rect 520142 160058 520226 160294
rect 520462 160058 520494 160294
rect 519874 142614 520494 160058
rect 519874 142378 519906 142614
rect 520142 142378 520226 142614
rect 520462 142378 520494 142614
rect 519874 142294 520494 142378
rect 519874 142058 519906 142294
rect 520142 142058 520226 142294
rect 520462 142058 520494 142294
rect 519874 124614 520494 142058
rect 519874 124378 519906 124614
rect 520142 124378 520226 124614
rect 520462 124378 520494 124614
rect 519874 124294 520494 124378
rect 519874 124058 519906 124294
rect 520142 124058 520226 124294
rect 520462 124058 520494 124294
rect 519874 106614 520494 124058
rect 519874 106378 519906 106614
rect 520142 106378 520226 106614
rect 520462 106378 520494 106614
rect 519874 106294 520494 106378
rect 519874 106058 519906 106294
rect 520142 106058 520226 106294
rect 520462 106058 520494 106294
rect 519874 88614 520494 106058
rect 519874 88378 519906 88614
rect 520142 88378 520226 88614
rect 520462 88378 520494 88614
rect 519874 88294 520494 88378
rect 519874 88058 519906 88294
rect 520142 88058 520226 88294
rect 520462 88058 520494 88294
rect 519874 70614 520494 88058
rect 519874 70378 519906 70614
rect 520142 70378 520226 70614
rect 520462 70378 520494 70614
rect 519874 70294 520494 70378
rect 519874 70058 519906 70294
rect 520142 70058 520226 70294
rect 520462 70058 520494 70294
rect 519874 52614 520494 70058
rect 519874 52378 519906 52614
rect 520142 52378 520226 52614
rect 520462 52378 520494 52614
rect 519874 52294 520494 52378
rect 519874 52058 519906 52294
rect 520142 52058 520226 52294
rect 520462 52058 520494 52294
rect 519874 34614 520494 52058
rect 519874 34378 519906 34614
rect 520142 34378 520226 34614
rect 520462 34378 520494 34614
rect 519874 34294 520494 34378
rect 519874 34058 519906 34294
rect 520142 34058 520226 34294
rect 520462 34058 520494 34294
rect 519874 16614 520494 34058
rect 519874 16378 519906 16614
rect 520142 16378 520226 16614
rect 520462 16378 520494 16614
rect 519874 16294 520494 16378
rect 519874 16058 519906 16294
rect 520142 16058 520226 16294
rect 520462 16058 520494 16294
rect 519874 880 520494 16058
rect 526714 461092 527334 464004
rect 526714 460856 526746 461092
rect 526982 460856 527066 461092
rect 527302 460856 527334 461092
rect 526714 460772 527334 460856
rect 526714 460536 526746 460772
rect 526982 460536 527066 460772
rect 527302 460536 527334 460772
rect 526714 455454 527334 460536
rect 526714 455218 526746 455454
rect 526982 455218 527066 455454
rect 527302 455218 527334 455454
rect 526714 455134 527334 455218
rect 526714 454898 526746 455134
rect 526982 454898 527066 455134
rect 527302 454898 527334 455134
rect 526714 437454 527334 454898
rect 526714 437218 526746 437454
rect 526982 437218 527066 437454
rect 527302 437218 527334 437454
rect 526714 437134 527334 437218
rect 526714 436898 526746 437134
rect 526982 436898 527066 437134
rect 527302 436898 527334 437134
rect 526714 419454 527334 436898
rect 526714 419218 526746 419454
rect 526982 419218 527066 419454
rect 527302 419218 527334 419454
rect 526714 419134 527334 419218
rect 526714 418898 526746 419134
rect 526982 418898 527066 419134
rect 527302 418898 527334 419134
rect 526714 401454 527334 418898
rect 526714 401218 526746 401454
rect 526982 401218 527066 401454
rect 527302 401218 527334 401454
rect 526714 401134 527334 401218
rect 526714 400898 526746 401134
rect 526982 400898 527066 401134
rect 527302 400898 527334 401134
rect 526714 383454 527334 400898
rect 526714 383218 526746 383454
rect 526982 383218 527066 383454
rect 527302 383218 527334 383454
rect 526714 383134 527334 383218
rect 526714 382898 526746 383134
rect 526982 382898 527066 383134
rect 527302 382898 527334 383134
rect 526714 365454 527334 382898
rect 526714 365218 526746 365454
rect 526982 365218 527066 365454
rect 527302 365218 527334 365454
rect 526714 365134 527334 365218
rect 526714 364898 526746 365134
rect 526982 364898 527066 365134
rect 527302 364898 527334 365134
rect 526714 347454 527334 364898
rect 526714 347218 526746 347454
rect 526982 347218 527066 347454
rect 527302 347218 527334 347454
rect 526714 347134 527334 347218
rect 526714 346898 526746 347134
rect 526982 346898 527066 347134
rect 527302 346898 527334 347134
rect 526714 329454 527334 346898
rect 526714 329218 526746 329454
rect 526982 329218 527066 329454
rect 527302 329218 527334 329454
rect 526714 329134 527334 329218
rect 526714 328898 526746 329134
rect 526982 328898 527066 329134
rect 527302 328898 527334 329134
rect 526714 311454 527334 328898
rect 526714 311218 526746 311454
rect 526982 311218 527066 311454
rect 527302 311218 527334 311454
rect 526714 311134 527334 311218
rect 526714 310898 526746 311134
rect 526982 310898 527066 311134
rect 527302 310898 527334 311134
rect 526714 293454 527334 310898
rect 526714 293218 526746 293454
rect 526982 293218 527066 293454
rect 527302 293218 527334 293454
rect 526714 293134 527334 293218
rect 526714 292898 526746 293134
rect 526982 292898 527066 293134
rect 527302 292898 527334 293134
rect 526714 275454 527334 292898
rect 526714 275218 526746 275454
rect 526982 275218 527066 275454
rect 527302 275218 527334 275454
rect 526714 275134 527334 275218
rect 526714 274898 526746 275134
rect 526982 274898 527066 275134
rect 527302 274898 527334 275134
rect 526714 257454 527334 274898
rect 526714 257218 526746 257454
rect 526982 257218 527066 257454
rect 527302 257218 527334 257454
rect 526714 257134 527334 257218
rect 526714 256898 526746 257134
rect 526982 256898 527066 257134
rect 527302 256898 527334 257134
rect 526714 239454 527334 256898
rect 526714 239218 526746 239454
rect 526982 239218 527066 239454
rect 527302 239218 527334 239454
rect 526714 239134 527334 239218
rect 526714 238898 526746 239134
rect 526982 238898 527066 239134
rect 527302 238898 527334 239134
rect 526714 221454 527334 238898
rect 526714 221218 526746 221454
rect 526982 221218 527066 221454
rect 527302 221218 527334 221454
rect 526714 221134 527334 221218
rect 526714 220898 526746 221134
rect 526982 220898 527066 221134
rect 527302 220898 527334 221134
rect 526714 203454 527334 220898
rect 526714 203218 526746 203454
rect 526982 203218 527066 203454
rect 527302 203218 527334 203454
rect 526714 203134 527334 203218
rect 526714 202898 526746 203134
rect 526982 202898 527066 203134
rect 527302 202898 527334 203134
rect 526714 185454 527334 202898
rect 526714 185218 526746 185454
rect 526982 185218 527066 185454
rect 527302 185218 527334 185454
rect 526714 185134 527334 185218
rect 526714 184898 526746 185134
rect 526982 184898 527066 185134
rect 527302 184898 527334 185134
rect 526714 167454 527334 184898
rect 526714 167218 526746 167454
rect 526982 167218 527066 167454
rect 527302 167218 527334 167454
rect 526714 167134 527334 167218
rect 526714 166898 526746 167134
rect 526982 166898 527066 167134
rect 527302 166898 527334 167134
rect 526714 149454 527334 166898
rect 526714 149218 526746 149454
rect 526982 149218 527066 149454
rect 527302 149218 527334 149454
rect 526714 149134 527334 149218
rect 526714 148898 526746 149134
rect 526982 148898 527066 149134
rect 527302 148898 527334 149134
rect 526714 131454 527334 148898
rect 526714 131218 526746 131454
rect 526982 131218 527066 131454
rect 527302 131218 527334 131454
rect 526714 131134 527334 131218
rect 526714 130898 526746 131134
rect 526982 130898 527066 131134
rect 527302 130898 527334 131134
rect 526714 113454 527334 130898
rect 526714 113218 526746 113454
rect 526982 113218 527066 113454
rect 527302 113218 527334 113454
rect 526714 113134 527334 113218
rect 526714 112898 526746 113134
rect 526982 112898 527066 113134
rect 527302 112898 527334 113134
rect 526714 95454 527334 112898
rect 526714 95218 526746 95454
rect 526982 95218 527066 95454
rect 527302 95218 527334 95454
rect 526714 95134 527334 95218
rect 526714 94898 526746 95134
rect 526982 94898 527066 95134
rect 527302 94898 527334 95134
rect 526714 77454 527334 94898
rect 526714 77218 526746 77454
rect 526982 77218 527066 77454
rect 527302 77218 527334 77454
rect 526714 77134 527334 77218
rect 526714 76898 526746 77134
rect 526982 76898 527066 77134
rect 527302 76898 527334 77134
rect 526714 59454 527334 76898
rect 526714 59218 526746 59454
rect 526982 59218 527066 59454
rect 527302 59218 527334 59454
rect 526714 59134 527334 59218
rect 526714 58898 526746 59134
rect 526982 58898 527066 59134
rect 527302 58898 527334 59134
rect 526714 41454 527334 58898
rect 526714 41218 526746 41454
rect 526982 41218 527066 41454
rect 527302 41218 527334 41454
rect 526714 41134 527334 41218
rect 526714 40898 526746 41134
rect 526982 40898 527066 41134
rect 527302 40898 527334 41134
rect 526714 23454 527334 40898
rect 526714 23218 526746 23454
rect 526982 23218 527066 23454
rect 527302 23218 527334 23454
rect 526714 23134 527334 23218
rect 526714 22898 526746 23134
rect 526982 22898 527066 23134
rect 527302 22898 527334 23134
rect 526714 5454 527334 22898
rect 526714 5218 526746 5454
rect 526982 5218 527066 5454
rect 527302 5218 527334 5454
rect 526714 5134 527334 5218
rect 526714 4898 526746 5134
rect 526982 4898 527066 5134
rect 527302 4898 527334 5134
rect 526714 880 527334 4898
rect 530434 462052 531054 464004
rect 530434 461816 530466 462052
rect 530702 461816 530786 462052
rect 531022 461816 531054 462052
rect 530434 461732 531054 461816
rect 530434 461496 530466 461732
rect 530702 461496 530786 461732
rect 531022 461496 531054 461732
rect 530434 441174 531054 461496
rect 530434 440938 530466 441174
rect 530702 440938 530786 441174
rect 531022 440938 531054 441174
rect 530434 440854 531054 440938
rect 530434 440618 530466 440854
rect 530702 440618 530786 440854
rect 531022 440618 531054 440854
rect 530434 423174 531054 440618
rect 530434 422938 530466 423174
rect 530702 422938 530786 423174
rect 531022 422938 531054 423174
rect 530434 422854 531054 422938
rect 530434 422618 530466 422854
rect 530702 422618 530786 422854
rect 531022 422618 531054 422854
rect 530434 405174 531054 422618
rect 530434 404938 530466 405174
rect 530702 404938 530786 405174
rect 531022 404938 531054 405174
rect 530434 404854 531054 404938
rect 530434 404618 530466 404854
rect 530702 404618 530786 404854
rect 531022 404618 531054 404854
rect 530434 387174 531054 404618
rect 530434 386938 530466 387174
rect 530702 386938 530786 387174
rect 531022 386938 531054 387174
rect 530434 386854 531054 386938
rect 530434 386618 530466 386854
rect 530702 386618 530786 386854
rect 531022 386618 531054 386854
rect 530434 369174 531054 386618
rect 530434 368938 530466 369174
rect 530702 368938 530786 369174
rect 531022 368938 531054 369174
rect 530434 368854 531054 368938
rect 530434 368618 530466 368854
rect 530702 368618 530786 368854
rect 531022 368618 531054 368854
rect 530434 351174 531054 368618
rect 530434 350938 530466 351174
rect 530702 350938 530786 351174
rect 531022 350938 531054 351174
rect 530434 350854 531054 350938
rect 530434 350618 530466 350854
rect 530702 350618 530786 350854
rect 531022 350618 531054 350854
rect 530434 333174 531054 350618
rect 530434 332938 530466 333174
rect 530702 332938 530786 333174
rect 531022 332938 531054 333174
rect 530434 332854 531054 332938
rect 530434 332618 530466 332854
rect 530702 332618 530786 332854
rect 531022 332618 531054 332854
rect 530434 315174 531054 332618
rect 530434 314938 530466 315174
rect 530702 314938 530786 315174
rect 531022 314938 531054 315174
rect 530434 314854 531054 314938
rect 530434 314618 530466 314854
rect 530702 314618 530786 314854
rect 531022 314618 531054 314854
rect 530434 297174 531054 314618
rect 530434 296938 530466 297174
rect 530702 296938 530786 297174
rect 531022 296938 531054 297174
rect 530434 296854 531054 296938
rect 530434 296618 530466 296854
rect 530702 296618 530786 296854
rect 531022 296618 531054 296854
rect 530434 279174 531054 296618
rect 530434 278938 530466 279174
rect 530702 278938 530786 279174
rect 531022 278938 531054 279174
rect 530434 278854 531054 278938
rect 530434 278618 530466 278854
rect 530702 278618 530786 278854
rect 531022 278618 531054 278854
rect 530434 261174 531054 278618
rect 530434 260938 530466 261174
rect 530702 260938 530786 261174
rect 531022 260938 531054 261174
rect 530434 260854 531054 260938
rect 530434 260618 530466 260854
rect 530702 260618 530786 260854
rect 531022 260618 531054 260854
rect 530434 243174 531054 260618
rect 530434 242938 530466 243174
rect 530702 242938 530786 243174
rect 531022 242938 531054 243174
rect 530434 242854 531054 242938
rect 530434 242618 530466 242854
rect 530702 242618 530786 242854
rect 531022 242618 531054 242854
rect 530434 225174 531054 242618
rect 530434 224938 530466 225174
rect 530702 224938 530786 225174
rect 531022 224938 531054 225174
rect 530434 224854 531054 224938
rect 530434 224618 530466 224854
rect 530702 224618 530786 224854
rect 531022 224618 531054 224854
rect 530434 207174 531054 224618
rect 530434 206938 530466 207174
rect 530702 206938 530786 207174
rect 531022 206938 531054 207174
rect 530434 206854 531054 206938
rect 530434 206618 530466 206854
rect 530702 206618 530786 206854
rect 531022 206618 531054 206854
rect 530434 189174 531054 206618
rect 530434 188938 530466 189174
rect 530702 188938 530786 189174
rect 531022 188938 531054 189174
rect 530434 188854 531054 188938
rect 530434 188618 530466 188854
rect 530702 188618 530786 188854
rect 531022 188618 531054 188854
rect 530434 171174 531054 188618
rect 530434 170938 530466 171174
rect 530702 170938 530786 171174
rect 531022 170938 531054 171174
rect 530434 170854 531054 170938
rect 530434 170618 530466 170854
rect 530702 170618 530786 170854
rect 531022 170618 531054 170854
rect 530434 153174 531054 170618
rect 530434 152938 530466 153174
rect 530702 152938 530786 153174
rect 531022 152938 531054 153174
rect 530434 152854 531054 152938
rect 530434 152618 530466 152854
rect 530702 152618 530786 152854
rect 531022 152618 531054 152854
rect 530434 135174 531054 152618
rect 530434 134938 530466 135174
rect 530702 134938 530786 135174
rect 531022 134938 531054 135174
rect 530434 134854 531054 134938
rect 530434 134618 530466 134854
rect 530702 134618 530786 134854
rect 531022 134618 531054 134854
rect 530434 117174 531054 134618
rect 530434 116938 530466 117174
rect 530702 116938 530786 117174
rect 531022 116938 531054 117174
rect 530434 116854 531054 116938
rect 530434 116618 530466 116854
rect 530702 116618 530786 116854
rect 531022 116618 531054 116854
rect 530434 99174 531054 116618
rect 530434 98938 530466 99174
rect 530702 98938 530786 99174
rect 531022 98938 531054 99174
rect 530434 98854 531054 98938
rect 530434 98618 530466 98854
rect 530702 98618 530786 98854
rect 531022 98618 531054 98854
rect 530434 81174 531054 98618
rect 530434 80938 530466 81174
rect 530702 80938 530786 81174
rect 531022 80938 531054 81174
rect 530434 80854 531054 80938
rect 530434 80618 530466 80854
rect 530702 80618 530786 80854
rect 531022 80618 531054 80854
rect 530434 63174 531054 80618
rect 530434 62938 530466 63174
rect 530702 62938 530786 63174
rect 531022 62938 531054 63174
rect 530434 62854 531054 62938
rect 530434 62618 530466 62854
rect 530702 62618 530786 62854
rect 531022 62618 531054 62854
rect 530434 45174 531054 62618
rect 530434 44938 530466 45174
rect 530702 44938 530786 45174
rect 531022 44938 531054 45174
rect 530434 44854 531054 44938
rect 530434 44618 530466 44854
rect 530702 44618 530786 44854
rect 531022 44618 531054 44854
rect 530434 27174 531054 44618
rect 530434 26938 530466 27174
rect 530702 26938 530786 27174
rect 531022 26938 531054 27174
rect 530434 26854 531054 26938
rect 530434 26618 530466 26854
rect 530702 26618 530786 26854
rect 531022 26618 531054 26854
rect 530434 9174 531054 26618
rect 530434 8938 530466 9174
rect 530702 8938 530786 9174
rect 531022 8938 531054 9174
rect 530434 8854 531054 8938
rect 530434 8618 530466 8854
rect 530702 8618 530786 8854
rect 531022 8618 531054 8854
rect 530434 880 531054 8618
rect 534154 463012 534774 464004
rect 534154 462776 534186 463012
rect 534422 462776 534506 463012
rect 534742 462776 534774 463012
rect 534154 462692 534774 462776
rect 534154 462456 534186 462692
rect 534422 462456 534506 462692
rect 534742 462456 534774 462692
rect 534154 444894 534774 462456
rect 534154 444658 534186 444894
rect 534422 444658 534506 444894
rect 534742 444658 534774 444894
rect 534154 444574 534774 444658
rect 534154 444338 534186 444574
rect 534422 444338 534506 444574
rect 534742 444338 534774 444574
rect 534154 426894 534774 444338
rect 534154 426658 534186 426894
rect 534422 426658 534506 426894
rect 534742 426658 534774 426894
rect 534154 426574 534774 426658
rect 534154 426338 534186 426574
rect 534422 426338 534506 426574
rect 534742 426338 534774 426574
rect 534154 408894 534774 426338
rect 534154 408658 534186 408894
rect 534422 408658 534506 408894
rect 534742 408658 534774 408894
rect 534154 408574 534774 408658
rect 534154 408338 534186 408574
rect 534422 408338 534506 408574
rect 534742 408338 534774 408574
rect 534154 390894 534774 408338
rect 534154 390658 534186 390894
rect 534422 390658 534506 390894
rect 534742 390658 534774 390894
rect 534154 390574 534774 390658
rect 534154 390338 534186 390574
rect 534422 390338 534506 390574
rect 534742 390338 534774 390574
rect 534154 372894 534774 390338
rect 534154 372658 534186 372894
rect 534422 372658 534506 372894
rect 534742 372658 534774 372894
rect 534154 372574 534774 372658
rect 534154 372338 534186 372574
rect 534422 372338 534506 372574
rect 534742 372338 534774 372574
rect 534154 354894 534774 372338
rect 534154 354658 534186 354894
rect 534422 354658 534506 354894
rect 534742 354658 534774 354894
rect 534154 354574 534774 354658
rect 534154 354338 534186 354574
rect 534422 354338 534506 354574
rect 534742 354338 534774 354574
rect 534154 336894 534774 354338
rect 534154 336658 534186 336894
rect 534422 336658 534506 336894
rect 534742 336658 534774 336894
rect 534154 336574 534774 336658
rect 534154 336338 534186 336574
rect 534422 336338 534506 336574
rect 534742 336338 534774 336574
rect 534154 318894 534774 336338
rect 534154 318658 534186 318894
rect 534422 318658 534506 318894
rect 534742 318658 534774 318894
rect 534154 318574 534774 318658
rect 534154 318338 534186 318574
rect 534422 318338 534506 318574
rect 534742 318338 534774 318574
rect 534154 300894 534774 318338
rect 534154 300658 534186 300894
rect 534422 300658 534506 300894
rect 534742 300658 534774 300894
rect 534154 300574 534774 300658
rect 534154 300338 534186 300574
rect 534422 300338 534506 300574
rect 534742 300338 534774 300574
rect 534154 282894 534774 300338
rect 534154 282658 534186 282894
rect 534422 282658 534506 282894
rect 534742 282658 534774 282894
rect 534154 282574 534774 282658
rect 534154 282338 534186 282574
rect 534422 282338 534506 282574
rect 534742 282338 534774 282574
rect 534154 264894 534774 282338
rect 534154 264658 534186 264894
rect 534422 264658 534506 264894
rect 534742 264658 534774 264894
rect 534154 264574 534774 264658
rect 534154 264338 534186 264574
rect 534422 264338 534506 264574
rect 534742 264338 534774 264574
rect 534154 246894 534774 264338
rect 534154 246658 534186 246894
rect 534422 246658 534506 246894
rect 534742 246658 534774 246894
rect 534154 246574 534774 246658
rect 534154 246338 534186 246574
rect 534422 246338 534506 246574
rect 534742 246338 534774 246574
rect 534154 228894 534774 246338
rect 534154 228658 534186 228894
rect 534422 228658 534506 228894
rect 534742 228658 534774 228894
rect 534154 228574 534774 228658
rect 534154 228338 534186 228574
rect 534422 228338 534506 228574
rect 534742 228338 534774 228574
rect 534154 210894 534774 228338
rect 534154 210658 534186 210894
rect 534422 210658 534506 210894
rect 534742 210658 534774 210894
rect 534154 210574 534774 210658
rect 534154 210338 534186 210574
rect 534422 210338 534506 210574
rect 534742 210338 534774 210574
rect 534154 192894 534774 210338
rect 534154 192658 534186 192894
rect 534422 192658 534506 192894
rect 534742 192658 534774 192894
rect 534154 192574 534774 192658
rect 534154 192338 534186 192574
rect 534422 192338 534506 192574
rect 534742 192338 534774 192574
rect 534154 174894 534774 192338
rect 534154 174658 534186 174894
rect 534422 174658 534506 174894
rect 534742 174658 534774 174894
rect 534154 174574 534774 174658
rect 534154 174338 534186 174574
rect 534422 174338 534506 174574
rect 534742 174338 534774 174574
rect 534154 156894 534774 174338
rect 534154 156658 534186 156894
rect 534422 156658 534506 156894
rect 534742 156658 534774 156894
rect 534154 156574 534774 156658
rect 534154 156338 534186 156574
rect 534422 156338 534506 156574
rect 534742 156338 534774 156574
rect 534154 138894 534774 156338
rect 534154 138658 534186 138894
rect 534422 138658 534506 138894
rect 534742 138658 534774 138894
rect 534154 138574 534774 138658
rect 534154 138338 534186 138574
rect 534422 138338 534506 138574
rect 534742 138338 534774 138574
rect 534154 120894 534774 138338
rect 534154 120658 534186 120894
rect 534422 120658 534506 120894
rect 534742 120658 534774 120894
rect 534154 120574 534774 120658
rect 534154 120338 534186 120574
rect 534422 120338 534506 120574
rect 534742 120338 534774 120574
rect 534154 102894 534774 120338
rect 534154 102658 534186 102894
rect 534422 102658 534506 102894
rect 534742 102658 534774 102894
rect 534154 102574 534774 102658
rect 534154 102338 534186 102574
rect 534422 102338 534506 102574
rect 534742 102338 534774 102574
rect 534154 84894 534774 102338
rect 534154 84658 534186 84894
rect 534422 84658 534506 84894
rect 534742 84658 534774 84894
rect 534154 84574 534774 84658
rect 534154 84338 534186 84574
rect 534422 84338 534506 84574
rect 534742 84338 534774 84574
rect 534154 66894 534774 84338
rect 534154 66658 534186 66894
rect 534422 66658 534506 66894
rect 534742 66658 534774 66894
rect 534154 66574 534774 66658
rect 534154 66338 534186 66574
rect 534422 66338 534506 66574
rect 534742 66338 534774 66574
rect 534154 48894 534774 66338
rect 534154 48658 534186 48894
rect 534422 48658 534506 48894
rect 534742 48658 534774 48894
rect 534154 48574 534774 48658
rect 534154 48338 534186 48574
rect 534422 48338 534506 48574
rect 534742 48338 534774 48574
rect 534154 30894 534774 48338
rect 534154 30658 534186 30894
rect 534422 30658 534506 30894
rect 534742 30658 534774 30894
rect 534154 30574 534774 30658
rect 534154 30338 534186 30574
rect 534422 30338 534506 30574
rect 534742 30338 534774 30574
rect 534154 12894 534774 30338
rect 534154 12658 534186 12894
rect 534422 12658 534506 12894
rect 534742 12658 534774 12894
rect 534154 12574 534774 12658
rect 534154 12338 534186 12574
rect 534422 12338 534506 12574
rect 534742 12338 534774 12574
rect 534154 880 534774 12338
rect 537874 463972 538494 464004
rect 537874 463736 537906 463972
rect 538142 463736 538226 463972
rect 538462 463736 538494 463972
rect 537874 463652 538494 463736
rect 537874 463416 537906 463652
rect 538142 463416 538226 463652
rect 538462 463416 538494 463652
rect 537874 448614 538494 463416
rect 547852 463972 548472 464004
rect 547852 463736 547884 463972
rect 548120 463736 548204 463972
rect 548440 463736 548472 463972
rect 547852 463652 548472 463736
rect 547852 463416 547884 463652
rect 548120 463416 548204 463652
rect 548440 463416 548472 463652
rect 546892 463012 547512 463044
rect 546892 462776 546924 463012
rect 547160 462776 547244 463012
rect 547480 462776 547512 463012
rect 546892 462692 547512 462776
rect 546892 462456 546924 462692
rect 547160 462456 547244 462692
rect 547480 462456 547512 462692
rect 545932 462052 546552 462084
rect 545932 461816 545964 462052
rect 546200 461816 546284 462052
rect 546520 461816 546552 462052
rect 545932 461732 546552 461816
rect 545932 461496 545964 461732
rect 546200 461496 546284 461732
rect 546520 461496 546552 461732
rect 537874 448378 537906 448614
rect 538142 448378 538226 448614
rect 538462 448378 538494 448614
rect 537874 448294 538494 448378
rect 537874 448058 537906 448294
rect 538142 448058 538226 448294
rect 538462 448058 538494 448294
rect 537874 430614 538494 448058
rect 537874 430378 537906 430614
rect 538142 430378 538226 430614
rect 538462 430378 538494 430614
rect 537874 430294 538494 430378
rect 537874 430058 537906 430294
rect 538142 430058 538226 430294
rect 538462 430058 538494 430294
rect 537874 412614 538494 430058
rect 537874 412378 537906 412614
rect 538142 412378 538226 412614
rect 538462 412378 538494 412614
rect 537874 412294 538494 412378
rect 537874 412058 537906 412294
rect 538142 412058 538226 412294
rect 538462 412058 538494 412294
rect 537874 394614 538494 412058
rect 537874 394378 537906 394614
rect 538142 394378 538226 394614
rect 538462 394378 538494 394614
rect 537874 394294 538494 394378
rect 537874 394058 537906 394294
rect 538142 394058 538226 394294
rect 538462 394058 538494 394294
rect 537874 376614 538494 394058
rect 537874 376378 537906 376614
rect 538142 376378 538226 376614
rect 538462 376378 538494 376614
rect 537874 376294 538494 376378
rect 537874 376058 537906 376294
rect 538142 376058 538226 376294
rect 538462 376058 538494 376294
rect 537874 358614 538494 376058
rect 537874 358378 537906 358614
rect 538142 358378 538226 358614
rect 538462 358378 538494 358614
rect 537874 358294 538494 358378
rect 537874 358058 537906 358294
rect 538142 358058 538226 358294
rect 538462 358058 538494 358294
rect 537874 340614 538494 358058
rect 537874 340378 537906 340614
rect 538142 340378 538226 340614
rect 538462 340378 538494 340614
rect 537874 340294 538494 340378
rect 537874 340058 537906 340294
rect 538142 340058 538226 340294
rect 538462 340058 538494 340294
rect 537874 322614 538494 340058
rect 537874 322378 537906 322614
rect 538142 322378 538226 322614
rect 538462 322378 538494 322614
rect 537874 322294 538494 322378
rect 537874 322058 537906 322294
rect 538142 322058 538226 322294
rect 538462 322058 538494 322294
rect 537874 304614 538494 322058
rect 537874 304378 537906 304614
rect 538142 304378 538226 304614
rect 538462 304378 538494 304614
rect 537874 304294 538494 304378
rect 537874 304058 537906 304294
rect 538142 304058 538226 304294
rect 538462 304058 538494 304294
rect 537874 286614 538494 304058
rect 537874 286378 537906 286614
rect 538142 286378 538226 286614
rect 538462 286378 538494 286614
rect 537874 286294 538494 286378
rect 537874 286058 537906 286294
rect 538142 286058 538226 286294
rect 538462 286058 538494 286294
rect 537874 268614 538494 286058
rect 537874 268378 537906 268614
rect 538142 268378 538226 268614
rect 538462 268378 538494 268614
rect 537874 268294 538494 268378
rect 537874 268058 537906 268294
rect 538142 268058 538226 268294
rect 538462 268058 538494 268294
rect 537874 250614 538494 268058
rect 537874 250378 537906 250614
rect 538142 250378 538226 250614
rect 538462 250378 538494 250614
rect 537874 250294 538494 250378
rect 537874 250058 537906 250294
rect 538142 250058 538226 250294
rect 538462 250058 538494 250294
rect 537874 232614 538494 250058
rect 537874 232378 537906 232614
rect 538142 232378 538226 232614
rect 538462 232378 538494 232614
rect 537874 232294 538494 232378
rect 537874 232058 537906 232294
rect 538142 232058 538226 232294
rect 538462 232058 538494 232294
rect 537874 214614 538494 232058
rect 537874 214378 537906 214614
rect 538142 214378 538226 214614
rect 538462 214378 538494 214614
rect 537874 214294 538494 214378
rect 537874 214058 537906 214294
rect 538142 214058 538226 214294
rect 538462 214058 538494 214294
rect 537874 196614 538494 214058
rect 537874 196378 537906 196614
rect 538142 196378 538226 196614
rect 538462 196378 538494 196614
rect 537874 196294 538494 196378
rect 537874 196058 537906 196294
rect 538142 196058 538226 196294
rect 538462 196058 538494 196294
rect 537874 178614 538494 196058
rect 537874 178378 537906 178614
rect 538142 178378 538226 178614
rect 538462 178378 538494 178614
rect 537874 178294 538494 178378
rect 537874 178058 537906 178294
rect 538142 178058 538226 178294
rect 538462 178058 538494 178294
rect 537874 160614 538494 178058
rect 537874 160378 537906 160614
rect 538142 160378 538226 160614
rect 538462 160378 538494 160614
rect 537874 160294 538494 160378
rect 537874 160058 537906 160294
rect 538142 160058 538226 160294
rect 538462 160058 538494 160294
rect 537874 142614 538494 160058
rect 537874 142378 537906 142614
rect 538142 142378 538226 142614
rect 538462 142378 538494 142614
rect 537874 142294 538494 142378
rect 537874 142058 537906 142294
rect 538142 142058 538226 142294
rect 538462 142058 538494 142294
rect 537874 124614 538494 142058
rect 537874 124378 537906 124614
rect 538142 124378 538226 124614
rect 538462 124378 538494 124614
rect 537874 124294 538494 124378
rect 537874 124058 537906 124294
rect 538142 124058 538226 124294
rect 538462 124058 538494 124294
rect 537874 106614 538494 124058
rect 537874 106378 537906 106614
rect 538142 106378 538226 106614
rect 538462 106378 538494 106614
rect 537874 106294 538494 106378
rect 537874 106058 537906 106294
rect 538142 106058 538226 106294
rect 538462 106058 538494 106294
rect 537874 88614 538494 106058
rect 537874 88378 537906 88614
rect 538142 88378 538226 88614
rect 538462 88378 538494 88614
rect 537874 88294 538494 88378
rect 537874 88058 537906 88294
rect 538142 88058 538226 88294
rect 538462 88058 538494 88294
rect 537874 70614 538494 88058
rect 537874 70378 537906 70614
rect 538142 70378 538226 70614
rect 538462 70378 538494 70614
rect 537874 70294 538494 70378
rect 537874 70058 537906 70294
rect 538142 70058 538226 70294
rect 538462 70058 538494 70294
rect 537874 52614 538494 70058
rect 537874 52378 537906 52614
rect 538142 52378 538226 52614
rect 538462 52378 538494 52614
rect 537874 52294 538494 52378
rect 537874 52058 537906 52294
rect 538142 52058 538226 52294
rect 538462 52058 538494 52294
rect 537874 34614 538494 52058
rect 537874 34378 537906 34614
rect 538142 34378 538226 34614
rect 538462 34378 538494 34614
rect 537874 34294 538494 34378
rect 537874 34058 537906 34294
rect 538142 34058 538226 34294
rect 538462 34058 538494 34294
rect 537874 16614 538494 34058
rect 537874 16378 537906 16614
rect 538142 16378 538226 16614
rect 538462 16378 538494 16614
rect 537874 16294 538494 16378
rect 537874 16058 537906 16294
rect 538142 16058 538226 16294
rect 538462 16058 538494 16294
rect 537874 880 538494 16058
rect 544972 461092 545592 461124
rect 544972 460856 545004 461092
rect 545240 460856 545324 461092
rect 545560 460856 545592 461092
rect 544972 460772 545592 460856
rect 544972 460536 545004 460772
rect 545240 460536 545324 460772
rect 545560 460536 545592 460772
rect 544972 455454 545592 460536
rect 544972 455218 545004 455454
rect 545240 455218 545324 455454
rect 545560 455218 545592 455454
rect 544972 455134 545592 455218
rect 544972 454898 545004 455134
rect 545240 454898 545324 455134
rect 545560 454898 545592 455134
rect 544972 437454 545592 454898
rect 544972 437218 545004 437454
rect 545240 437218 545324 437454
rect 545560 437218 545592 437454
rect 544972 437134 545592 437218
rect 544972 436898 545004 437134
rect 545240 436898 545324 437134
rect 545560 436898 545592 437134
rect 544972 419454 545592 436898
rect 544972 419218 545004 419454
rect 545240 419218 545324 419454
rect 545560 419218 545592 419454
rect 544972 419134 545592 419218
rect 544972 418898 545004 419134
rect 545240 418898 545324 419134
rect 545560 418898 545592 419134
rect 544972 401454 545592 418898
rect 544972 401218 545004 401454
rect 545240 401218 545324 401454
rect 545560 401218 545592 401454
rect 544972 401134 545592 401218
rect 544972 400898 545004 401134
rect 545240 400898 545324 401134
rect 545560 400898 545592 401134
rect 544972 383454 545592 400898
rect 544972 383218 545004 383454
rect 545240 383218 545324 383454
rect 545560 383218 545592 383454
rect 544972 383134 545592 383218
rect 544972 382898 545004 383134
rect 545240 382898 545324 383134
rect 545560 382898 545592 383134
rect 544972 365454 545592 382898
rect 544972 365218 545004 365454
rect 545240 365218 545324 365454
rect 545560 365218 545592 365454
rect 544972 365134 545592 365218
rect 544972 364898 545004 365134
rect 545240 364898 545324 365134
rect 545560 364898 545592 365134
rect 544972 347454 545592 364898
rect 544972 347218 545004 347454
rect 545240 347218 545324 347454
rect 545560 347218 545592 347454
rect 544972 347134 545592 347218
rect 544972 346898 545004 347134
rect 545240 346898 545324 347134
rect 545560 346898 545592 347134
rect 544972 329454 545592 346898
rect 544972 329218 545004 329454
rect 545240 329218 545324 329454
rect 545560 329218 545592 329454
rect 544972 329134 545592 329218
rect 544972 328898 545004 329134
rect 545240 328898 545324 329134
rect 545560 328898 545592 329134
rect 544972 311454 545592 328898
rect 544972 311218 545004 311454
rect 545240 311218 545324 311454
rect 545560 311218 545592 311454
rect 544972 311134 545592 311218
rect 544972 310898 545004 311134
rect 545240 310898 545324 311134
rect 545560 310898 545592 311134
rect 544972 293454 545592 310898
rect 544972 293218 545004 293454
rect 545240 293218 545324 293454
rect 545560 293218 545592 293454
rect 544972 293134 545592 293218
rect 544972 292898 545004 293134
rect 545240 292898 545324 293134
rect 545560 292898 545592 293134
rect 544972 275454 545592 292898
rect 544972 275218 545004 275454
rect 545240 275218 545324 275454
rect 545560 275218 545592 275454
rect 544972 275134 545592 275218
rect 544972 274898 545004 275134
rect 545240 274898 545324 275134
rect 545560 274898 545592 275134
rect 544972 257454 545592 274898
rect 544972 257218 545004 257454
rect 545240 257218 545324 257454
rect 545560 257218 545592 257454
rect 544972 257134 545592 257218
rect 544972 256898 545004 257134
rect 545240 256898 545324 257134
rect 545560 256898 545592 257134
rect 544972 239454 545592 256898
rect 544972 239218 545004 239454
rect 545240 239218 545324 239454
rect 545560 239218 545592 239454
rect 544972 239134 545592 239218
rect 544972 238898 545004 239134
rect 545240 238898 545324 239134
rect 545560 238898 545592 239134
rect 544972 221454 545592 238898
rect 544972 221218 545004 221454
rect 545240 221218 545324 221454
rect 545560 221218 545592 221454
rect 544972 221134 545592 221218
rect 544972 220898 545004 221134
rect 545240 220898 545324 221134
rect 545560 220898 545592 221134
rect 544972 203454 545592 220898
rect 544972 203218 545004 203454
rect 545240 203218 545324 203454
rect 545560 203218 545592 203454
rect 544972 203134 545592 203218
rect 544972 202898 545004 203134
rect 545240 202898 545324 203134
rect 545560 202898 545592 203134
rect 544972 185454 545592 202898
rect 544972 185218 545004 185454
rect 545240 185218 545324 185454
rect 545560 185218 545592 185454
rect 544972 185134 545592 185218
rect 544972 184898 545004 185134
rect 545240 184898 545324 185134
rect 545560 184898 545592 185134
rect 544972 167454 545592 184898
rect 544972 167218 545004 167454
rect 545240 167218 545324 167454
rect 545560 167218 545592 167454
rect 544972 167134 545592 167218
rect 544972 166898 545004 167134
rect 545240 166898 545324 167134
rect 545560 166898 545592 167134
rect 544972 149454 545592 166898
rect 544972 149218 545004 149454
rect 545240 149218 545324 149454
rect 545560 149218 545592 149454
rect 544972 149134 545592 149218
rect 544972 148898 545004 149134
rect 545240 148898 545324 149134
rect 545560 148898 545592 149134
rect 544972 131454 545592 148898
rect 544972 131218 545004 131454
rect 545240 131218 545324 131454
rect 545560 131218 545592 131454
rect 544972 131134 545592 131218
rect 544972 130898 545004 131134
rect 545240 130898 545324 131134
rect 545560 130898 545592 131134
rect 544972 113454 545592 130898
rect 544972 113218 545004 113454
rect 545240 113218 545324 113454
rect 545560 113218 545592 113454
rect 544972 113134 545592 113218
rect 544972 112898 545004 113134
rect 545240 112898 545324 113134
rect 545560 112898 545592 113134
rect 544972 95454 545592 112898
rect 544972 95218 545004 95454
rect 545240 95218 545324 95454
rect 545560 95218 545592 95454
rect 544972 95134 545592 95218
rect 544972 94898 545004 95134
rect 545240 94898 545324 95134
rect 545560 94898 545592 95134
rect 544972 77454 545592 94898
rect 544972 77218 545004 77454
rect 545240 77218 545324 77454
rect 545560 77218 545592 77454
rect 544972 77134 545592 77218
rect 544972 76898 545004 77134
rect 545240 76898 545324 77134
rect 545560 76898 545592 77134
rect 544972 59454 545592 76898
rect 544972 59218 545004 59454
rect 545240 59218 545324 59454
rect 545560 59218 545592 59454
rect 544972 59134 545592 59218
rect 544972 58898 545004 59134
rect 545240 58898 545324 59134
rect 545560 58898 545592 59134
rect 544972 41454 545592 58898
rect 544972 41218 545004 41454
rect 545240 41218 545324 41454
rect 545560 41218 545592 41454
rect 544972 41134 545592 41218
rect 544972 40898 545004 41134
rect 545240 40898 545324 41134
rect 545560 40898 545592 41134
rect 544972 23454 545592 40898
rect 544972 23218 545004 23454
rect 545240 23218 545324 23454
rect 545560 23218 545592 23454
rect 544972 23134 545592 23218
rect 544972 22898 545004 23134
rect 545240 22898 545324 23134
rect 545560 22898 545592 23134
rect 544972 5454 545592 22898
rect 544972 5218 545004 5454
rect 545240 5218 545324 5454
rect 545560 5218 545592 5454
rect 544972 5134 545592 5218
rect 544972 4898 545004 5134
rect 545240 4898 545324 5134
rect 545560 4898 545592 5134
rect 500302 0 505082 638
rect 510281 0 515061 638
rect 524302 0 529082 638
rect 534281 0 539061 638
rect 544972 -856 545592 4898
rect 544972 -1092 545004 -856
rect 545240 -1092 545324 -856
rect 545560 -1092 545592 -856
rect 544972 -1176 545592 -1092
rect 544972 -1412 545004 -1176
rect 545240 -1412 545324 -1176
rect 545560 -1412 545592 -1176
rect 544972 -1444 545592 -1412
rect 545932 441174 546552 461496
rect 545932 440938 545964 441174
rect 546200 440938 546284 441174
rect 546520 440938 546552 441174
rect 545932 440854 546552 440938
rect 545932 440618 545964 440854
rect 546200 440618 546284 440854
rect 546520 440618 546552 440854
rect 545932 423174 546552 440618
rect 545932 422938 545964 423174
rect 546200 422938 546284 423174
rect 546520 422938 546552 423174
rect 545932 422854 546552 422938
rect 545932 422618 545964 422854
rect 546200 422618 546284 422854
rect 546520 422618 546552 422854
rect 545932 405174 546552 422618
rect 545932 404938 545964 405174
rect 546200 404938 546284 405174
rect 546520 404938 546552 405174
rect 545932 404854 546552 404938
rect 545932 404618 545964 404854
rect 546200 404618 546284 404854
rect 546520 404618 546552 404854
rect 545932 387174 546552 404618
rect 545932 386938 545964 387174
rect 546200 386938 546284 387174
rect 546520 386938 546552 387174
rect 545932 386854 546552 386938
rect 545932 386618 545964 386854
rect 546200 386618 546284 386854
rect 546520 386618 546552 386854
rect 545932 369174 546552 386618
rect 545932 368938 545964 369174
rect 546200 368938 546284 369174
rect 546520 368938 546552 369174
rect 545932 368854 546552 368938
rect 545932 368618 545964 368854
rect 546200 368618 546284 368854
rect 546520 368618 546552 368854
rect 545932 351174 546552 368618
rect 545932 350938 545964 351174
rect 546200 350938 546284 351174
rect 546520 350938 546552 351174
rect 545932 350854 546552 350938
rect 545932 350618 545964 350854
rect 546200 350618 546284 350854
rect 546520 350618 546552 350854
rect 545932 333174 546552 350618
rect 545932 332938 545964 333174
rect 546200 332938 546284 333174
rect 546520 332938 546552 333174
rect 545932 332854 546552 332938
rect 545932 332618 545964 332854
rect 546200 332618 546284 332854
rect 546520 332618 546552 332854
rect 545932 315174 546552 332618
rect 545932 314938 545964 315174
rect 546200 314938 546284 315174
rect 546520 314938 546552 315174
rect 545932 314854 546552 314938
rect 545932 314618 545964 314854
rect 546200 314618 546284 314854
rect 546520 314618 546552 314854
rect 545932 297174 546552 314618
rect 545932 296938 545964 297174
rect 546200 296938 546284 297174
rect 546520 296938 546552 297174
rect 545932 296854 546552 296938
rect 545932 296618 545964 296854
rect 546200 296618 546284 296854
rect 546520 296618 546552 296854
rect 545932 279174 546552 296618
rect 545932 278938 545964 279174
rect 546200 278938 546284 279174
rect 546520 278938 546552 279174
rect 545932 278854 546552 278938
rect 545932 278618 545964 278854
rect 546200 278618 546284 278854
rect 546520 278618 546552 278854
rect 545932 261174 546552 278618
rect 545932 260938 545964 261174
rect 546200 260938 546284 261174
rect 546520 260938 546552 261174
rect 545932 260854 546552 260938
rect 545932 260618 545964 260854
rect 546200 260618 546284 260854
rect 546520 260618 546552 260854
rect 545932 243174 546552 260618
rect 545932 242938 545964 243174
rect 546200 242938 546284 243174
rect 546520 242938 546552 243174
rect 545932 242854 546552 242938
rect 545932 242618 545964 242854
rect 546200 242618 546284 242854
rect 546520 242618 546552 242854
rect 545932 225174 546552 242618
rect 545932 224938 545964 225174
rect 546200 224938 546284 225174
rect 546520 224938 546552 225174
rect 545932 224854 546552 224938
rect 545932 224618 545964 224854
rect 546200 224618 546284 224854
rect 546520 224618 546552 224854
rect 545932 207174 546552 224618
rect 545932 206938 545964 207174
rect 546200 206938 546284 207174
rect 546520 206938 546552 207174
rect 545932 206854 546552 206938
rect 545932 206618 545964 206854
rect 546200 206618 546284 206854
rect 546520 206618 546552 206854
rect 545932 189174 546552 206618
rect 545932 188938 545964 189174
rect 546200 188938 546284 189174
rect 546520 188938 546552 189174
rect 545932 188854 546552 188938
rect 545932 188618 545964 188854
rect 546200 188618 546284 188854
rect 546520 188618 546552 188854
rect 545932 171174 546552 188618
rect 545932 170938 545964 171174
rect 546200 170938 546284 171174
rect 546520 170938 546552 171174
rect 545932 170854 546552 170938
rect 545932 170618 545964 170854
rect 546200 170618 546284 170854
rect 546520 170618 546552 170854
rect 545932 153174 546552 170618
rect 545932 152938 545964 153174
rect 546200 152938 546284 153174
rect 546520 152938 546552 153174
rect 545932 152854 546552 152938
rect 545932 152618 545964 152854
rect 546200 152618 546284 152854
rect 546520 152618 546552 152854
rect 545932 135174 546552 152618
rect 545932 134938 545964 135174
rect 546200 134938 546284 135174
rect 546520 134938 546552 135174
rect 545932 134854 546552 134938
rect 545932 134618 545964 134854
rect 546200 134618 546284 134854
rect 546520 134618 546552 134854
rect 545932 117174 546552 134618
rect 545932 116938 545964 117174
rect 546200 116938 546284 117174
rect 546520 116938 546552 117174
rect 545932 116854 546552 116938
rect 545932 116618 545964 116854
rect 546200 116618 546284 116854
rect 546520 116618 546552 116854
rect 545932 99174 546552 116618
rect 545932 98938 545964 99174
rect 546200 98938 546284 99174
rect 546520 98938 546552 99174
rect 545932 98854 546552 98938
rect 545932 98618 545964 98854
rect 546200 98618 546284 98854
rect 546520 98618 546552 98854
rect 545932 81174 546552 98618
rect 545932 80938 545964 81174
rect 546200 80938 546284 81174
rect 546520 80938 546552 81174
rect 545932 80854 546552 80938
rect 545932 80618 545964 80854
rect 546200 80618 546284 80854
rect 546520 80618 546552 80854
rect 545932 63174 546552 80618
rect 545932 62938 545964 63174
rect 546200 62938 546284 63174
rect 546520 62938 546552 63174
rect 545932 62854 546552 62938
rect 545932 62618 545964 62854
rect 546200 62618 546284 62854
rect 546520 62618 546552 62854
rect 545932 45174 546552 62618
rect 545932 44938 545964 45174
rect 546200 44938 546284 45174
rect 546520 44938 546552 45174
rect 545932 44854 546552 44938
rect 545932 44618 545964 44854
rect 546200 44618 546284 44854
rect 546520 44618 546552 44854
rect 545932 27174 546552 44618
rect 545932 26938 545964 27174
rect 546200 26938 546284 27174
rect 546520 26938 546552 27174
rect 545932 26854 546552 26938
rect 545932 26618 545964 26854
rect 546200 26618 546284 26854
rect 546520 26618 546552 26854
rect 545932 9174 546552 26618
rect 545932 8938 545964 9174
rect 546200 8938 546284 9174
rect 546520 8938 546552 9174
rect 545932 8854 546552 8938
rect 545932 8618 545964 8854
rect 546200 8618 546284 8854
rect 546520 8618 546552 8854
rect 545932 -1816 546552 8618
rect 545932 -2052 545964 -1816
rect 546200 -2052 546284 -1816
rect 546520 -2052 546552 -1816
rect 545932 -2136 546552 -2052
rect 545932 -2372 545964 -2136
rect 546200 -2372 546284 -2136
rect 546520 -2372 546552 -2136
rect 545932 -2404 546552 -2372
rect 546892 444894 547512 462456
rect 546892 444658 546924 444894
rect 547160 444658 547244 444894
rect 547480 444658 547512 444894
rect 546892 444574 547512 444658
rect 546892 444338 546924 444574
rect 547160 444338 547244 444574
rect 547480 444338 547512 444574
rect 546892 426894 547512 444338
rect 546892 426658 546924 426894
rect 547160 426658 547244 426894
rect 547480 426658 547512 426894
rect 546892 426574 547512 426658
rect 546892 426338 546924 426574
rect 547160 426338 547244 426574
rect 547480 426338 547512 426574
rect 546892 408894 547512 426338
rect 546892 408658 546924 408894
rect 547160 408658 547244 408894
rect 547480 408658 547512 408894
rect 546892 408574 547512 408658
rect 546892 408338 546924 408574
rect 547160 408338 547244 408574
rect 547480 408338 547512 408574
rect 546892 390894 547512 408338
rect 546892 390658 546924 390894
rect 547160 390658 547244 390894
rect 547480 390658 547512 390894
rect 546892 390574 547512 390658
rect 546892 390338 546924 390574
rect 547160 390338 547244 390574
rect 547480 390338 547512 390574
rect 546892 372894 547512 390338
rect 546892 372658 546924 372894
rect 547160 372658 547244 372894
rect 547480 372658 547512 372894
rect 546892 372574 547512 372658
rect 546892 372338 546924 372574
rect 547160 372338 547244 372574
rect 547480 372338 547512 372574
rect 546892 354894 547512 372338
rect 546892 354658 546924 354894
rect 547160 354658 547244 354894
rect 547480 354658 547512 354894
rect 546892 354574 547512 354658
rect 546892 354338 546924 354574
rect 547160 354338 547244 354574
rect 547480 354338 547512 354574
rect 546892 336894 547512 354338
rect 546892 336658 546924 336894
rect 547160 336658 547244 336894
rect 547480 336658 547512 336894
rect 546892 336574 547512 336658
rect 546892 336338 546924 336574
rect 547160 336338 547244 336574
rect 547480 336338 547512 336574
rect 546892 318894 547512 336338
rect 546892 318658 546924 318894
rect 547160 318658 547244 318894
rect 547480 318658 547512 318894
rect 546892 318574 547512 318658
rect 546892 318338 546924 318574
rect 547160 318338 547244 318574
rect 547480 318338 547512 318574
rect 546892 300894 547512 318338
rect 546892 300658 546924 300894
rect 547160 300658 547244 300894
rect 547480 300658 547512 300894
rect 546892 300574 547512 300658
rect 546892 300338 546924 300574
rect 547160 300338 547244 300574
rect 547480 300338 547512 300574
rect 546892 282894 547512 300338
rect 546892 282658 546924 282894
rect 547160 282658 547244 282894
rect 547480 282658 547512 282894
rect 546892 282574 547512 282658
rect 546892 282338 546924 282574
rect 547160 282338 547244 282574
rect 547480 282338 547512 282574
rect 546892 264894 547512 282338
rect 546892 264658 546924 264894
rect 547160 264658 547244 264894
rect 547480 264658 547512 264894
rect 546892 264574 547512 264658
rect 546892 264338 546924 264574
rect 547160 264338 547244 264574
rect 547480 264338 547512 264574
rect 546892 246894 547512 264338
rect 546892 246658 546924 246894
rect 547160 246658 547244 246894
rect 547480 246658 547512 246894
rect 546892 246574 547512 246658
rect 546892 246338 546924 246574
rect 547160 246338 547244 246574
rect 547480 246338 547512 246574
rect 546892 228894 547512 246338
rect 546892 228658 546924 228894
rect 547160 228658 547244 228894
rect 547480 228658 547512 228894
rect 546892 228574 547512 228658
rect 546892 228338 546924 228574
rect 547160 228338 547244 228574
rect 547480 228338 547512 228574
rect 546892 210894 547512 228338
rect 546892 210658 546924 210894
rect 547160 210658 547244 210894
rect 547480 210658 547512 210894
rect 546892 210574 547512 210658
rect 546892 210338 546924 210574
rect 547160 210338 547244 210574
rect 547480 210338 547512 210574
rect 546892 192894 547512 210338
rect 546892 192658 546924 192894
rect 547160 192658 547244 192894
rect 547480 192658 547512 192894
rect 546892 192574 547512 192658
rect 546892 192338 546924 192574
rect 547160 192338 547244 192574
rect 547480 192338 547512 192574
rect 546892 174894 547512 192338
rect 546892 174658 546924 174894
rect 547160 174658 547244 174894
rect 547480 174658 547512 174894
rect 546892 174574 547512 174658
rect 546892 174338 546924 174574
rect 547160 174338 547244 174574
rect 547480 174338 547512 174574
rect 546892 156894 547512 174338
rect 546892 156658 546924 156894
rect 547160 156658 547244 156894
rect 547480 156658 547512 156894
rect 546892 156574 547512 156658
rect 546892 156338 546924 156574
rect 547160 156338 547244 156574
rect 547480 156338 547512 156574
rect 546892 138894 547512 156338
rect 546892 138658 546924 138894
rect 547160 138658 547244 138894
rect 547480 138658 547512 138894
rect 546892 138574 547512 138658
rect 546892 138338 546924 138574
rect 547160 138338 547244 138574
rect 547480 138338 547512 138574
rect 546892 120894 547512 138338
rect 546892 120658 546924 120894
rect 547160 120658 547244 120894
rect 547480 120658 547512 120894
rect 546892 120574 547512 120658
rect 546892 120338 546924 120574
rect 547160 120338 547244 120574
rect 547480 120338 547512 120574
rect 546892 102894 547512 120338
rect 546892 102658 546924 102894
rect 547160 102658 547244 102894
rect 547480 102658 547512 102894
rect 546892 102574 547512 102658
rect 546892 102338 546924 102574
rect 547160 102338 547244 102574
rect 547480 102338 547512 102574
rect 546892 84894 547512 102338
rect 546892 84658 546924 84894
rect 547160 84658 547244 84894
rect 547480 84658 547512 84894
rect 546892 84574 547512 84658
rect 546892 84338 546924 84574
rect 547160 84338 547244 84574
rect 547480 84338 547512 84574
rect 546892 66894 547512 84338
rect 546892 66658 546924 66894
rect 547160 66658 547244 66894
rect 547480 66658 547512 66894
rect 546892 66574 547512 66658
rect 546892 66338 546924 66574
rect 547160 66338 547244 66574
rect 547480 66338 547512 66574
rect 546892 48894 547512 66338
rect 546892 48658 546924 48894
rect 547160 48658 547244 48894
rect 547480 48658 547512 48894
rect 546892 48574 547512 48658
rect 546892 48338 546924 48574
rect 547160 48338 547244 48574
rect 547480 48338 547512 48574
rect 546892 30894 547512 48338
rect 546892 30658 546924 30894
rect 547160 30658 547244 30894
rect 547480 30658 547512 30894
rect 546892 30574 547512 30658
rect 546892 30338 546924 30574
rect 547160 30338 547244 30574
rect 547480 30338 547512 30574
rect 546892 12894 547512 30338
rect 546892 12658 546924 12894
rect 547160 12658 547244 12894
rect 547480 12658 547512 12894
rect 546892 12574 547512 12658
rect 546892 12338 546924 12574
rect 547160 12338 547244 12574
rect 547480 12338 547512 12574
rect 498154 -3012 498186 -2776
rect 498422 -3012 498506 -2776
rect 498742 -3012 498774 -2776
rect 498154 -3096 498774 -3012
rect 498154 -3332 498186 -3096
rect 498422 -3332 498506 -3096
rect 498742 -3332 498774 -3096
rect 498154 -4324 498774 -3332
rect 546892 -2776 547512 12338
rect 546892 -3012 546924 -2776
rect 547160 -3012 547244 -2776
rect 547480 -3012 547512 -2776
rect 546892 -3096 547512 -3012
rect 546892 -3332 546924 -3096
rect 547160 -3332 547244 -3096
rect 547480 -3332 547512 -3096
rect 546892 -3364 547512 -3332
rect 547852 448614 548472 463416
rect 547852 448378 547884 448614
rect 548120 448378 548204 448614
rect 548440 448378 548472 448614
rect 547852 448294 548472 448378
rect 547852 448058 547884 448294
rect 548120 448058 548204 448294
rect 548440 448058 548472 448294
rect 547852 430614 548472 448058
rect 547852 430378 547884 430614
rect 548120 430378 548204 430614
rect 548440 430378 548472 430614
rect 547852 430294 548472 430378
rect 547852 430058 547884 430294
rect 548120 430058 548204 430294
rect 548440 430058 548472 430294
rect 547852 412614 548472 430058
rect 547852 412378 547884 412614
rect 548120 412378 548204 412614
rect 548440 412378 548472 412614
rect 547852 412294 548472 412378
rect 547852 412058 547884 412294
rect 548120 412058 548204 412294
rect 548440 412058 548472 412294
rect 547852 394614 548472 412058
rect 547852 394378 547884 394614
rect 548120 394378 548204 394614
rect 548440 394378 548472 394614
rect 547852 394294 548472 394378
rect 547852 394058 547884 394294
rect 548120 394058 548204 394294
rect 548440 394058 548472 394294
rect 547852 376614 548472 394058
rect 547852 376378 547884 376614
rect 548120 376378 548204 376614
rect 548440 376378 548472 376614
rect 547852 376294 548472 376378
rect 547852 376058 547884 376294
rect 548120 376058 548204 376294
rect 548440 376058 548472 376294
rect 547852 358614 548472 376058
rect 547852 358378 547884 358614
rect 548120 358378 548204 358614
rect 548440 358378 548472 358614
rect 547852 358294 548472 358378
rect 547852 358058 547884 358294
rect 548120 358058 548204 358294
rect 548440 358058 548472 358294
rect 547852 340614 548472 358058
rect 547852 340378 547884 340614
rect 548120 340378 548204 340614
rect 548440 340378 548472 340614
rect 547852 340294 548472 340378
rect 547852 340058 547884 340294
rect 548120 340058 548204 340294
rect 548440 340058 548472 340294
rect 547852 322614 548472 340058
rect 547852 322378 547884 322614
rect 548120 322378 548204 322614
rect 548440 322378 548472 322614
rect 547852 322294 548472 322378
rect 547852 322058 547884 322294
rect 548120 322058 548204 322294
rect 548440 322058 548472 322294
rect 547852 304614 548472 322058
rect 547852 304378 547884 304614
rect 548120 304378 548204 304614
rect 548440 304378 548472 304614
rect 547852 304294 548472 304378
rect 547852 304058 547884 304294
rect 548120 304058 548204 304294
rect 548440 304058 548472 304294
rect 547852 286614 548472 304058
rect 547852 286378 547884 286614
rect 548120 286378 548204 286614
rect 548440 286378 548472 286614
rect 547852 286294 548472 286378
rect 547852 286058 547884 286294
rect 548120 286058 548204 286294
rect 548440 286058 548472 286294
rect 547852 268614 548472 286058
rect 547852 268378 547884 268614
rect 548120 268378 548204 268614
rect 548440 268378 548472 268614
rect 547852 268294 548472 268378
rect 547852 268058 547884 268294
rect 548120 268058 548204 268294
rect 548440 268058 548472 268294
rect 547852 250614 548472 268058
rect 547852 250378 547884 250614
rect 548120 250378 548204 250614
rect 548440 250378 548472 250614
rect 547852 250294 548472 250378
rect 547852 250058 547884 250294
rect 548120 250058 548204 250294
rect 548440 250058 548472 250294
rect 547852 232614 548472 250058
rect 547852 232378 547884 232614
rect 548120 232378 548204 232614
rect 548440 232378 548472 232614
rect 547852 232294 548472 232378
rect 547852 232058 547884 232294
rect 548120 232058 548204 232294
rect 548440 232058 548472 232294
rect 547852 214614 548472 232058
rect 547852 214378 547884 214614
rect 548120 214378 548204 214614
rect 548440 214378 548472 214614
rect 547852 214294 548472 214378
rect 547852 214058 547884 214294
rect 548120 214058 548204 214294
rect 548440 214058 548472 214294
rect 547852 196614 548472 214058
rect 547852 196378 547884 196614
rect 548120 196378 548204 196614
rect 548440 196378 548472 196614
rect 547852 196294 548472 196378
rect 547852 196058 547884 196294
rect 548120 196058 548204 196294
rect 548440 196058 548472 196294
rect 547852 178614 548472 196058
rect 547852 178378 547884 178614
rect 548120 178378 548204 178614
rect 548440 178378 548472 178614
rect 547852 178294 548472 178378
rect 547852 178058 547884 178294
rect 548120 178058 548204 178294
rect 548440 178058 548472 178294
rect 547852 160614 548472 178058
rect 547852 160378 547884 160614
rect 548120 160378 548204 160614
rect 548440 160378 548472 160614
rect 547852 160294 548472 160378
rect 547852 160058 547884 160294
rect 548120 160058 548204 160294
rect 548440 160058 548472 160294
rect 547852 142614 548472 160058
rect 547852 142378 547884 142614
rect 548120 142378 548204 142614
rect 548440 142378 548472 142614
rect 547852 142294 548472 142378
rect 547852 142058 547884 142294
rect 548120 142058 548204 142294
rect 548440 142058 548472 142294
rect 547852 124614 548472 142058
rect 547852 124378 547884 124614
rect 548120 124378 548204 124614
rect 548440 124378 548472 124614
rect 547852 124294 548472 124378
rect 547852 124058 547884 124294
rect 548120 124058 548204 124294
rect 548440 124058 548472 124294
rect 547852 106614 548472 124058
rect 547852 106378 547884 106614
rect 548120 106378 548204 106614
rect 548440 106378 548472 106614
rect 547852 106294 548472 106378
rect 547852 106058 547884 106294
rect 548120 106058 548204 106294
rect 548440 106058 548472 106294
rect 547852 88614 548472 106058
rect 547852 88378 547884 88614
rect 548120 88378 548204 88614
rect 548440 88378 548472 88614
rect 547852 88294 548472 88378
rect 547852 88058 547884 88294
rect 548120 88058 548204 88294
rect 548440 88058 548472 88294
rect 547852 70614 548472 88058
rect 547852 70378 547884 70614
rect 548120 70378 548204 70614
rect 548440 70378 548472 70614
rect 547852 70294 548472 70378
rect 547852 70058 547884 70294
rect 548120 70058 548204 70294
rect 548440 70058 548472 70294
rect 547852 52614 548472 70058
rect 547852 52378 547884 52614
rect 548120 52378 548204 52614
rect 548440 52378 548472 52614
rect 547852 52294 548472 52378
rect 547852 52058 547884 52294
rect 548120 52058 548204 52294
rect 548440 52058 548472 52294
rect 547852 34614 548472 52058
rect 547852 34378 547884 34614
rect 548120 34378 548204 34614
rect 548440 34378 548472 34614
rect 547852 34294 548472 34378
rect 547852 34058 547884 34294
rect 548120 34058 548204 34294
rect 548440 34058 548472 34294
rect 547852 16614 548472 34058
rect 547852 16378 547884 16614
rect 548120 16378 548204 16614
rect 548440 16378 548472 16614
rect 547852 16294 548472 16378
rect 547852 16058 547884 16294
rect 548120 16058 548204 16294
rect 548440 16058 548472 16294
rect 547852 -3736 548472 16058
rect 547852 -3972 547884 -3736
rect 548120 -3972 548204 -3736
rect 548440 -3972 548472 -3736
rect 547852 -4056 548472 -3972
rect 547852 -4292 547884 -4056
rect 548120 -4292 548204 -4056
rect 548440 -4292 548472 -4056
rect 547852 -4324 548472 -4292
<< via4 >>
rect -4444 463736 -4208 463972
rect -4124 463736 -3888 463972
rect -4444 463416 -4208 463652
rect -4124 463416 -3888 463652
rect -4444 448378 -4208 448614
rect -4124 448378 -3888 448614
rect -4444 448058 -4208 448294
rect -4124 448058 -3888 448294
rect -4444 430378 -4208 430614
rect -4124 430378 -3888 430614
rect -4444 430058 -4208 430294
rect -4124 430058 -3888 430294
rect -4444 412378 -4208 412614
rect -4124 412378 -3888 412614
rect -4444 412058 -4208 412294
rect -4124 412058 -3888 412294
rect -4444 394378 -4208 394614
rect -4124 394378 -3888 394614
rect -4444 394058 -4208 394294
rect -4124 394058 -3888 394294
rect -4444 376378 -4208 376614
rect -4124 376378 -3888 376614
rect -4444 376058 -4208 376294
rect -4124 376058 -3888 376294
rect -4444 358378 -4208 358614
rect -4124 358378 -3888 358614
rect -4444 358058 -4208 358294
rect -4124 358058 -3888 358294
rect -4444 340378 -4208 340614
rect -4124 340378 -3888 340614
rect -4444 340058 -4208 340294
rect -4124 340058 -3888 340294
rect -4444 322378 -4208 322614
rect -4124 322378 -3888 322614
rect -4444 322058 -4208 322294
rect -4124 322058 -3888 322294
rect -4444 304378 -4208 304614
rect -4124 304378 -3888 304614
rect -4444 304058 -4208 304294
rect -4124 304058 -3888 304294
rect -4444 286378 -4208 286614
rect -4124 286378 -3888 286614
rect -4444 286058 -4208 286294
rect -4124 286058 -3888 286294
rect -4444 268378 -4208 268614
rect -4124 268378 -3888 268614
rect -4444 268058 -4208 268294
rect -4124 268058 -3888 268294
rect -4444 250378 -4208 250614
rect -4124 250378 -3888 250614
rect -4444 250058 -4208 250294
rect -4124 250058 -3888 250294
rect -4444 232378 -4208 232614
rect -4124 232378 -3888 232614
rect -4444 232058 -4208 232294
rect -4124 232058 -3888 232294
rect -4444 214378 -4208 214614
rect -4124 214378 -3888 214614
rect -4444 214058 -4208 214294
rect -4124 214058 -3888 214294
rect -4444 196378 -4208 196614
rect -4124 196378 -3888 196614
rect -4444 196058 -4208 196294
rect -4124 196058 -3888 196294
rect -4444 178378 -4208 178614
rect -4124 178378 -3888 178614
rect -4444 178058 -4208 178294
rect -4124 178058 -3888 178294
rect -4444 160378 -4208 160614
rect -4124 160378 -3888 160614
rect -4444 160058 -4208 160294
rect -4124 160058 -3888 160294
rect -4444 142378 -4208 142614
rect -4124 142378 -3888 142614
rect -4444 142058 -4208 142294
rect -4124 142058 -3888 142294
rect -4444 124378 -4208 124614
rect -4124 124378 -3888 124614
rect -4444 124058 -4208 124294
rect -4124 124058 -3888 124294
rect -4444 106378 -4208 106614
rect -4124 106378 -3888 106614
rect -4444 106058 -4208 106294
rect -4124 106058 -3888 106294
rect -4444 88378 -4208 88614
rect -4124 88378 -3888 88614
rect -4444 88058 -4208 88294
rect -4124 88058 -3888 88294
rect -4444 70378 -4208 70614
rect -4124 70378 -3888 70614
rect -4444 70058 -4208 70294
rect -4124 70058 -3888 70294
rect -4444 52378 -4208 52614
rect -4124 52378 -3888 52614
rect -4444 52058 -4208 52294
rect -4124 52058 -3888 52294
rect -4444 34378 -4208 34614
rect -4124 34378 -3888 34614
rect -4444 34058 -4208 34294
rect -4124 34058 -3888 34294
rect -4444 16378 -4208 16614
rect -4124 16378 -3888 16614
rect -4444 16058 -4208 16294
rect -4124 16058 -3888 16294
rect -3484 462776 -3248 463012
rect -3164 462776 -2928 463012
rect -3484 462456 -3248 462692
rect -3164 462456 -2928 462692
rect -3484 444658 -3248 444894
rect -3164 444658 -2928 444894
rect -3484 444338 -3248 444574
rect -3164 444338 -2928 444574
rect -3484 426658 -3248 426894
rect -3164 426658 -2928 426894
rect -3484 426338 -3248 426574
rect -3164 426338 -2928 426574
rect -3484 408658 -3248 408894
rect -3164 408658 -2928 408894
rect -3484 408338 -3248 408574
rect -3164 408338 -2928 408574
rect -3484 390658 -3248 390894
rect -3164 390658 -2928 390894
rect -3484 390338 -3248 390574
rect -3164 390338 -2928 390574
rect -3484 372658 -3248 372894
rect -3164 372658 -2928 372894
rect -3484 372338 -3248 372574
rect -3164 372338 -2928 372574
rect -3484 354658 -3248 354894
rect -3164 354658 -2928 354894
rect -3484 354338 -3248 354574
rect -3164 354338 -2928 354574
rect -3484 336658 -3248 336894
rect -3164 336658 -2928 336894
rect -3484 336338 -3248 336574
rect -3164 336338 -2928 336574
rect -3484 318658 -3248 318894
rect -3164 318658 -2928 318894
rect -3484 318338 -3248 318574
rect -3164 318338 -2928 318574
rect -3484 300658 -3248 300894
rect -3164 300658 -2928 300894
rect -3484 300338 -3248 300574
rect -3164 300338 -2928 300574
rect -3484 282658 -3248 282894
rect -3164 282658 -2928 282894
rect -3484 282338 -3248 282574
rect -3164 282338 -2928 282574
rect -3484 264658 -3248 264894
rect -3164 264658 -2928 264894
rect -3484 264338 -3248 264574
rect -3164 264338 -2928 264574
rect -3484 246658 -3248 246894
rect -3164 246658 -2928 246894
rect -3484 246338 -3248 246574
rect -3164 246338 -2928 246574
rect -3484 228658 -3248 228894
rect -3164 228658 -2928 228894
rect -3484 228338 -3248 228574
rect -3164 228338 -2928 228574
rect -3484 210658 -3248 210894
rect -3164 210658 -2928 210894
rect -3484 210338 -3248 210574
rect -3164 210338 -2928 210574
rect -3484 192658 -3248 192894
rect -3164 192658 -2928 192894
rect -3484 192338 -3248 192574
rect -3164 192338 -2928 192574
rect -3484 174658 -3248 174894
rect -3164 174658 -2928 174894
rect -3484 174338 -3248 174574
rect -3164 174338 -2928 174574
rect -3484 156658 -3248 156894
rect -3164 156658 -2928 156894
rect -3484 156338 -3248 156574
rect -3164 156338 -2928 156574
rect -3484 138658 -3248 138894
rect -3164 138658 -2928 138894
rect -3484 138338 -3248 138574
rect -3164 138338 -2928 138574
rect -3484 120658 -3248 120894
rect -3164 120658 -2928 120894
rect -3484 120338 -3248 120574
rect -3164 120338 -2928 120574
rect -3484 102658 -3248 102894
rect -3164 102658 -2928 102894
rect -3484 102338 -3248 102574
rect -3164 102338 -2928 102574
rect -3484 84658 -3248 84894
rect -3164 84658 -2928 84894
rect -3484 84338 -3248 84574
rect -3164 84338 -2928 84574
rect -3484 66658 -3248 66894
rect -3164 66658 -2928 66894
rect -3484 66338 -3248 66574
rect -3164 66338 -2928 66574
rect -3484 48658 -3248 48894
rect -3164 48658 -2928 48894
rect -3484 48338 -3248 48574
rect -3164 48338 -2928 48574
rect -3484 30658 -3248 30894
rect -3164 30658 -2928 30894
rect -3484 30338 -3248 30574
rect -3164 30338 -2928 30574
rect -3484 12658 -3248 12894
rect -3164 12658 -2928 12894
rect -3484 12338 -3248 12574
rect -3164 12338 -2928 12574
rect -2524 461816 -2288 462052
rect -2204 461816 -1968 462052
rect -2524 461496 -2288 461732
rect -2204 461496 -1968 461732
rect -2524 440938 -2288 441174
rect -2204 440938 -1968 441174
rect -2524 440618 -2288 440854
rect -2204 440618 -1968 440854
rect -2524 422938 -2288 423174
rect -2204 422938 -1968 423174
rect -2524 422618 -2288 422854
rect -2204 422618 -1968 422854
rect -2524 404938 -2288 405174
rect -2204 404938 -1968 405174
rect -2524 404618 -2288 404854
rect -2204 404618 -1968 404854
rect -2524 386938 -2288 387174
rect -2204 386938 -1968 387174
rect -2524 386618 -2288 386854
rect -2204 386618 -1968 386854
rect -2524 368938 -2288 369174
rect -2204 368938 -1968 369174
rect -2524 368618 -2288 368854
rect -2204 368618 -1968 368854
rect -2524 350938 -2288 351174
rect -2204 350938 -1968 351174
rect -2524 350618 -2288 350854
rect -2204 350618 -1968 350854
rect -2524 332938 -2288 333174
rect -2204 332938 -1968 333174
rect -2524 332618 -2288 332854
rect -2204 332618 -1968 332854
rect -2524 314938 -2288 315174
rect -2204 314938 -1968 315174
rect -2524 314618 -2288 314854
rect -2204 314618 -1968 314854
rect -2524 296938 -2288 297174
rect -2204 296938 -1968 297174
rect -2524 296618 -2288 296854
rect -2204 296618 -1968 296854
rect -2524 278938 -2288 279174
rect -2204 278938 -1968 279174
rect -2524 278618 -2288 278854
rect -2204 278618 -1968 278854
rect -2524 260938 -2288 261174
rect -2204 260938 -1968 261174
rect -2524 260618 -2288 260854
rect -2204 260618 -1968 260854
rect -2524 242938 -2288 243174
rect -2204 242938 -1968 243174
rect -2524 242618 -2288 242854
rect -2204 242618 -1968 242854
rect -2524 224938 -2288 225174
rect -2204 224938 -1968 225174
rect -2524 224618 -2288 224854
rect -2204 224618 -1968 224854
rect -2524 206938 -2288 207174
rect -2204 206938 -1968 207174
rect -2524 206618 -2288 206854
rect -2204 206618 -1968 206854
rect -2524 188938 -2288 189174
rect -2204 188938 -1968 189174
rect -2524 188618 -2288 188854
rect -2204 188618 -1968 188854
rect -2524 170938 -2288 171174
rect -2204 170938 -1968 171174
rect -2524 170618 -2288 170854
rect -2204 170618 -1968 170854
rect -2524 152938 -2288 153174
rect -2204 152938 -1968 153174
rect -2524 152618 -2288 152854
rect -2204 152618 -1968 152854
rect -2524 134938 -2288 135174
rect -2204 134938 -1968 135174
rect -2524 134618 -2288 134854
rect -2204 134618 -1968 134854
rect -2524 116938 -2288 117174
rect -2204 116938 -1968 117174
rect -2524 116618 -2288 116854
rect -2204 116618 -1968 116854
rect -2524 98938 -2288 99174
rect -2204 98938 -1968 99174
rect -2524 98618 -2288 98854
rect -2204 98618 -1968 98854
rect -2524 80938 -2288 81174
rect -2204 80938 -1968 81174
rect -2524 80618 -2288 80854
rect -2204 80618 -1968 80854
rect -2524 62938 -2288 63174
rect -2204 62938 -1968 63174
rect -2524 62618 -2288 62854
rect -2204 62618 -1968 62854
rect -2524 44938 -2288 45174
rect -2204 44938 -1968 45174
rect -2524 44618 -2288 44854
rect -2204 44618 -1968 44854
rect -2524 26938 -2288 27174
rect -2204 26938 -1968 27174
rect -2524 26618 -2288 26854
rect -2204 26618 -1968 26854
rect -2524 8938 -2288 9174
rect -2204 8938 -1968 9174
rect -2524 8618 -2288 8854
rect -2204 8618 -1968 8854
rect -1564 460856 -1328 461092
rect -1244 460856 -1008 461092
rect -1564 460536 -1328 460772
rect -1244 460536 -1008 460772
rect -1564 455218 -1328 455454
rect -1244 455218 -1008 455454
rect -1564 454898 -1328 455134
rect -1244 454898 -1008 455134
rect -1564 437218 -1328 437454
rect -1244 437218 -1008 437454
rect -1564 436898 -1328 437134
rect -1244 436898 -1008 437134
rect -1564 419218 -1328 419454
rect -1244 419218 -1008 419454
rect -1564 418898 -1328 419134
rect -1244 418898 -1008 419134
rect -1564 401218 -1328 401454
rect -1244 401218 -1008 401454
rect -1564 400898 -1328 401134
rect -1244 400898 -1008 401134
rect -1564 383218 -1328 383454
rect -1244 383218 -1008 383454
rect -1564 382898 -1328 383134
rect -1244 382898 -1008 383134
rect -1564 365218 -1328 365454
rect -1244 365218 -1008 365454
rect -1564 364898 -1328 365134
rect -1244 364898 -1008 365134
rect -1564 347218 -1328 347454
rect -1244 347218 -1008 347454
rect -1564 346898 -1328 347134
rect -1244 346898 -1008 347134
rect -1564 329218 -1328 329454
rect -1244 329218 -1008 329454
rect -1564 328898 -1328 329134
rect -1244 328898 -1008 329134
rect -1564 311218 -1328 311454
rect -1244 311218 -1008 311454
rect -1564 310898 -1328 311134
rect -1244 310898 -1008 311134
rect -1564 293218 -1328 293454
rect -1244 293218 -1008 293454
rect -1564 292898 -1328 293134
rect -1244 292898 -1008 293134
rect 4746 460856 4982 461092
rect 5066 460856 5302 461092
rect 4746 460536 4982 460772
rect 5066 460536 5302 460772
rect 4746 455218 4982 455454
rect 5066 455218 5302 455454
rect 4746 454898 4982 455134
rect 5066 454898 5302 455134
rect 4746 437218 4982 437454
rect 5066 437218 5302 437454
rect 4746 436898 4982 437134
rect 5066 436898 5302 437134
rect 4746 419218 4982 419454
rect 5066 419218 5302 419454
rect 4746 418898 4982 419134
rect 5066 418898 5302 419134
rect 4746 401218 4982 401454
rect 5066 401218 5302 401454
rect 4746 400898 4982 401134
rect 5066 400898 5302 401134
rect 4746 383218 4982 383454
rect 5066 383218 5302 383454
rect 4746 382898 4982 383134
rect 5066 382898 5302 383134
rect 4746 365218 4982 365454
rect 5066 365218 5302 365454
rect 4746 364898 4982 365134
rect 5066 364898 5302 365134
rect 4746 347218 4982 347454
rect 5066 347218 5302 347454
rect 4746 346898 4982 347134
rect 5066 346898 5302 347134
rect 4746 329218 4982 329454
rect 5066 329218 5302 329454
rect 4746 328898 4982 329134
rect 5066 328898 5302 329134
rect 4746 311218 4982 311454
rect 5066 311218 5302 311454
rect 4746 310898 4982 311134
rect 5066 310898 5302 311134
rect 4746 293218 4982 293454
rect 5066 293218 5302 293454
rect 4746 292898 4982 293134
rect 5066 292898 5302 293134
rect -1564 275218 -1328 275454
rect -1244 275218 -1008 275454
rect -1564 274898 -1328 275134
rect -1244 274898 -1008 275134
rect -1564 257218 -1328 257454
rect -1244 257218 -1008 257454
rect -1564 256898 -1328 257134
rect -1244 256898 -1008 257134
rect -1564 239218 -1328 239454
rect -1244 239218 -1008 239454
rect -1564 238898 -1328 239134
rect -1244 238898 -1008 239134
rect -1564 221218 -1328 221454
rect -1244 221218 -1008 221454
rect -1564 220898 -1328 221134
rect -1244 220898 -1008 221134
rect -1564 203218 -1328 203454
rect -1244 203218 -1008 203454
rect -1564 202898 -1328 203134
rect -1244 202898 -1008 203134
rect -1564 185218 -1328 185454
rect -1244 185218 -1008 185454
rect -1564 184898 -1328 185134
rect -1244 184898 -1008 185134
rect -1564 167218 -1328 167454
rect -1244 167218 -1008 167454
rect -1564 166898 -1328 167134
rect -1244 166898 -1008 167134
rect -1564 149218 -1328 149454
rect -1244 149218 -1008 149454
rect -1564 148898 -1328 149134
rect -1244 148898 -1008 149134
rect -1564 131218 -1328 131454
rect -1244 131218 -1008 131454
rect -1564 130898 -1328 131134
rect -1244 130898 -1008 131134
rect -1564 113218 -1328 113454
rect -1244 113218 -1008 113454
rect -1564 112898 -1328 113134
rect -1244 112898 -1008 113134
rect -1564 95218 -1328 95454
rect -1244 95218 -1008 95454
rect -1564 94898 -1328 95134
rect -1244 94898 -1008 95134
rect -1564 77218 -1328 77454
rect -1244 77218 -1008 77454
rect -1564 76898 -1328 77134
rect -1244 76898 -1008 77134
rect 4746 275218 4982 275454
rect 5066 275218 5302 275454
rect 4746 274898 4982 275134
rect 5066 274898 5302 275134
rect 4746 257218 4982 257454
rect 5066 257218 5302 257454
rect 4746 256898 4982 257134
rect 5066 256898 5302 257134
rect 4746 239218 4982 239454
rect 5066 239218 5302 239454
rect 4746 238898 4982 239134
rect 5066 238898 5302 239134
rect 4746 221218 4982 221454
rect 5066 221218 5302 221454
rect 4746 220898 4982 221134
rect 5066 220898 5302 221134
rect 4746 203218 4982 203454
rect 5066 203218 5302 203454
rect 4746 202898 4982 203134
rect 5066 202898 5302 203134
rect 4746 185218 4982 185454
rect 5066 185218 5302 185454
rect 4746 184898 4982 185134
rect 5066 184898 5302 185134
rect 4746 167218 4982 167454
rect 5066 167218 5302 167454
rect 4746 166898 4982 167134
rect 5066 166898 5302 167134
rect 4746 149218 4982 149454
rect 5066 149218 5302 149454
rect 4746 148898 4982 149134
rect 5066 148898 5302 149134
rect 4746 131218 4982 131454
rect 5066 131218 5302 131454
rect 4746 130898 4982 131134
rect 5066 130898 5302 131134
rect 4746 113218 4982 113454
rect 5066 113218 5302 113454
rect 4746 112898 4982 113134
rect 5066 112898 5302 113134
rect 4746 95218 4982 95454
rect 5066 95218 5302 95454
rect 4746 94898 4982 95134
rect 5066 94898 5302 95134
rect 4746 77218 4982 77454
rect 5066 77218 5302 77454
rect 4746 76898 4982 77134
rect 5066 76898 5302 77134
rect 158 60062 394 60298
rect -1564 59218 -1328 59454
rect -1244 59218 -1008 59454
rect -1564 58898 -1328 59134
rect -1244 58898 -1008 59134
rect -1564 41218 -1328 41454
rect -1244 41218 -1008 41454
rect -1564 40898 -1328 41134
rect -1244 40898 -1008 41134
rect -1564 23218 -1328 23454
rect -1244 23218 -1008 23454
rect -1564 22898 -1328 23134
rect -1244 22898 -1008 23134
rect -1564 5218 -1328 5454
rect -1244 5218 -1008 5454
rect -1564 4898 -1328 5134
rect -1244 4898 -1008 5134
rect 4746 59218 4982 59454
rect 5066 59218 5302 59454
rect 4746 58898 4982 59134
rect 5066 58898 5302 59134
rect 4746 41218 4982 41454
rect 5066 41218 5302 41454
rect 4746 40898 4982 41134
rect 5066 40898 5302 41134
rect 4746 23218 4982 23454
rect 5066 23218 5302 23454
rect 4746 22898 4982 23134
rect 5066 22898 5302 23134
rect 4746 5218 4982 5454
rect 5066 5218 5302 5454
rect 4746 4898 4982 5134
rect 5066 4898 5302 5134
rect 8466 461816 8702 462052
rect 8786 461816 9022 462052
rect 8466 461496 8702 461732
rect 8786 461496 9022 461732
rect 8466 440938 8702 441174
rect 8786 440938 9022 441174
rect 8466 440618 8702 440854
rect 8786 440618 9022 440854
rect 8466 422938 8702 423174
rect 8786 422938 9022 423174
rect 8466 422618 8702 422854
rect 8786 422618 9022 422854
rect 8466 404938 8702 405174
rect 8786 404938 9022 405174
rect 8466 404618 8702 404854
rect 8786 404618 9022 404854
rect 8466 386938 8702 387174
rect 8786 386938 9022 387174
rect 8466 386618 8702 386854
rect 8786 386618 9022 386854
rect 8466 368938 8702 369174
rect 8786 368938 9022 369174
rect 8466 368618 8702 368854
rect 8786 368618 9022 368854
rect 8466 350938 8702 351174
rect 8786 350938 9022 351174
rect 8466 350618 8702 350854
rect 8786 350618 9022 350854
rect 8466 332938 8702 333174
rect 8786 332938 9022 333174
rect 8466 332618 8702 332854
rect 8786 332618 9022 332854
rect 8466 314938 8702 315174
rect 8786 314938 9022 315174
rect 8466 314618 8702 314854
rect 8786 314618 9022 314854
rect 8466 296938 8702 297174
rect 8786 296938 9022 297174
rect 8466 296618 8702 296854
rect 8786 296618 9022 296854
rect 8466 278938 8702 279174
rect 8786 278938 9022 279174
rect 8466 278618 8702 278854
rect 8786 278618 9022 278854
rect 8466 260938 8702 261174
rect 8786 260938 9022 261174
rect 8466 260618 8702 260854
rect 8786 260618 9022 260854
rect 8466 242938 8702 243174
rect 8786 242938 9022 243174
rect 8466 242618 8702 242854
rect 8786 242618 9022 242854
rect 8466 224938 8702 225174
rect 8786 224938 9022 225174
rect 8466 224618 8702 224854
rect 8786 224618 9022 224854
rect 8466 206938 8702 207174
rect 8786 206938 9022 207174
rect 8466 206618 8702 206854
rect 8786 206618 9022 206854
rect 8466 188938 8702 189174
rect 8786 188938 9022 189174
rect 8466 188618 8702 188854
rect 8786 188618 9022 188854
rect 8466 170938 8702 171174
rect 8786 170938 9022 171174
rect 8466 170618 8702 170854
rect 8786 170618 9022 170854
rect 8466 152938 8702 153174
rect 8786 152938 9022 153174
rect 8466 152618 8702 152854
rect 8786 152618 9022 152854
rect 8466 134938 8702 135174
rect 8786 134938 9022 135174
rect 8466 134618 8702 134854
rect 8786 134618 9022 134854
rect 8466 116938 8702 117174
rect 8786 116938 9022 117174
rect 8466 116618 8702 116854
rect 8786 116618 9022 116854
rect 8466 98938 8702 99174
rect 8786 98938 9022 99174
rect 8466 98618 8702 98854
rect 8786 98618 9022 98854
rect 8466 80938 8702 81174
rect 8786 80938 9022 81174
rect 8466 80618 8702 80854
rect 8786 80618 9022 80854
rect 8466 62938 8702 63174
rect 8786 62938 9022 63174
rect 8466 62618 8702 62854
rect 8786 62618 9022 62854
rect 8466 44938 8702 45174
rect 8786 44938 9022 45174
rect 8466 44618 8702 44854
rect 8786 44618 9022 44854
rect 8466 26938 8702 27174
rect 8786 26938 9022 27174
rect 8466 26618 8702 26854
rect 8786 26618 9022 26854
rect 8466 8938 8702 9174
rect 8786 8938 9022 9174
rect 8466 8618 8702 8854
rect 8786 8618 9022 8854
rect 12186 462776 12422 463012
rect 12506 462776 12742 463012
rect 12186 462456 12422 462692
rect 12506 462456 12742 462692
rect 12186 444658 12422 444894
rect 12506 444658 12742 444894
rect 12186 444338 12422 444574
rect 12506 444338 12742 444574
rect 12186 426658 12422 426894
rect 12506 426658 12742 426894
rect 12186 426338 12422 426574
rect 12506 426338 12742 426574
rect 12186 408658 12422 408894
rect 12506 408658 12742 408894
rect 12186 408338 12422 408574
rect 12506 408338 12742 408574
rect 12186 390658 12422 390894
rect 12506 390658 12742 390894
rect 12186 390338 12422 390574
rect 12506 390338 12742 390574
rect 12186 372658 12422 372894
rect 12506 372658 12742 372894
rect 12186 372338 12422 372574
rect 12506 372338 12742 372574
rect 12186 354658 12422 354894
rect 12506 354658 12742 354894
rect 12186 354338 12422 354574
rect 12506 354338 12742 354574
rect 12186 336658 12422 336894
rect 12506 336658 12742 336894
rect 12186 336338 12422 336574
rect 12506 336338 12742 336574
rect 12186 318658 12422 318894
rect 12506 318658 12742 318894
rect 12186 318338 12422 318574
rect 12506 318338 12742 318574
rect 12186 300658 12422 300894
rect 12506 300658 12742 300894
rect 12186 300338 12422 300574
rect 12506 300338 12742 300574
rect 12186 282658 12422 282894
rect 12506 282658 12742 282894
rect 12186 282338 12422 282574
rect 12506 282338 12742 282574
rect 12186 264658 12422 264894
rect 12506 264658 12742 264894
rect 12186 264338 12422 264574
rect 12506 264338 12742 264574
rect 12186 246658 12422 246894
rect 12506 246658 12742 246894
rect 12186 246338 12422 246574
rect 12506 246338 12742 246574
rect 12186 228658 12422 228894
rect 12506 228658 12742 228894
rect 12186 228338 12422 228574
rect 12506 228338 12742 228574
rect 12186 210658 12422 210894
rect 12506 210658 12742 210894
rect 12186 210338 12422 210574
rect 12506 210338 12742 210574
rect 12186 192658 12422 192894
rect 12506 192658 12742 192894
rect 12186 192338 12422 192574
rect 12506 192338 12742 192574
rect 12186 174658 12422 174894
rect 12506 174658 12742 174894
rect 12186 174338 12422 174574
rect 12506 174338 12742 174574
rect 12186 156658 12422 156894
rect 12506 156658 12742 156894
rect 12186 156338 12422 156574
rect 12506 156338 12742 156574
rect 12186 138658 12422 138894
rect 12506 138658 12742 138894
rect 12186 138338 12422 138574
rect 12506 138338 12742 138574
rect 12186 120658 12422 120894
rect 12506 120658 12742 120894
rect 12186 120338 12422 120574
rect 12506 120338 12742 120574
rect 12186 102658 12422 102894
rect 12506 102658 12742 102894
rect 12186 102338 12422 102574
rect 12506 102338 12742 102574
rect 12186 84658 12422 84894
rect 12506 84658 12742 84894
rect 12186 84338 12422 84574
rect 12506 84338 12742 84574
rect 12186 66658 12422 66894
rect 12506 66658 12742 66894
rect 12186 66338 12422 66574
rect 12506 66338 12742 66574
rect 12186 48658 12422 48894
rect 12506 48658 12742 48894
rect 12186 48338 12422 48574
rect 12506 48338 12742 48574
rect 12186 30658 12422 30894
rect 12506 30658 12742 30894
rect 12186 30338 12422 30574
rect 12506 30338 12742 30574
rect 12186 12658 12422 12894
rect 12506 12658 12742 12894
rect 12186 12338 12422 12574
rect 12506 12338 12742 12574
rect 15906 463736 16142 463972
rect 16226 463736 16462 463972
rect 15906 463416 16142 463652
rect 16226 463416 16462 463652
rect 15906 448378 16142 448614
rect 16226 448378 16462 448614
rect 15906 448058 16142 448294
rect 16226 448058 16462 448294
rect 15906 430378 16142 430614
rect 16226 430378 16462 430614
rect 15906 430058 16142 430294
rect 16226 430058 16462 430294
rect 15906 412378 16142 412614
rect 16226 412378 16462 412614
rect 15906 412058 16142 412294
rect 16226 412058 16462 412294
rect 15906 394378 16142 394614
rect 16226 394378 16462 394614
rect 15906 394058 16142 394294
rect 16226 394058 16462 394294
rect 15906 376378 16142 376614
rect 16226 376378 16462 376614
rect 15906 376058 16142 376294
rect 16226 376058 16462 376294
rect 15906 358378 16142 358614
rect 16226 358378 16462 358614
rect 15906 358058 16142 358294
rect 16226 358058 16462 358294
rect 15906 340378 16142 340614
rect 16226 340378 16462 340614
rect 15906 340058 16142 340294
rect 16226 340058 16462 340294
rect 15906 322378 16142 322614
rect 16226 322378 16462 322614
rect 15906 322058 16142 322294
rect 16226 322058 16462 322294
rect 15906 304378 16142 304614
rect 16226 304378 16462 304614
rect 15906 304058 16142 304294
rect 16226 304058 16462 304294
rect 15906 286378 16142 286614
rect 16226 286378 16462 286614
rect 15906 286058 16142 286294
rect 16226 286058 16462 286294
rect 15906 268378 16142 268614
rect 16226 268378 16462 268614
rect 15906 268058 16142 268294
rect 16226 268058 16462 268294
rect 15906 250378 16142 250614
rect 16226 250378 16462 250614
rect 15906 250058 16142 250294
rect 16226 250058 16462 250294
rect 15906 232378 16142 232614
rect 16226 232378 16462 232614
rect 15906 232058 16142 232294
rect 16226 232058 16462 232294
rect 15906 214378 16142 214614
rect 16226 214378 16462 214614
rect 15906 214058 16142 214294
rect 16226 214058 16462 214294
rect 15906 196378 16142 196614
rect 16226 196378 16462 196614
rect 15906 196058 16142 196294
rect 16226 196058 16462 196294
rect 15906 178378 16142 178614
rect 16226 178378 16462 178614
rect 15906 178058 16142 178294
rect 16226 178058 16462 178294
rect 15906 160378 16142 160614
rect 16226 160378 16462 160614
rect 15906 160058 16142 160294
rect 16226 160058 16462 160294
rect 15906 142378 16142 142614
rect 16226 142378 16462 142614
rect 15906 142058 16142 142294
rect 16226 142058 16462 142294
rect 15906 124378 16142 124614
rect 16226 124378 16462 124614
rect 15906 124058 16142 124294
rect 16226 124058 16462 124294
rect 15906 106378 16142 106614
rect 16226 106378 16462 106614
rect 15906 106058 16142 106294
rect 16226 106058 16462 106294
rect 15906 88378 16142 88614
rect 16226 88378 16462 88614
rect 15906 88058 16142 88294
rect 16226 88058 16462 88294
rect 15906 70378 16142 70614
rect 16226 70378 16462 70614
rect 15906 70058 16142 70294
rect 16226 70058 16462 70294
rect 15906 52378 16142 52614
rect 16226 52378 16462 52614
rect 15906 52058 16142 52294
rect 16226 52058 16462 52294
rect 15906 34378 16142 34614
rect 16226 34378 16462 34614
rect 15906 34058 16142 34294
rect 16226 34058 16462 34294
rect 15906 16378 16142 16614
rect 16226 16378 16462 16614
rect 15906 16058 16142 16294
rect 16226 16058 16462 16294
rect 22746 460856 22982 461092
rect 23066 460856 23302 461092
rect 22746 460536 22982 460772
rect 23066 460536 23302 460772
rect 22746 455218 22982 455454
rect 23066 455218 23302 455454
rect 22746 454898 22982 455134
rect 23066 454898 23302 455134
rect 22746 437218 22982 437454
rect 23066 437218 23302 437454
rect 22746 436898 22982 437134
rect 23066 436898 23302 437134
rect 22746 419218 22982 419454
rect 23066 419218 23302 419454
rect 22746 418898 22982 419134
rect 23066 418898 23302 419134
rect 22746 401218 22982 401454
rect 23066 401218 23302 401454
rect 22746 400898 22982 401134
rect 23066 400898 23302 401134
rect 22746 383218 22982 383454
rect 23066 383218 23302 383454
rect 22746 382898 22982 383134
rect 23066 382898 23302 383134
rect 22746 365218 22982 365454
rect 23066 365218 23302 365454
rect 22746 364898 22982 365134
rect 23066 364898 23302 365134
rect 22746 347218 22982 347454
rect 23066 347218 23302 347454
rect 22746 346898 22982 347134
rect 23066 346898 23302 347134
rect 22746 329218 22982 329454
rect 23066 329218 23302 329454
rect 22746 328898 22982 329134
rect 23066 328898 23302 329134
rect 22746 311218 22982 311454
rect 23066 311218 23302 311454
rect 22746 310898 22982 311134
rect 23066 310898 23302 311134
rect 22746 293218 22982 293454
rect 23066 293218 23302 293454
rect 22746 292898 22982 293134
rect 23066 292898 23302 293134
rect 22746 275218 22982 275454
rect 23066 275218 23302 275454
rect 22746 274898 22982 275134
rect 23066 274898 23302 275134
rect 22746 257218 22982 257454
rect 23066 257218 23302 257454
rect 22746 256898 22982 257134
rect 23066 256898 23302 257134
rect 22746 239218 22982 239454
rect 23066 239218 23302 239454
rect 22746 238898 22982 239134
rect 23066 238898 23302 239134
rect 22746 221218 22982 221454
rect 23066 221218 23302 221454
rect 22746 220898 22982 221134
rect 23066 220898 23302 221134
rect 22746 203218 22982 203454
rect 23066 203218 23302 203454
rect 22746 202898 22982 203134
rect 23066 202898 23302 203134
rect 22746 185218 22982 185454
rect 23066 185218 23302 185454
rect 22746 184898 22982 185134
rect 23066 184898 23302 185134
rect 22746 167218 22982 167454
rect 23066 167218 23302 167454
rect 22746 166898 22982 167134
rect 23066 166898 23302 167134
rect 22746 149218 22982 149454
rect 23066 149218 23302 149454
rect 22746 148898 22982 149134
rect 23066 148898 23302 149134
rect 22746 131218 22982 131454
rect 23066 131218 23302 131454
rect 22746 130898 22982 131134
rect 23066 130898 23302 131134
rect 22746 113218 22982 113454
rect 23066 113218 23302 113454
rect 22746 112898 22982 113134
rect 23066 112898 23302 113134
rect 22746 95218 22982 95454
rect 23066 95218 23302 95454
rect 22746 94898 22982 95134
rect 23066 94898 23302 95134
rect 22746 77218 22982 77454
rect 23066 77218 23302 77454
rect 22746 76898 22982 77134
rect 23066 76898 23302 77134
rect 22746 59218 22982 59454
rect 23066 59218 23302 59454
rect 22746 58898 22982 59134
rect 23066 58898 23302 59134
rect 22746 41218 22982 41454
rect 23066 41218 23302 41454
rect 22746 40898 22982 41134
rect 23066 40898 23302 41134
rect 22746 23218 22982 23454
rect 23066 23218 23302 23454
rect 22746 22898 22982 23134
rect 23066 22898 23302 23134
rect 22746 5218 22982 5454
rect 23066 5218 23302 5454
rect 22746 4898 22982 5134
rect 23066 4898 23302 5134
rect 26466 461816 26702 462052
rect 26786 461816 27022 462052
rect 26466 461496 26702 461732
rect 26786 461496 27022 461732
rect 26466 440938 26702 441174
rect 26786 440938 27022 441174
rect 26466 440618 26702 440854
rect 26786 440618 27022 440854
rect 26466 422938 26702 423174
rect 26786 422938 27022 423174
rect 26466 422618 26702 422854
rect 26786 422618 27022 422854
rect 26466 404938 26702 405174
rect 26786 404938 27022 405174
rect 26466 404618 26702 404854
rect 26786 404618 27022 404854
rect 26466 386938 26702 387174
rect 26786 386938 27022 387174
rect 26466 386618 26702 386854
rect 26786 386618 27022 386854
rect 26466 368938 26702 369174
rect 26786 368938 27022 369174
rect 26466 368618 26702 368854
rect 26786 368618 27022 368854
rect 26466 350938 26702 351174
rect 26786 350938 27022 351174
rect 26466 350618 26702 350854
rect 26786 350618 27022 350854
rect 26466 332938 26702 333174
rect 26786 332938 27022 333174
rect 26466 332618 26702 332854
rect 26786 332618 27022 332854
rect 26466 314938 26702 315174
rect 26786 314938 27022 315174
rect 26466 314618 26702 314854
rect 26786 314618 27022 314854
rect 26466 296938 26702 297174
rect 26786 296938 27022 297174
rect 26466 296618 26702 296854
rect 26786 296618 27022 296854
rect 26466 278938 26702 279174
rect 26786 278938 27022 279174
rect 26466 278618 26702 278854
rect 26786 278618 27022 278854
rect 26466 260938 26702 261174
rect 26786 260938 27022 261174
rect 26466 260618 26702 260854
rect 26786 260618 27022 260854
rect 26466 242938 26702 243174
rect 26786 242938 27022 243174
rect 26466 242618 26702 242854
rect 26786 242618 27022 242854
rect 26466 224938 26702 225174
rect 26786 224938 27022 225174
rect 26466 224618 26702 224854
rect 26786 224618 27022 224854
rect 26466 206938 26702 207174
rect 26786 206938 27022 207174
rect 26466 206618 26702 206854
rect 26786 206618 27022 206854
rect 26466 188938 26702 189174
rect 26786 188938 27022 189174
rect 26466 188618 26702 188854
rect 26786 188618 27022 188854
rect 26466 170938 26702 171174
rect 26786 170938 27022 171174
rect 26466 170618 26702 170854
rect 26786 170618 27022 170854
rect 26466 152938 26702 153174
rect 26786 152938 27022 153174
rect 26466 152618 26702 152854
rect 26786 152618 27022 152854
rect 26466 134938 26702 135174
rect 26786 134938 27022 135174
rect 26466 134618 26702 134854
rect 26786 134618 27022 134854
rect 26466 116938 26702 117174
rect 26786 116938 27022 117174
rect 26466 116618 26702 116854
rect 26786 116618 27022 116854
rect 26466 98938 26702 99174
rect 26786 98938 27022 99174
rect 26466 98618 26702 98854
rect 26786 98618 27022 98854
rect 26466 80938 26702 81174
rect 26786 80938 27022 81174
rect 26466 80618 26702 80854
rect 26786 80618 27022 80854
rect 26466 62938 26702 63174
rect 26786 62938 27022 63174
rect 26466 62618 26702 62854
rect 26786 62618 27022 62854
rect 26466 44938 26702 45174
rect 26786 44938 27022 45174
rect 26466 44618 26702 44854
rect 26786 44618 27022 44854
rect 26466 26938 26702 27174
rect 26786 26938 27022 27174
rect 26466 26618 26702 26854
rect 26786 26618 27022 26854
rect 26466 8938 26702 9174
rect 26786 8938 27022 9174
rect 26466 8618 26702 8854
rect 26786 8618 27022 8854
rect 30186 462776 30422 463012
rect 30506 462776 30742 463012
rect 30186 462456 30422 462692
rect 30506 462456 30742 462692
rect 30186 444658 30422 444894
rect 30506 444658 30742 444894
rect 30186 444338 30422 444574
rect 30506 444338 30742 444574
rect 30186 426658 30422 426894
rect 30506 426658 30742 426894
rect 30186 426338 30422 426574
rect 30506 426338 30742 426574
rect 30186 408658 30422 408894
rect 30506 408658 30742 408894
rect 30186 408338 30422 408574
rect 30506 408338 30742 408574
rect 30186 390658 30422 390894
rect 30506 390658 30742 390894
rect 30186 390338 30422 390574
rect 30506 390338 30742 390574
rect 30186 372658 30422 372894
rect 30506 372658 30742 372894
rect 30186 372338 30422 372574
rect 30506 372338 30742 372574
rect 30186 354658 30422 354894
rect 30506 354658 30742 354894
rect 30186 354338 30422 354574
rect 30506 354338 30742 354574
rect 30186 336658 30422 336894
rect 30506 336658 30742 336894
rect 30186 336338 30422 336574
rect 30506 336338 30742 336574
rect 30186 318658 30422 318894
rect 30506 318658 30742 318894
rect 30186 318338 30422 318574
rect 30506 318338 30742 318574
rect 30186 300658 30422 300894
rect 30506 300658 30742 300894
rect 30186 300338 30422 300574
rect 30506 300338 30742 300574
rect 30186 282658 30422 282894
rect 30506 282658 30742 282894
rect 30186 282338 30422 282574
rect 30506 282338 30742 282574
rect 30186 264658 30422 264894
rect 30506 264658 30742 264894
rect 30186 264338 30422 264574
rect 30506 264338 30742 264574
rect 30186 246658 30422 246894
rect 30506 246658 30742 246894
rect 30186 246338 30422 246574
rect 30506 246338 30742 246574
rect 30186 228658 30422 228894
rect 30506 228658 30742 228894
rect 30186 228338 30422 228574
rect 30506 228338 30742 228574
rect 30186 210658 30422 210894
rect 30506 210658 30742 210894
rect 30186 210338 30422 210574
rect 30506 210338 30742 210574
rect 30186 192658 30422 192894
rect 30506 192658 30742 192894
rect 30186 192338 30422 192574
rect 30506 192338 30742 192574
rect 30186 174658 30422 174894
rect 30506 174658 30742 174894
rect 30186 174338 30422 174574
rect 30506 174338 30742 174574
rect 30186 156658 30422 156894
rect 30506 156658 30742 156894
rect 30186 156338 30422 156574
rect 30506 156338 30742 156574
rect 30186 138658 30422 138894
rect 30506 138658 30742 138894
rect 30186 138338 30422 138574
rect 30506 138338 30742 138574
rect 30186 120658 30422 120894
rect 30506 120658 30742 120894
rect 30186 120338 30422 120574
rect 30506 120338 30742 120574
rect 30186 102658 30422 102894
rect 30506 102658 30742 102894
rect 30186 102338 30422 102574
rect 30506 102338 30742 102574
rect 30186 84658 30422 84894
rect 30506 84658 30742 84894
rect 30186 84338 30422 84574
rect 30506 84338 30742 84574
rect 30186 66658 30422 66894
rect 30506 66658 30742 66894
rect 30186 66338 30422 66574
rect 30506 66338 30742 66574
rect 30186 48658 30422 48894
rect 30506 48658 30742 48894
rect 30186 48338 30422 48574
rect 30506 48338 30742 48574
rect 30186 30658 30422 30894
rect 30506 30658 30742 30894
rect 30186 30338 30422 30574
rect 30506 30338 30742 30574
rect 30186 12658 30422 12894
rect 30506 12658 30742 12894
rect 30186 12338 30422 12574
rect 30506 12338 30742 12574
rect 33906 463736 34142 463972
rect 34226 463736 34462 463972
rect 33906 463416 34142 463652
rect 34226 463416 34462 463652
rect 33906 448378 34142 448614
rect 34226 448378 34462 448614
rect 33906 448058 34142 448294
rect 34226 448058 34462 448294
rect 33906 430378 34142 430614
rect 34226 430378 34462 430614
rect 33906 430058 34142 430294
rect 34226 430058 34462 430294
rect 33906 412378 34142 412614
rect 34226 412378 34462 412614
rect 33906 412058 34142 412294
rect 34226 412058 34462 412294
rect 33906 394378 34142 394614
rect 34226 394378 34462 394614
rect 33906 394058 34142 394294
rect 34226 394058 34462 394294
rect 33906 376378 34142 376614
rect 34226 376378 34462 376614
rect 33906 376058 34142 376294
rect 34226 376058 34462 376294
rect 33906 358378 34142 358614
rect 34226 358378 34462 358614
rect 33906 358058 34142 358294
rect 34226 358058 34462 358294
rect 33906 340378 34142 340614
rect 34226 340378 34462 340614
rect 33906 340058 34142 340294
rect 34226 340058 34462 340294
rect 33906 322378 34142 322614
rect 34226 322378 34462 322614
rect 33906 322058 34142 322294
rect 34226 322058 34462 322294
rect 33906 304378 34142 304614
rect 34226 304378 34462 304614
rect 33906 304058 34142 304294
rect 34226 304058 34462 304294
rect 33906 286378 34142 286614
rect 34226 286378 34462 286614
rect 33906 286058 34142 286294
rect 34226 286058 34462 286294
rect 33906 268378 34142 268614
rect 34226 268378 34462 268614
rect 33906 268058 34142 268294
rect 34226 268058 34462 268294
rect 33906 250378 34142 250614
rect 34226 250378 34462 250614
rect 33906 250058 34142 250294
rect 34226 250058 34462 250294
rect 33906 232378 34142 232614
rect 34226 232378 34462 232614
rect 33906 232058 34142 232294
rect 34226 232058 34462 232294
rect 33906 214378 34142 214614
rect 34226 214378 34462 214614
rect 33906 214058 34142 214294
rect 34226 214058 34462 214294
rect 33906 196378 34142 196614
rect 34226 196378 34462 196614
rect 33906 196058 34142 196294
rect 34226 196058 34462 196294
rect 33906 178378 34142 178614
rect 34226 178378 34462 178614
rect 33906 178058 34142 178294
rect 34226 178058 34462 178294
rect 33906 160378 34142 160614
rect 34226 160378 34462 160614
rect 33906 160058 34142 160294
rect 34226 160058 34462 160294
rect 33906 142378 34142 142614
rect 34226 142378 34462 142614
rect 33906 142058 34142 142294
rect 34226 142058 34462 142294
rect 33906 124378 34142 124614
rect 34226 124378 34462 124614
rect 33906 124058 34142 124294
rect 34226 124058 34462 124294
rect 33906 106378 34142 106614
rect 34226 106378 34462 106614
rect 33906 106058 34142 106294
rect 34226 106058 34462 106294
rect 33906 88378 34142 88614
rect 34226 88378 34462 88614
rect 33906 88058 34142 88294
rect 34226 88058 34462 88294
rect 33906 70378 34142 70614
rect 34226 70378 34462 70614
rect 33906 70058 34142 70294
rect 34226 70058 34462 70294
rect 33906 52378 34142 52614
rect 34226 52378 34462 52614
rect 33906 52058 34142 52294
rect 34226 52058 34462 52294
rect 33906 34378 34142 34614
rect 34226 34378 34462 34614
rect 33906 34058 34142 34294
rect 34226 34058 34462 34294
rect 33906 16378 34142 16614
rect 34226 16378 34462 16614
rect 33906 16058 34142 16294
rect 34226 16058 34462 16294
rect 40746 460856 40982 461092
rect 41066 460856 41302 461092
rect 40746 460536 40982 460772
rect 41066 460536 41302 460772
rect 40746 455218 40982 455454
rect 41066 455218 41302 455454
rect 40746 454898 40982 455134
rect 41066 454898 41302 455134
rect 40746 437218 40982 437454
rect 41066 437218 41302 437454
rect 40746 436898 40982 437134
rect 41066 436898 41302 437134
rect 40746 419218 40982 419454
rect 41066 419218 41302 419454
rect 40746 418898 40982 419134
rect 41066 418898 41302 419134
rect 40746 401218 40982 401454
rect 41066 401218 41302 401454
rect 40746 400898 40982 401134
rect 41066 400898 41302 401134
rect 40746 383218 40982 383454
rect 41066 383218 41302 383454
rect 40746 382898 40982 383134
rect 41066 382898 41302 383134
rect 40746 365218 40982 365454
rect 41066 365218 41302 365454
rect 40746 364898 40982 365134
rect 41066 364898 41302 365134
rect 40746 347218 40982 347454
rect 41066 347218 41302 347454
rect 40746 346898 40982 347134
rect 41066 346898 41302 347134
rect 40746 329218 40982 329454
rect 41066 329218 41302 329454
rect 40746 328898 40982 329134
rect 41066 328898 41302 329134
rect 40746 311218 40982 311454
rect 41066 311218 41302 311454
rect 40746 310898 40982 311134
rect 41066 310898 41302 311134
rect 40746 293218 40982 293454
rect 41066 293218 41302 293454
rect 40746 292898 40982 293134
rect 41066 292898 41302 293134
rect 40746 275218 40982 275454
rect 41066 275218 41302 275454
rect 40746 274898 40982 275134
rect 41066 274898 41302 275134
rect 40746 257218 40982 257454
rect 41066 257218 41302 257454
rect 40746 256898 40982 257134
rect 41066 256898 41302 257134
rect 40746 239218 40982 239454
rect 41066 239218 41302 239454
rect 40746 238898 40982 239134
rect 41066 238898 41302 239134
rect 40746 221218 40982 221454
rect 41066 221218 41302 221454
rect 40746 220898 40982 221134
rect 41066 220898 41302 221134
rect 40746 203218 40982 203454
rect 41066 203218 41302 203454
rect 40746 202898 40982 203134
rect 41066 202898 41302 203134
rect 40746 185218 40982 185454
rect 41066 185218 41302 185454
rect 40746 184898 40982 185134
rect 41066 184898 41302 185134
rect 40746 167218 40982 167454
rect 41066 167218 41302 167454
rect 40746 166898 40982 167134
rect 41066 166898 41302 167134
rect 40746 149218 40982 149454
rect 41066 149218 41302 149454
rect 40746 148898 40982 149134
rect 41066 148898 41302 149134
rect 40746 131218 40982 131454
rect 41066 131218 41302 131454
rect 40746 130898 40982 131134
rect 41066 130898 41302 131134
rect 40746 113218 40982 113454
rect 41066 113218 41302 113454
rect 40746 112898 40982 113134
rect 41066 112898 41302 113134
rect 40746 95218 40982 95454
rect 41066 95218 41302 95454
rect 40746 94898 40982 95134
rect 41066 94898 41302 95134
rect 40746 77218 40982 77454
rect 41066 77218 41302 77454
rect 40746 76898 40982 77134
rect 41066 76898 41302 77134
rect 40746 59218 40982 59454
rect 41066 59218 41302 59454
rect 40746 58898 40982 59134
rect 41066 58898 41302 59134
rect 40746 41218 40982 41454
rect 41066 41218 41302 41454
rect 40746 40898 40982 41134
rect 41066 40898 41302 41134
rect 40746 23218 40982 23454
rect 41066 23218 41302 23454
rect 40746 22898 40982 23134
rect 41066 22898 41302 23134
rect 40746 5218 40982 5454
rect 41066 5218 41302 5454
rect 40746 4898 40982 5134
rect 41066 4898 41302 5134
rect 44466 461816 44702 462052
rect 44786 461816 45022 462052
rect 44466 461496 44702 461732
rect 44786 461496 45022 461732
rect 44466 440938 44702 441174
rect 44786 440938 45022 441174
rect 44466 440618 44702 440854
rect 44786 440618 45022 440854
rect 44466 422938 44702 423174
rect 44786 422938 45022 423174
rect 44466 422618 44702 422854
rect 44786 422618 45022 422854
rect 44466 404938 44702 405174
rect 44786 404938 45022 405174
rect 44466 404618 44702 404854
rect 44786 404618 45022 404854
rect 44466 386938 44702 387174
rect 44786 386938 45022 387174
rect 44466 386618 44702 386854
rect 44786 386618 45022 386854
rect 44466 368938 44702 369174
rect 44786 368938 45022 369174
rect 44466 368618 44702 368854
rect 44786 368618 45022 368854
rect 44466 350938 44702 351174
rect 44786 350938 45022 351174
rect 44466 350618 44702 350854
rect 44786 350618 45022 350854
rect 44466 332938 44702 333174
rect 44786 332938 45022 333174
rect 44466 332618 44702 332854
rect 44786 332618 45022 332854
rect 44466 314938 44702 315174
rect 44786 314938 45022 315174
rect 44466 314618 44702 314854
rect 44786 314618 45022 314854
rect 44466 296938 44702 297174
rect 44786 296938 45022 297174
rect 44466 296618 44702 296854
rect 44786 296618 45022 296854
rect 44466 278938 44702 279174
rect 44786 278938 45022 279174
rect 44466 278618 44702 278854
rect 44786 278618 45022 278854
rect 44466 260938 44702 261174
rect 44786 260938 45022 261174
rect 44466 260618 44702 260854
rect 44786 260618 45022 260854
rect 44466 242938 44702 243174
rect 44786 242938 45022 243174
rect 44466 242618 44702 242854
rect 44786 242618 45022 242854
rect 44466 224938 44702 225174
rect 44786 224938 45022 225174
rect 44466 224618 44702 224854
rect 44786 224618 45022 224854
rect 44466 206938 44702 207174
rect 44786 206938 45022 207174
rect 44466 206618 44702 206854
rect 44786 206618 45022 206854
rect 44466 188938 44702 189174
rect 44786 188938 45022 189174
rect 44466 188618 44702 188854
rect 44786 188618 45022 188854
rect 44466 170938 44702 171174
rect 44786 170938 45022 171174
rect 44466 170618 44702 170854
rect 44786 170618 45022 170854
rect 44466 152938 44702 153174
rect 44786 152938 45022 153174
rect 44466 152618 44702 152854
rect 44786 152618 45022 152854
rect 44466 134938 44702 135174
rect 44786 134938 45022 135174
rect 44466 134618 44702 134854
rect 44786 134618 45022 134854
rect 44466 116938 44702 117174
rect 44786 116938 45022 117174
rect 44466 116618 44702 116854
rect 44786 116618 45022 116854
rect 44466 98938 44702 99174
rect 44786 98938 45022 99174
rect 44466 98618 44702 98854
rect 44786 98618 45022 98854
rect 44466 80938 44702 81174
rect 44786 80938 45022 81174
rect 44466 80618 44702 80854
rect 44786 80618 45022 80854
rect 44466 62938 44702 63174
rect 44786 62938 45022 63174
rect 44466 62618 44702 62854
rect 44786 62618 45022 62854
rect 44466 44938 44702 45174
rect 44786 44938 45022 45174
rect 44466 44618 44702 44854
rect 44786 44618 45022 44854
rect 44466 26938 44702 27174
rect 44786 26938 45022 27174
rect 44466 26618 44702 26854
rect 44786 26618 45022 26854
rect 44466 8938 44702 9174
rect 44786 8938 45022 9174
rect 44466 8618 44702 8854
rect 44786 8618 45022 8854
rect 48186 462776 48422 463012
rect 48506 462776 48742 463012
rect 48186 462456 48422 462692
rect 48506 462456 48742 462692
rect 48186 444658 48422 444894
rect 48506 444658 48742 444894
rect 48186 444338 48422 444574
rect 48506 444338 48742 444574
rect 48186 426658 48422 426894
rect 48506 426658 48742 426894
rect 48186 426338 48422 426574
rect 48506 426338 48742 426574
rect 48186 408658 48422 408894
rect 48506 408658 48742 408894
rect 48186 408338 48422 408574
rect 48506 408338 48742 408574
rect 48186 390658 48422 390894
rect 48506 390658 48742 390894
rect 48186 390338 48422 390574
rect 48506 390338 48742 390574
rect 48186 372658 48422 372894
rect 48506 372658 48742 372894
rect 48186 372338 48422 372574
rect 48506 372338 48742 372574
rect 48186 354658 48422 354894
rect 48506 354658 48742 354894
rect 48186 354338 48422 354574
rect 48506 354338 48742 354574
rect 48186 336658 48422 336894
rect 48506 336658 48742 336894
rect 48186 336338 48422 336574
rect 48506 336338 48742 336574
rect 48186 318658 48422 318894
rect 48506 318658 48742 318894
rect 48186 318338 48422 318574
rect 48506 318338 48742 318574
rect 48186 300658 48422 300894
rect 48506 300658 48742 300894
rect 48186 300338 48422 300574
rect 48506 300338 48742 300574
rect 48186 282658 48422 282894
rect 48506 282658 48742 282894
rect 48186 282338 48422 282574
rect 48506 282338 48742 282574
rect 48186 264658 48422 264894
rect 48506 264658 48742 264894
rect 48186 264338 48422 264574
rect 48506 264338 48742 264574
rect 48186 246658 48422 246894
rect 48506 246658 48742 246894
rect 48186 246338 48422 246574
rect 48506 246338 48742 246574
rect 48186 228658 48422 228894
rect 48506 228658 48742 228894
rect 48186 228338 48422 228574
rect 48506 228338 48742 228574
rect 48186 210658 48422 210894
rect 48506 210658 48742 210894
rect 48186 210338 48422 210574
rect 48506 210338 48742 210574
rect 48186 192658 48422 192894
rect 48506 192658 48742 192894
rect 48186 192338 48422 192574
rect 48506 192338 48742 192574
rect 48186 174658 48422 174894
rect 48506 174658 48742 174894
rect 48186 174338 48422 174574
rect 48506 174338 48742 174574
rect 48186 156658 48422 156894
rect 48506 156658 48742 156894
rect 48186 156338 48422 156574
rect 48506 156338 48742 156574
rect 48186 138658 48422 138894
rect 48506 138658 48742 138894
rect 48186 138338 48422 138574
rect 48506 138338 48742 138574
rect 48186 120658 48422 120894
rect 48506 120658 48742 120894
rect 48186 120338 48422 120574
rect 48506 120338 48742 120574
rect 48186 102658 48422 102894
rect 48506 102658 48742 102894
rect 48186 102338 48422 102574
rect 48506 102338 48742 102574
rect 48186 84658 48422 84894
rect 48506 84658 48742 84894
rect 48186 84338 48422 84574
rect 48506 84338 48742 84574
rect 48186 66658 48422 66894
rect 48506 66658 48742 66894
rect 48186 66338 48422 66574
rect 48506 66338 48742 66574
rect 48186 48658 48422 48894
rect 48506 48658 48742 48894
rect 48186 48338 48422 48574
rect 48506 48338 48742 48574
rect 48186 30658 48422 30894
rect 48506 30658 48742 30894
rect 48186 30338 48422 30574
rect 48506 30338 48742 30574
rect 48186 12658 48422 12894
rect 48506 12658 48742 12894
rect 48186 12338 48422 12574
rect 48506 12338 48742 12574
rect -1564 -1092 -1328 -856
rect -1244 -1092 -1008 -856
rect -1564 -1412 -1328 -1176
rect -1244 -1412 -1008 -1176
rect -2524 -2052 -2288 -1816
rect -2204 -2052 -1968 -1816
rect -2524 -2372 -2288 -2136
rect -2204 -2372 -1968 -2136
rect -3484 -3012 -3248 -2776
rect -3164 -3012 -2928 -2776
rect -3484 -3332 -3248 -3096
rect -3164 -3332 -2928 -3096
rect 48186 -3012 48422 -2776
rect 48506 -3012 48742 -2776
rect 48186 -3332 48422 -3096
rect 48506 -3332 48742 -3096
rect -4444 -3972 -4208 -3736
rect -4124 -3972 -3888 -3736
rect -4444 -4292 -4208 -4056
rect -4124 -4292 -3888 -4056
rect 51906 463736 52142 463972
rect 52226 463736 52462 463972
rect 51906 463416 52142 463652
rect 52226 463416 52462 463652
rect 51906 448378 52142 448614
rect 52226 448378 52462 448614
rect 51906 448058 52142 448294
rect 52226 448058 52462 448294
rect 51906 430378 52142 430614
rect 52226 430378 52462 430614
rect 51906 430058 52142 430294
rect 52226 430058 52462 430294
rect 51906 412378 52142 412614
rect 52226 412378 52462 412614
rect 51906 412058 52142 412294
rect 52226 412058 52462 412294
rect 51906 394378 52142 394614
rect 52226 394378 52462 394614
rect 51906 394058 52142 394294
rect 52226 394058 52462 394294
rect 51906 376378 52142 376614
rect 52226 376378 52462 376614
rect 51906 376058 52142 376294
rect 52226 376058 52462 376294
rect 51906 358378 52142 358614
rect 52226 358378 52462 358614
rect 51906 358058 52142 358294
rect 52226 358058 52462 358294
rect 51906 340378 52142 340614
rect 52226 340378 52462 340614
rect 51906 340058 52142 340294
rect 52226 340058 52462 340294
rect 51906 322378 52142 322614
rect 52226 322378 52462 322614
rect 51906 322058 52142 322294
rect 52226 322058 52462 322294
rect 51906 304378 52142 304614
rect 52226 304378 52462 304614
rect 51906 304058 52142 304294
rect 52226 304058 52462 304294
rect 51906 286378 52142 286614
rect 52226 286378 52462 286614
rect 51906 286058 52142 286294
rect 52226 286058 52462 286294
rect 51906 268378 52142 268614
rect 52226 268378 52462 268614
rect 51906 268058 52142 268294
rect 52226 268058 52462 268294
rect 51906 250378 52142 250614
rect 52226 250378 52462 250614
rect 51906 250058 52142 250294
rect 52226 250058 52462 250294
rect 51906 232378 52142 232614
rect 52226 232378 52462 232614
rect 51906 232058 52142 232294
rect 52226 232058 52462 232294
rect 51906 214378 52142 214614
rect 52226 214378 52462 214614
rect 51906 214058 52142 214294
rect 52226 214058 52462 214294
rect 51906 196378 52142 196614
rect 52226 196378 52462 196614
rect 51906 196058 52142 196294
rect 52226 196058 52462 196294
rect 51906 178378 52142 178614
rect 52226 178378 52462 178614
rect 51906 178058 52142 178294
rect 52226 178058 52462 178294
rect 51906 160378 52142 160614
rect 52226 160378 52462 160614
rect 51906 160058 52142 160294
rect 52226 160058 52462 160294
rect 51906 142378 52142 142614
rect 52226 142378 52462 142614
rect 51906 142058 52142 142294
rect 52226 142058 52462 142294
rect 51906 124378 52142 124614
rect 52226 124378 52462 124614
rect 51906 124058 52142 124294
rect 52226 124058 52462 124294
rect 51906 106378 52142 106614
rect 52226 106378 52462 106614
rect 51906 106058 52142 106294
rect 52226 106058 52462 106294
rect 51906 88378 52142 88614
rect 52226 88378 52462 88614
rect 51906 88058 52142 88294
rect 52226 88058 52462 88294
rect 51906 70378 52142 70614
rect 52226 70378 52462 70614
rect 51906 70058 52142 70294
rect 52226 70058 52462 70294
rect 51906 52378 52142 52614
rect 52226 52378 52462 52614
rect 51906 52058 52142 52294
rect 52226 52058 52462 52294
rect 51906 34378 52142 34614
rect 52226 34378 52462 34614
rect 51906 34058 52142 34294
rect 52226 34058 52462 34294
rect 51906 16378 52142 16614
rect 52226 16378 52462 16614
rect 51906 16058 52142 16294
rect 52226 16058 52462 16294
rect 51906 -3972 52142 -3736
rect 52226 -3972 52462 -3736
rect 51906 -4292 52142 -4056
rect 52226 -4292 52462 -4056
rect 58746 460856 58982 461092
rect 59066 460856 59302 461092
rect 58746 460536 58982 460772
rect 59066 460536 59302 460772
rect 58746 455218 58982 455454
rect 59066 455218 59302 455454
rect 58746 454898 58982 455134
rect 59066 454898 59302 455134
rect 58746 437218 58982 437454
rect 59066 437218 59302 437454
rect 58746 436898 58982 437134
rect 59066 436898 59302 437134
rect 58746 419218 58982 419454
rect 59066 419218 59302 419454
rect 58746 418898 58982 419134
rect 59066 418898 59302 419134
rect 58746 401218 58982 401454
rect 59066 401218 59302 401454
rect 58746 400898 58982 401134
rect 59066 400898 59302 401134
rect 58746 383218 58982 383454
rect 59066 383218 59302 383454
rect 58746 382898 58982 383134
rect 59066 382898 59302 383134
rect 58746 365218 58982 365454
rect 59066 365218 59302 365454
rect 58746 364898 58982 365134
rect 59066 364898 59302 365134
rect 58746 347218 58982 347454
rect 59066 347218 59302 347454
rect 58746 346898 58982 347134
rect 59066 346898 59302 347134
rect 58746 329218 58982 329454
rect 59066 329218 59302 329454
rect 58746 328898 58982 329134
rect 59066 328898 59302 329134
rect 58746 311218 58982 311454
rect 59066 311218 59302 311454
rect 58746 310898 58982 311134
rect 59066 310898 59302 311134
rect 58746 293218 58982 293454
rect 59066 293218 59302 293454
rect 58746 292898 58982 293134
rect 59066 292898 59302 293134
rect 58746 275218 58982 275454
rect 59066 275218 59302 275454
rect 58746 274898 58982 275134
rect 59066 274898 59302 275134
rect 58746 257218 58982 257454
rect 59066 257218 59302 257454
rect 58746 256898 58982 257134
rect 59066 256898 59302 257134
rect 58746 239218 58982 239454
rect 59066 239218 59302 239454
rect 58746 238898 58982 239134
rect 59066 238898 59302 239134
rect 58746 221218 58982 221454
rect 59066 221218 59302 221454
rect 58746 220898 58982 221134
rect 59066 220898 59302 221134
rect 58746 203218 58982 203454
rect 59066 203218 59302 203454
rect 58746 202898 58982 203134
rect 59066 202898 59302 203134
rect 58746 185218 58982 185454
rect 59066 185218 59302 185454
rect 58746 184898 58982 185134
rect 59066 184898 59302 185134
rect 58746 167218 58982 167454
rect 59066 167218 59302 167454
rect 58746 166898 58982 167134
rect 59066 166898 59302 167134
rect 58746 149218 58982 149454
rect 59066 149218 59302 149454
rect 58746 148898 58982 149134
rect 59066 148898 59302 149134
rect 58746 131218 58982 131454
rect 59066 131218 59302 131454
rect 58746 130898 58982 131134
rect 59066 130898 59302 131134
rect 58746 113218 58982 113454
rect 59066 113218 59302 113454
rect 58746 112898 58982 113134
rect 59066 112898 59302 113134
rect 58746 95218 58982 95454
rect 59066 95218 59302 95454
rect 58746 94898 58982 95134
rect 59066 94898 59302 95134
rect 58746 77218 58982 77454
rect 59066 77218 59302 77454
rect 58746 76898 58982 77134
rect 59066 76898 59302 77134
rect 58746 59218 58982 59454
rect 59066 59218 59302 59454
rect 58746 58898 58982 59134
rect 59066 58898 59302 59134
rect 58746 41218 58982 41454
rect 59066 41218 59302 41454
rect 58746 40898 58982 41134
rect 59066 40898 59302 41134
rect 58746 23218 58982 23454
rect 59066 23218 59302 23454
rect 58746 22898 58982 23134
rect 59066 22898 59302 23134
rect 58746 5218 58982 5454
rect 59066 5218 59302 5454
rect 58746 4898 58982 5134
rect 59066 4898 59302 5134
rect 58746 -1092 58982 -856
rect 59066 -1092 59302 -856
rect 58746 -1412 58982 -1176
rect 59066 -1412 59302 -1176
rect 62466 461816 62702 462052
rect 62786 461816 63022 462052
rect 62466 461496 62702 461732
rect 62786 461496 63022 461732
rect 62466 440938 62702 441174
rect 62786 440938 63022 441174
rect 62466 440618 62702 440854
rect 62786 440618 63022 440854
rect 62466 422938 62702 423174
rect 62786 422938 63022 423174
rect 62466 422618 62702 422854
rect 62786 422618 63022 422854
rect 62466 404938 62702 405174
rect 62786 404938 63022 405174
rect 62466 404618 62702 404854
rect 62786 404618 63022 404854
rect 62466 386938 62702 387174
rect 62786 386938 63022 387174
rect 62466 386618 62702 386854
rect 62786 386618 63022 386854
rect 62466 368938 62702 369174
rect 62786 368938 63022 369174
rect 62466 368618 62702 368854
rect 62786 368618 63022 368854
rect 62466 350938 62702 351174
rect 62786 350938 63022 351174
rect 62466 350618 62702 350854
rect 62786 350618 63022 350854
rect 62466 332938 62702 333174
rect 62786 332938 63022 333174
rect 62466 332618 62702 332854
rect 62786 332618 63022 332854
rect 62466 314938 62702 315174
rect 62786 314938 63022 315174
rect 62466 314618 62702 314854
rect 62786 314618 63022 314854
rect 62466 296938 62702 297174
rect 62786 296938 63022 297174
rect 62466 296618 62702 296854
rect 62786 296618 63022 296854
rect 62466 278938 62702 279174
rect 62786 278938 63022 279174
rect 62466 278618 62702 278854
rect 62786 278618 63022 278854
rect 62466 260938 62702 261174
rect 62786 260938 63022 261174
rect 62466 260618 62702 260854
rect 62786 260618 63022 260854
rect 62466 242938 62702 243174
rect 62786 242938 63022 243174
rect 62466 242618 62702 242854
rect 62786 242618 63022 242854
rect 62466 224938 62702 225174
rect 62786 224938 63022 225174
rect 62466 224618 62702 224854
rect 62786 224618 63022 224854
rect 62466 206938 62702 207174
rect 62786 206938 63022 207174
rect 62466 206618 62702 206854
rect 62786 206618 63022 206854
rect 62466 188938 62702 189174
rect 62786 188938 63022 189174
rect 62466 188618 62702 188854
rect 62786 188618 63022 188854
rect 62466 170938 62702 171174
rect 62786 170938 63022 171174
rect 62466 170618 62702 170854
rect 62786 170618 63022 170854
rect 62466 152938 62702 153174
rect 62786 152938 63022 153174
rect 62466 152618 62702 152854
rect 62786 152618 63022 152854
rect 62466 134938 62702 135174
rect 62786 134938 63022 135174
rect 62466 134618 62702 134854
rect 62786 134618 63022 134854
rect 62466 116938 62702 117174
rect 62786 116938 63022 117174
rect 62466 116618 62702 116854
rect 62786 116618 63022 116854
rect 62466 98938 62702 99174
rect 62786 98938 63022 99174
rect 62466 98618 62702 98854
rect 62786 98618 63022 98854
rect 62466 80938 62702 81174
rect 62786 80938 63022 81174
rect 62466 80618 62702 80854
rect 62786 80618 63022 80854
rect 62466 62938 62702 63174
rect 62786 62938 63022 63174
rect 62466 62618 62702 62854
rect 62786 62618 63022 62854
rect 62466 44938 62702 45174
rect 62786 44938 63022 45174
rect 62466 44618 62702 44854
rect 62786 44618 63022 44854
rect 62466 26938 62702 27174
rect 62786 26938 63022 27174
rect 62466 26618 62702 26854
rect 62786 26618 63022 26854
rect 62466 8938 62702 9174
rect 62786 8938 63022 9174
rect 62466 8618 62702 8854
rect 62786 8618 63022 8854
rect 62466 -2052 62702 -1816
rect 62786 -2052 63022 -1816
rect 62466 -2372 62702 -2136
rect 62786 -2372 63022 -2136
rect 66186 462776 66422 463012
rect 66506 462776 66742 463012
rect 66186 462456 66422 462692
rect 66506 462456 66742 462692
rect 66186 444658 66422 444894
rect 66506 444658 66742 444894
rect 66186 444338 66422 444574
rect 66506 444338 66742 444574
rect 66186 426658 66422 426894
rect 66506 426658 66742 426894
rect 66186 426338 66422 426574
rect 66506 426338 66742 426574
rect 66186 408658 66422 408894
rect 66506 408658 66742 408894
rect 66186 408338 66422 408574
rect 66506 408338 66742 408574
rect 66186 390658 66422 390894
rect 66506 390658 66742 390894
rect 66186 390338 66422 390574
rect 66506 390338 66742 390574
rect 66186 372658 66422 372894
rect 66506 372658 66742 372894
rect 66186 372338 66422 372574
rect 66506 372338 66742 372574
rect 66186 354658 66422 354894
rect 66506 354658 66742 354894
rect 66186 354338 66422 354574
rect 66506 354338 66742 354574
rect 66186 336658 66422 336894
rect 66506 336658 66742 336894
rect 66186 336338 66422 336574
rect 66506 336338 66742 336574
rect 66186 318658 66422 318894
rect 66506 318658 66742 318894
rect 66186 318338 66422 318574
rect 66506 318338 66742 318574
rect 66186 300658 66422 300894
rect 66506 300658 66742 300894
rect 66186 300338 66422 300574
rect 66506 300338 66742 300574
rect 66186 282658 66422 282894
rect 66506 282658 66742 282894
rect 66186 282338 66422 282574
rect 66506 282338 66742 282574
rect 66186 264658 66422 264894
rect 66506 264658 66742 264894
rect 66186 264338 66422 264574
rect 66506 264338 66742 264574
rect 66186 246658 66422 246894
rect 66506 246658 66742 246894
rect 66186 246338 66422 246574
rect 66506 246338 66742 246574
rect 66186 228658 66422 228894
rect 66506 228658 66742 228894
rect 66186 228338 66422 228574
rect 66506 228338 66742 228574
rect 66186 210658 66422 210894
rect 66506 210658 66742 210894
rect 66186 210338 66422 210574
rect 66506 210338 66742 210574
rect 66186 192658 66422 192894
rect 66506 192658 66742 192894
rect 66186 192338 66422 192574
rect 66506 192338 66742 192574
rect 66186 174658 66422 174894
rect 66506 174658 66742 174894
rect 66186 174338 66422 174574
rect 66506 174338 66742 174574
rect 66186 156658 66422 156894
rect 66506 156658 66742 156894
rect 66186 156338 66422 156574
rect 66506 156338 66742 156574
rect 66186 138658 66422 138894
rect 66506 138658 66742 138894
rect 66186 138338 66422 138574
rect 66506 138338 66742 138574
rect 66186 120658 66422 120894
rect 66506 120658 66742 120894
rect 66186 120338 66422 120574
rect 66506 120338 66742 120574
rect 66186 102658 66422 102894
rect 66506 102658 66742 102894
rect 66186 102338 66422 102574
rect 66506 102338 66742 102574
rect 66186 84658 66422 84894
rect 66506 84658 66742 84894
rect 66186 84338 66422 84574
rect 66506 84338 66742 84574
rect 66186 66658 66422 66894
rect 66506 66658 66742 66894
rect 66186 66338 66422 66574
rect 66506 66338 66742 66574
rect 66186 48658 66422 48894
rect 66506 48658 66742 48894
rect 66186 48338 66422 48574
rect 66506 48338 66742 48574
rect 66186 30658 66422 30894
rect 66506 30658 66742 30894
rect 66186 30338 66422 30574
rect 66506 30338 66742 30574
rect 66186 12658 66422 12894
rect 66506 12658 66742 12894
rect 66186 12338 66422 12574
rect 66506 12338 66742 12574
rect 66186 -3012 66422 -2776
rect 66506 -3012 66742 -2776
rect 66186 -3332 66422 -3096
rect 66506 -3332 66742 -3096
rect 69906 463736 70142 463972
rect 70226 463736 70462 463972
rect 69906 463416 70142 463652
rect 70226 463416 70462 463652
rect 69906 448378 70142 448614
rect 70226 448378 70462 448614
rect 69906 448058 70142 448294
rect 70226 448058 70462 448294
rect 69906 430378 70142 430614
rect 70226 430378 70462 430614
rect 69906 430058 70142 430294
rect 70226 430058 70462 430294
rect 69906 412378 70142 412614
rect 70226 412378 70462 412614
rect 69906 412058 70142 412294
rect 70226 412058 70462 412294
rect 69906 394378 70142 394614
rect 70226 394378 70462 394614
rect 69906 394058 70142 394294
rect 70226 394058 70462 394294
rect 69906 376378 70142 376614
rect 70226 376378 70462 376614
rect 69906 376058 70142 376294
rect 70226 376058 70462 376294
rect 69906 358378 70142 358614
rect 70226 358378 70462 358614
rect 69906 358058 70142 358294
rect 70226 358058 70462 358294
rect 69906 340378 70142 340614
rect 70226 340378 70462 340614
rect 69906 340058 70142 340294
rect 70226 340058 70462 340294
rect 69906 322378 70142 322614
rect 70226 322378 70462 322614
rect 69906 322058 70142 322294
rect 70226 322058 70462 322294
rect 69906 304378 70142 304614
rect 70226 304378 70462 304614
rect 69906 304058 70142 304294
rect 70226 304058 70462 304294
rect 69906 286378 70142 286614
rect 70226 286378 70462 286614
rect 69906 286058 70142 286294
rect 70226 286058 70462 286294
rect 69906 268378 70142 268614
rect 70226 268378 70462 268614
rect 69906 268058 70142 268294
rect 70226 268058 70462 268294
rect 69906 250378 70142 250614
rect 70226 250378 70462 250614
rect 69906 250058 70142 250294
rect 70226 250058 70462 250294
rect 69906 232378 70142 232614
rect 70226 232378 70462 232614
rect 69906 232058 70142 232294
rect 70226 232058 70462 232294
rect 69906 214378 70142 214614
rect 70226 214378 70462 214614
rect 69906 214058 70142 214294
rect 70226 214058 70462 214294
rect 69906 196378 70142 196614
rect 70226 196378 70462 196614
rect 69906 196058 70142 196294
rect 70226 196058 70462 196294
rect 69906 178378 70142 178614
rect 70226 178378 70462 178614
rect 69906 178058 70142 178294
rect 70226 178058 70462 178294
rect 69906 160378 70142 160614
rect 70226 160378 70462 160614
rect 69906 160058 70142 160294
rect 70226 160058 70462 160294
rect 69906 142378 70142 142614
rect 70226 142378 70462 142614
rect 69906 142058 70142 142294
rect 70226 142058 70462 142294
rect 69906 124378 70142 124614
rect 70226 124378 70462 124614
rect 69906 124058 70142 124294
rect 70226 124058 70462 124294
rect 69906 106378 70142 106614
rect 70226 106378 70462 106614
rect 69906 106058 70142 106294
rect 70226 106058 70462 106294
rect 69906 88378 70142 88614
rect 70226 88378 70462 88614
rect 69906 88058 70142 88294
rect 70226 88058 70462 88294
rect 69906 70378 70142 70614
rect 70226 70378 70462 70614
rect 69906 70058 70142 70294
rect 70226 70058 70462 70294
rect 69906 52378 70142 52614
rect 70226 52378 70462 52614
rect 69906 52058 70142 52294
rect 70226 52058 70462 52294
rect 69906 34378 70142 34614
rect 70226 34378 70462 34614
rect 69906 34058 70142 34294
rect 70226 34058 70462 34294
rect 69906 16378 70142 16614
rect 70226 16378 70462 16614
rect 69906 16058 70142 16294
rect 70226 16058 70462 16294
rect 69906 -3972 70142 -3736
rect 70226 -3972 70462 -3736
rect 69906 -4292 70142 -4056
rect 70226 -4292 70462 -4056
rect 76746 460856 76982 461092
rect 77066 460856 77302 461092
rect 76746 460536 76982 460772
rect 77066 460536 77302 460772
rect 76746 455218 76982 455454
rect 77066 455218 77302 455454
rect 76746 454898 76982 455134
rect 77066 454898 77302 455134
rect 76746 437218 76982 437454
rect 77066 437218 77302 437454
rect 76746 436898 76982 437134
rect 77066 436898 77302 437134
rect 76746 419218 76982 419454
rect 77066 419218 77302 419454
rect 76746 418898 76982 419134
rect 77066 418898 77302 419134
rect 76746 401218 76982 401454
rect 77066 401218 77302 401454
rect 76746 400898 76982 401134
rect 77066 400898 77302 401134
rect 76746 383218 76982 383454
rect 77066 383218 77302 383454
rect 76746 382898 76982 383134
rect 77066 382898 77302 383134
rect 76746 365218 76982 365454
rect 77066 365218 77302 365454
rect 76746 364898 76982 365134
rect 77066 364898 77302 365134
rect 76746 347218 76982 347454
rect 77066 347218 77302 347454
rect 76746 346898 76982 347134
rect 77066 346898 77302 347134
rect 76746 329218 76982 329454
rect 77066 329218 77302 329454
rect 76746 328898 76982 329134
rect 77066 328898 77302 329134
rect 76746 311218 76982 311454
rect 77066 311218 77302 311454
rect 76746 310898 76982 311134
rect 77066 310898 77302 311134
rect 76746 293218 76982 293454
rect 77066 293218 77302 293454
rect 76746 292898 76982 293134
rect 77066 292898 77302 293134
rect 76746 275218 76982 275454
rect 77066 275218 77302 275454
rect 76746 274898 76982 275134
rect 77066 274898 77302 275134
rect 76746 257218 76982 257454
rect 77066 257218 77302 257454
rect 76746 256898 76982 257134
rect 77066 256898 77302 257134
rect 76746 239218 76982 239454
rect 77066 239218 77302 239454
rect 76746 238898 76982 239134
rect 77066 238898 77302 239134
rect 76746 221218 76982 221454
rect 77066 221218 77302 221454
rect 76746 220898 76982 221134
rect 77066 220898 77302 221134
rect 76746 203218 76982 203454
rect 77066 203218 77302 203454
rect 76746 202898 76982 203134
rect 77066 202898 77302 203134
rect 76746 185218 76982 185454
rect 77066 185218 77302 185454
rect 76746 184898 76982 185134
rect 77066 184898 77302 185134
rect 76746 167218 76982 167454
rect 77066 167218 77302 167454
rect 76746 166898 76982 167134
rect 77066 166898 77302 167134
rect 76746 149218 76982 149454
rect 77066 149218 77302 149454
rect 76746 148898 76982 149134
rect 77066 148898 77302 149134
rect 76746 131218 76982 131454
rect 77066 131218 77302 131454
rect 76746 130898 76982 131134
rect 77066 130898 77302 131134
rect 76746 113218 76982 113454
rect 77066 113218 77302 113454
rect 76746 112898 76982 113134
rect 77066 112898 77302 113134
rect 76746 95218 76982 95454
rect 77066 95218 77302 95454
rect 76746 94898 76982 95134
rect 77066 94898 77302 95134
rect 76746 77218 76982 77454
rect 77066 77218 77302 77454
rect 76746 76898 76982 77134
rect 77066 76898 77302 77134
rect 76746 59218 76982 59454
rect 77066 59218 77302 59454
rect 76746 58898 76982 59134
rect 77066 58898 77302 59134
rect 76746 41218 76982 41454
rect 77066 41218 77302 41454
rect 76746 40898 76982 41134
rect 77066 40898 77302 41134
rect 76746 23218 76982 23454
rect 77066 23218 77302 23454
rect 76746 22898 76982 23134
rect 77066 22898 77302 23134
rect 76746 5218 76982 5454
rect 77066 5218 77302 5454
rect 76746 4898 76982 5134
rect 77066 4898 77302 5134
rect 76746 -1092 76982 -856
rect 77066 -1092 77302 -856
rect 76746 -1412 76982 -1176
rect 77066 -1412 77302 -1176
rect 80466 461816 80702 462052
rect 80786 461816 81022 462052
rect 80466 461496 80702 461732
rect 80786 461496 81022 461732
rect 80466 440938 80702 441174
rect 80786 440938 81022 441174
rect 80466 440618 80702 440854
rect 80786 440618 81022 440854
rect 80466 422938 80702 423174
rect 80786 422938 81022 423174
rect 80466 422618 80702 422854
rect 80786 422618 81022 422854
rect 80466 404938 80702 405174
rect 80786 404938 81022 405174
rect 80466 404618 80702 404854
rect 80786 404618 81022 404854
rect 80466 386938 80702 387174
rect 80786 386938 81022 387174
rect 80466 386618 80702 386854
rect 80786 386618 81022 386854
rect 80466 368938 80702 369174
rect 80786 368938 81022 369174
rect 80466 368618 80702 368854
rect 80786 368618 81022 368854
rect 80466 350938 80702 351174
rect 80786 350938 81022 351174
rect 80466 350618 80702 350854
rect 80786 350618 81022 350854
rect 80466 332938 80702 333174
rect 80786 332938 81022 333174
rect 80466 332618 80702 332854
rect 80786 332618 81022 332854
rect 80466 314938 80702 315174
rect 80786 314938 81022 315174
rect 80466 314618 80702 314854
rect 80786 314618 81022 314854
rect 80466 296938 80702 297174
rect 80786 296938 81022 297174
rect 80466 296618 80702 296854
rect 80786 296618 81022 296854
rect 80466 278938 80702 279174
rect 80786 278938 81022 279174
rect 80466 278618 80702 278854
rect 80786 278618 81022 278854
rect 80466 260938 80702 261174
rect 80786 260938 81022 261174
rect 80466 260618 80702 260854
rect 80786 260618 81022 260854
rect 80466 242938 80702 243174
rect 80786 242938 81022 243174
rect 80466 242618 80702 242854
rect 80786 242618 81022 242854
rect 80466 224938 80702 225174
rect 80786 224938 81022 225174
rect 80466 224618 80702 224854
rect 80786 224618 81022 224854
rect 80466 206938 80702 207174
rect 80786 206938 81022 207174
rect 80466 206618 80702 206854
rect 80786 206618 81022 206854
rect 80466 188938 80702 189174
rect 80786 188938 81022 189174
rect 80466 188618 80702 188854
rect 80786 188618 81022 188854
rect 80466 170938 80702 171174
rect 80786 170938 81022 171174
rect 80466 170618 80702 170854
rect 80786 170618 81022 170854
rect 80466 152938 80702 153174
rect 80786 152938 81022 153174
rect 80466 152618 80702 152854
rect 80786 152618 81022 152854
rect 80466 134938 80702 135174
rect 80786 134938 81022 135174
rect 80466 134618 80702 134854
rect 80786 134618 81022 134854
rect 80466 116938 80702 117174
rect 80786 116938 81022 117174
rect 80466 116618 80702 116854
rect 80786 116618 81022 116854
rect 80466 98938 80702 99174
rect 80786 98938 81022 99174
rect 80466 98618 80702 98854
rect 80786 98618 81022 98854
rect 80466 80938 80702 81174
rect 80786 80938 81022 81174
rect 80466 80618 80702 80854
rect 80786 80618 81022 80854
rect 80466 62938 80702 63174
rect 80786 62938 81022 63174
rect 80466 62618 80702 62854
rect 80786 62618 81022 62854
rect 80466 44938 80702 45174
rect 80786 44938 81022 45174
rect 80466 44618 80702 44854
rect 80786 44618 81022 44854
rect 80466 26938 80702 27174
rect 80786 26938 81022 27174
rect 80466 26618 80702 26854
rect 80786 26618 81022 26854
rect 80466 8938 80702 9174
rect 80786 8938 81022 9174
rect 80466 8618 80702 8854
rect 80786 8618 81022 8854
rect 80466 -2052 80702 -1816
rect 80786 -2052 81022 -1816
rect 80466 -2372 80702 -2136
rect 80786 -2372 81022 -2136
rect 84186 462776 84422 463012
rect 84506 462776 84742 463012
rect 84186 462456 84422 462692
rect 84506 462456 84742 462692
rect 84186 444658 84422 444894
rect 84506 444658 84742 444894
rect 84186 444338 84422 444574
rect 84506 444338 84742 444574
rect 84186 426658 84422 426894
rect 84506 426658 84742 426894
rect 84186 426338 84422 426574
rect 84506 426338 84742 426574
rect 84186 408658 84422 408894
rect 84506 408658 84742 408894
rect 84186 408338 84422 408574
rect 84506 408338 84742 408574
rect 84186 390658 84422 390894
rect 84506 390658 84742 390894
rect 84186 390338 84422 390574
rect 84506 390338 84742 390574
rect 84186 372658 84422 372894
rect 84506 372658 84742 372894
rect 84186 372338 84422 372574
rect 84506 372338 84742 372574
rect 84186 354658 84422 354894
rect 84506 354658 84742 354894
rect 84186 354338 84422 354574
rect 84506 354338 84742 354574
rect 84186 336658 84422 336894
rect 84506 336658 84742 336894
rect 84186 336338 84422 336574
rect 84506 336338 84742 336574
rect 84186 318658 84422 318894
rect 84506 318658 84742 318894
rect 84186 318338 84422 318574
rect 84506 318338 84742 318574
rect 84186 300658 84422 300894
rect 84506 300658 84742 300894
rect 84186 300338 84422 300574
rect 84506 300338 84742 300574
rect 84186 282658 84422 282894
rect 84506 282658 84742 282894
rect 84186 282338 84422 282574
rect 84506 282338 84742 282574
rect 84186 264658 84422 264894
rect 84506 264658 84742 264894
rect 84186 264338 84422 264574
rect 84506 264338 84742 264574
rect 84186 246658 84422 246894
rect 84506 246658 84742 246894
rect 84186 246338 84422 246574
rect 84506 246338 84742 246574
rect 84186 228658 84422 228894
rect 84506 228658 84742 228894
rect 84186 228338 84422 228574
rect 84506 228338 84742 228574
rect 84186 210658 84422 210894
rect 84506 210658 84742 210894
rect 84186 210338 84422 210574
rect 84506 210338 84742 210574
rect 84186 192658 84422 192894
rect 84506 192658 84742 192894
rect 84186 192338 84422 192574
rect 84506 192338 84742 192574
rect 84186 174658 84422 174894
rect 84506 174658 84742 174894
rect 84186 174338 84422 174574
rect 84506 174338 84742 174574
rect 84186 156658 84422 156894
rect 84506 156658 84742 156894
rect 84186 156338 84422 156574
rect 84506 156338 84742 156574
rect 84186 138658 84422 138894
rect 84506 138658 84742 138894
rect 84186 138338 84422 138574
rect 84506 138338 84742 138574
rect 84186 120658 84422 120894
rect 84506 120658 84742 120894
rect 84186 120338 84422 120574
rect 84506 120338 84742 120574
rect 84186 102658 84422 102894
rect 84506 102658 84742 102894
rect 84186 102338 84422 102574
rect 84506 102338 84742 102574
rect 84186 84658 84422 84894
rect 84506 84658 84742 84894
rect 84186 84338 84422 84574
rect 84506 84338 84742 84574
rect 84186 66658 84422 66894
rect 84506 66658 84742 66894
rect 84186 66338 84422 66574
rect 84506 66338 84742 66574
rect 84186 48658 84422 48894
rect 84506 48658 84742 48894
rect 84186 48338 84422 48574
rect 84506 48338 84742 48574
rect 84186 30658 84422 30894
rect 84506 30658 84742 30894
rect 84186 30338 84422 30574
rect 84506 30338 84742 30574
rect 84186 12658 84422 12894
rect 84506 12658 84742 12894
rect 84186 12338 84422 12574
rect 84506 12338 84742 12574
rect 84186 -3012 84422 -2776
rect 84506 -3012 84742 -2776
rect 84186 -3332 84422 -3096
rect 84506 -3332 84742 -3096
rect 87906 463736 88142 463972
rect 88226 463736 88462 463972
rect 87906 463416 88142 463652
rect 88226 463416 88462 463652
rect 87906 448378 88142 448614
rect 88226 448378 88462 448614
rect 87906 448058 88142 448294
rect 88226 448058 88462 448294
rect 87906 430378 88142 430614
rect 88226 430378 88462 430614
rect 87906 430058 88142 430294
rect 88226 430058 88462 430294
rect 87906 412378 88142 412614
rect 88226 412378 88462 412614
rect 87906 412058 88142 412294
rect 88226 412058 88462 412294
rect 87906 394378 88142 394614
rect 88226 394378 88462 394614
rect 87906 394058 88142 394294
rect 88226 394058 88462 394294
rect 87906 376378 88142 376614
rect 88226 376378 88462 376614
rect 87906 376058 88142 376294
rect 88226 376058 88462 376294
rect 87906 358378 88142 358614
rect 88226 358378 88462 358614
rect 87906 358058 88142 358294
rect 88226 358058 88462 358294
rect 87906 340378 88142 340614
rect 88226 340378 88462 340614
rect 87906 340058 88142 340294
rect 88226 340058 88462 340294
rect 87906 322378 88142 322614
rect 88226 322378 88462 322614
rect 87906 322058 88142 322294
rect 88226 322058 88462 322294
rect 87906 304378 88142 304614
rect 88226 304378 88462 304614
rect 87906 304058 88142 304294
rect 88226 304058 88462 304294
rect 87906 286378 88142 286614
rect 88226 286378 88462 286614
rect 87906 286058 88142 286294
rect 88226 286058 88462 286294
rect 87906 268378 88142 268614
rect 88226 268378 88462 268614
rect 87906 268058 88142 268294
rect 88226 268058 88462 268294
rect 87906 250378 88142 250614
rect 88226 250378 88462 250614
rect 87906 250058 88142 250294
rect 88226 250058 88462 250294
rect 87906 232378 88142 232614
rect 88226 232378 88462 232614
rect 87906 232058 88142 232294
rect 88226 232058 88462 232294
rect 87906 214378 88142 214614
rect 88226 214378 88462 214614
rect 87906 214058 88142 214294
rect 88226 214058 88462 214294
rect 87906 196378 88142 196614
rect 88226 196378 88462 196614
rect 87906 196058 88142 196294
rect 88226 196058 88462 196294
rect 87906 178378 88142 178614
rect 88226 178378 88462 178614
rect 87906 178058 88142 178294
rect 88226 178058 88462 178294
rect 87906 160378 88142 160614
rect 88226 160378 88462 160614
rect 87906 160058 88142 160294
rect 88226 160058 88462 160294
rect 87906 142378 88142 142614
rect 88226 142378 88462 142614
rect 87906 142058 88142 142294
rect 88226 142058 88462 142294
rect 87906 124378 88142 124614
rect 88226 124378 88462 124614
rect 87906 124058 88142 124294
rect 88226 124058 88462 124294
rect 87906 106378 88142 106614
rect 88226 106378 88462 106614
rect 87906 106058 88142 106294
rect 88226 106058 88462 106294
rect 87906 88378 88142 88614
rect 88226 88378 88462 88614
rect 87906 88058 88142 88294
rect 88226 88058 88462 88294
rect 87906 70378 88142 70614
rect 88226 70378 88462 70614
rect 87906 70058 88142 70294
rect 88226 70058 88462 70294
rect 94746 460856 94982 461092
rect 95066 460856 95302 461092
rect 94746 460536 94982 460772
rect 95066 460536 95302 460772
rect 94746 455218 94982 455454
rect 95066 455218 95302 455454
rect 94746 454898 94982 455134
rect 95066 454898 95302 455134
rect 94746 437218 94982 437454
rect 95066 437218 95302 437454
rect 94746 436898 94982 437134
rect 95066 436898 95302 437134
rect 94746 419218 94982 419454
rect 95066 419218 95302 419454
rect 94746 418898 94982 419134
rect 95066 418898 95302 419134
rect 94746 401218 94982 401454
rect 95066 401218 95302 401454
rect 94746 400898 94982 401134
rect 95066 400898 95302 401134
rect 94746 383218 94982 383454
rect 95066 383218 95302 383454
rect 94746 382898 94982 383134
rect 95066 382898 95302 383134
rect 94746 365218 94982 365454
rect 95066 365218 95302 365454
rect 94746 364898 94982 365134
rect 95066 364898 95302 365134
rect 94746 347218 94982 347454
rect 95066 347218 95302 347454
rect 94746 346898 94982 347134
rect 95066 346898 95302 347134
rect 94746 329218 94982 329454
rect 95066 329218 95302 329454
rect 94746 328898 94982 329134
rect 95066 328898 95302 329134
rect 94746 311218 94982 311454
rect 95066 311218 95302 311454
rect 94746 310898 94982 311134
rect 95066 310898 95302 311134
rect 94746 293218 94982 293454
rect 95066 293218 95302 293454
rect 94746 292898 94982 293134
rect 95066 292898 95302 293134
rect 94746 275218 94982 275454
rect 95066 275218 95302 275454
rect 94746 274898 94982 275134
rect 95066 274898 95302 275134
rect 94746 257218 94982 257454
rect 95066 257218 95302 257454
rect 94746 256898 94982 257134
rect 95066 256898 95302 257134
rect 94746 239218 94982 239454
rect 95066 239218 95302 239454
rect 94746 238898 94982 239134
rect 95066 238898 95302 239134
rect 94746 221218 94982 221454
rect 95066 221218 95302 221454
rect 94746 220898 94982 221134
rect 95066 220898 95302 221134
rect 94746 203218 94982 203454
rect 95066 203218 95302 203454
rect 94746 202898 94982 203134
rect 95066 202898 95302 203134
rect 94746 185218 94982 185454
rect 95066 185218 95302 185454
rect 94746 184898 94982 185134
rect 95066 184898 95302 185134
rect 94746 167218 94982 167454
rect 95066 167218 95302 167454
rect 94746 166898 94982 167134
rect 95066 166898 95302 167134
rect 94746 149218 94982 149454
rect 95066 149218 95302 149454
rect 94746 148898 94982 149134
rect 95066 148898 95302 149134
rect 94746 131218 94982 131454
rect 95066 131218 95302 131454
rect 94746 130898 94982 131134
rect 95066 130898 95302 131134
rect 94746 113218 94982 113454
rect 95066 113218 95302 113454
rect 94746 112898 94982 113134
rect 95066 112898 95302 113134
rect 94746 95218 94982 95454
rect 95066 95218 95302 95454
rect 94746 94898 94982 95134
rect 95066 94898 95302 95134
rect 94746 77218 94982 77454
rect 95066 77218 95302 77454
rect 94746 76898 94982 77134
rect 95066 76898 95302 77134
rect 98466 461816 98702 462052
rect 98786 461816 99022 462052
rect 98466 461496 98702 461732
rect 98786 461496 99022 461732
rect 98466 440938 98702 441174
rect 98786 440938 99022 441174
rect 98466 440618 98702 440854
rect 98786 440618 99022 440854
rect 98466 422938 98702 423174
rect 98786 422938 99022 423174
rect 98466 422618 98702 422854
rect 98786 422618 99022 422854
rect 98466 404938 98702 405174
rect 98786 404938 99022 405174
rect 98466 404618 98702 404854
rect 98786 404618 99022 404854
rect 98466 386938 98702 387174
rect 98786 386938 99022 387174
rect 98466 386618 98702 386854
rect 98786 386618 99022 386854
rect 98466 368938 98702 369174
rect 98786 368938 99022 369174
rect 98466 368618 98702 368854
rect 98786 368618 99022 368854
rect 98466 350938 98702 351174
rect 98786 350938 99022 351174
rect 98466 350618 98702 350854
rect 98786 350618 99022 350854
rect 98466 332938 98702 333174
rect 98786 332938 99022 333174
rect 98466 332618 98702 332854
rect 98786 332618 99022 332854
rect 98466 314938 98702 315174
rect 98786 314938 99022 315174
rect 98466 314618 98702 314854
rect 98786 314618 99022 314854
rect 98466 296938 98702 297174
rect 98786 296938 99022 297174
rect 98466 296618 98702 296854
rect 98786 296618 99022 296854
rect 98466 278938 98702 279174
rect 98786 278938 99022 279174
rect 98466 278618 98702 278854
rect 98786 278618 99022 278854
rect 98466 260938 98702 261174
rect 98786 260938 99022 261174
rect 98466 260618 98702 260854
rect 98786 260618 99022 260854
rect 98466 242938 98702 243174
rect 98786 242938 99022 243174
rect 98466 242618 98702 242854
rect 98786 242618 99022 242854
rect 98466 224938 98702 225174
rect 98786 224938 99022 225174
rect 98466 224618 98702 224854
rect 98786 224618 99022 224854
rect 98466 206938 98702 207174
rect 98786 206938 99022 207174
rect 98466 206618 98702 206854
rect 98786 206618 99022 206854
rect 98466 188938 98702 189174
rect 98786 188938 99022 189174
rect 98466 188618 98702 188854
rect 98786 188618 99022 188854
rect 98466 170938 98702 171174
rect 98786 170938 99022 171174
rect 98466 170618 98702 170854
rect 98786 170618 99022 170854
rect 98466 152938 98702 153174
rect 98786 152938 99022 153174
rect 98466 152618 98702 152854
rect 98786 152618 99022 152854
rect 98466 134938 98702 135174
rect 98786 134938 99022 135174
rect 98466 134618 98702 134854
rect 98786 134618 99022 134854
rect 98466 116938 98702 117174
rect 98786 116938 99022 117174
rect 98466 116618 98702 116854
rect 98786 116618 99022 116854
rect 98466 98938 98702 99174
rect 98786 98938 99022 99174
rect 98466 98618 98702 98854
rect 98786 98618 99022 98854
rect 98466 80938 98702 81174
rect 98786 80938 99022 81174
rect 98466 80618 98702 80854
rect 98786 80618 99022 80854
rect 98466 62938 98702 63174
rect 98786 62938 99022 63174
rect 98466 62618 98702 62854
rect 98786 62618 99022 62854
rect 102186 462776 102422 463012
rect 102506 462776 102742 463012
rect 102186 462456 102422 462692
rect 102506 462456 102742 462692
rect 102186 444658 102422 444894
rect 102506 444658 102742 444894
rect 102186 444338 102422 444574
rect 102506 444338 102742 444574
rect 102186 426658 102422 426894
rect 102506 426658 102742 426894
rect 102186 426338 102422 426574
rect 102506 426338 102742 426574
rect 102186 408658 102422 408894
rect 102506 408658 102742 408894
rect 102186 408338 102422 408574
rect 102506 408338 102742 408574
rect 102186 390658 102422 390894
rect 102506 390658 102742 390894
rect 102186 390338 102422 390574
rect 102506 390338 102742 390574
rect 102186 372658 102422 372894
rect 102506 372658 102742 372894
rect 102186 372338 102422 372574
rect 102506 372338 102742 372574
rect 102186 354658 102422 354894
rect 102506 354658 102742 354894
rect 102186 354338 102422 354574
rect 102506 354338 102742 354574
rect 102186 336658 102422 336894
rect 102506 336658 102742 336894
rect 102186 336338 102422 336574
rect 102506 336338 102742 336574
rect 102186 318658 102422 318894
rect 102506 318658 102742 318894
rect 102186 318338 102422 318574
rect 102506 318338 102742 318574
rect 102186 300658 102422 300894
rect 102506 300658 102742 300894
rect 102186 300338 102422 300574
rect 102506 300338 102742 300574
rect 102186 282658 102422 282894
rect 102506 282658 102742 282894
rect 102186 282338 102422 282574
rect 102506 282338 102742 282574
rect 102186 264658 102422 264894
rect 102506 264658 102742 264894
rect 102186 264338 102422 264574
rect 102506 264338 102742 264574
rect 102186 246658 102422 246894
rect 102506 246658 102742 246894
rect 102186 246338 102422 246574
rect 102506 246338 102742 246574
rect 102186 228658 102422 228894
rect 102506 228658 102742 228894
rect 102186 228338 102422 228574
rect 102506 228338 102742 228574
rect 102186 210658 102422 210894
rect 102506 210658 102742 210894
rect 102186 210338 102422 210574
rect 102506 210338 102742 210574
rect 102186 192658 102422 192894
rect 102506 192658 102742 192894
rect 102186 192338 102422 192574
rect 102506 192338 102742 192574
rect 102186 174658 102422 174894
rect 102506 174658 102742 174894
rect 102186 174338 102422 174574
rect 102506 174338 102742 174574
rect 102186 156658 102422 156894
rect 102506 156658 102742 156894
rect 102186 156338 102422 156574
rect 102506 156338 102742 156574
rect 102186 138658 102422 138894
rect 102506 138658 102742 138894
rect 102186 138338 102422 138574
rect 102506 138338 102742 138574
rect 102186 120658 102422 120894
rect 102506 120658 102742 120894
rect 102186 120338 102422 120574
rect 102506 120338 102742 120574
rect 102186 102658 102422 102894
rect 102506 102658 102742 102894
rect 102186 102338 102422 102574
rect 102506 102338 102742 102574
rect 102186 84658 102422 84894
rect 102506 84658 102742 84894
rect 102186 84338 102422 84574
rect 102506 84338 102742 84574
rect 102186 66658 102422 66894
rect 102506 66658 102742 66894
rect 102186 66338 102422 66574
rect 102506 66338 102742 66574
rect 105906 463736 106142 463972
rect 106226 463736 106462 463972
rect 105906 463416 106142 463652
rect 106226 463416 106462 463652
rect 105906 448378 106142 448614
rect 106226 448378 106462 448614
rect 105906 448058 106142 448294
rect 106226 448058 106462 448294
rect 105906 430378 106142 430614
rect 106226 430378 106462 430614
rect 105906 430058 106142 430294
rect 106226 430058 106462 430294
rect 105906 412378 106142 412614
rect 106226 412378 106462 412614
rect 105906 412058 106142 412294
rect 106226 412058 106462 412294
rect 105906 394378 106142 394614
rect 106226 394378 106462 394614
rect 105906 394058 106142 394294
rect 106226 394058 106462 394294
rect 105906 376378 106142 376614
rect 106226 376378 106462 376614
rect 105906 376058 106142 376294
rect 106226 376058 106462 376294
rect 105906 358378 106142 358614
rect 106226 358378 106462 358614
rect 105906 358058 106142 358294
rect 106226 358058 106462 358294
rect 105906 340378 106142 340614
rect 106226 340378 106462 340614
rect 105906 340058 106142 340294
rect 106226 340058 106462 340294
rect 105906 322378 106142 322614
rect 106226 322378 106462 322614
rect 105906 322058 106142 322294
rect 106226 322058 106462 322294
rect 105906 304378 106142 304614
rect 106226 304378 106462 304614
rect 105906 304058 106142 304294
rect 106226 304058 106462 304294
rect 105906 286378 106142 286614
rect 106226 286378 106462 286614
rect 105906 286058 106142 286294
rect 106226 286058 106462 286294
rect 105906 268378 106142 268614
rect 106226 268378 106462 268614
rect 105906 268058 106142 268294
rect 106226 268058 106462 268294
rect 105906 250378 106142 250614
rect 106226 250378 106462 250614
rect 105906 250058 106142 250294
rect 106226 250058 106462 250294
rect 105906 232378 106142 232614
rect 106226 232378 106462 232614
rect 105906 232058 106142 232294
rect 106226 232058 106462 232294
rect 105906 214378 106142 214614
rect 106226 214378 106462 214614
rect 105906 214058 106142 214294
rect 106226 214058 106462 214294
rect 105906 196378 106142 196614
rect 106226 196378 106462 196614
rect 105906 196058 106142 196294
rect 106226 196058 106462 196294
rect 105906 178378 106142 178614
rect 106226 178378 106462 178614
rect 105906 178058 106142 178294
rect 106226 178058 106462 178294
rect 105906 160378 106142 160614
rect 106226 160378 106462 160614
rect 105906 160058 106142 160294
rect 106226 160058 106462 160294
rect 105906 142378 106142 142614
rect 106226 142378 106462 142614
rect 105906 142058 106142 142294
rect 106226 142058 106462 142294
rect 105906 124378 106142 124614
rect 106226 124378 106462 124614
rect 105906 124058 106142 124294
rect 106226 124058 106462 124294
rect 105906 106378 106142 106614
rect 106226 106378 106462 106614
rect 105906 106058 106142 106294
rect 106226 106058 106462 106294
rect 105906 88378 106142 88614
rect 106226 88378 106462 88614
rect 105906 88058 106142 88294
rect 106226 88058 106462 88294
rect 105906 70378 106142 70614
rect 106226 70378 106462 70614
rect 105906 70058 106142 70294
rect 106226 70058 106462 70294
rect 112746 460856 112982 461092
rect 113066 460856 113302 461092
rect 112746 460536 112982 460772
rect 113066 460536 113302 460772
rect 112746 455218 112982 455454
rect 113066 455218 113302 455454
rect 112746 454898 112982 455134
rect 113066 454898 113302 455134
rect 112746 437218 112982 437454
rect 113066 437218 113302 437454
rect 112746 436898 112982 437134
rect 113066 436898 113302 437134
rect 112746 419218 112982 419454
rect 113066 419218 113302 419454
rect 112746 418898 112982 419134
rect 113066 418898 113302 419134
rect 112746 401218 112982 401454
rect 113066 401218 113302 401454
rect 112746 400898 112982 401134
rect 113066 400898 113302 401134
rect 112746 383218 112982 383454
rect 113066 383218 113302 383454
rect 112746 382898 112982 383134
rect 113066 382898 113302 383134
rect 112746 365218 112982 365454
rect 113066 365218 113302 365454
rect 112746 364898 112982 365134
rect 113066 364898 113302 365134
rect 112746 347218 112982 347454
rect 113066 347218 113302 347454
rect 112746 346898 112982 347134
rect 113066 346898 113302 347134
rect 112746 329218 112982 329454
rect 113066 329218 113302 329454
rect 112746 328898 112982 329134
rect 113066 328898 113302 329134
rect 112746 311218 112982 311454
rect 113066 311218 113302 311454
rect 112746 310898 112982 311134
rect 113066 310898 113302 311134
rect 112746 293218 112982 293454
rect 113066 293218 113302 293454
rect 112746 292898 112982 293134
rect 113066 292898 113302 293134
rect 112746 275218 112982 275454
rect 113066 275218 113302 275454
rect 112746 274898 112982 275134
rect 113066 274898 113302 275134
rect 112746 257218 112982 257454
rect 113066 257218 113302 257454
rect 112746 256898 112982 257134
rect 113066 256898 113302 257134
rect 112746 239218 112982 239454
rect 113066 239218 113302 239454
rect 112746 238898 112982 239134
rect 113066 238898 113302 239134
rect 112746 221218 112982 221454
rect 113066 221218 113302 221454
rect 112746 220898 112982 221134
rect 113066 220898 113302 221134
rect 112746 203218 112982 203454
rect 113066 203218 113302 203454
rect 112746 202898 112982 203134
rect 113066 202898 113302 203134
rect 112746 185218 112982 185454
rect 113066 185218 113302 185454
rect 112746 184898 112982 185134
rect 113066 184898 113302 185134
rect 112746 167218 112982 167454
rect 113066 167218 113302 167454
rect 112746 166898 112982 167134
rect 113066 166898 113302 167134
rect 112746 149218 112982 149454
rect 113066 149218 113302 149454
rect 112746 148898 112982 149134
rect 113066 148898 113302 149134
rect 112746 131218 112982 131454
rect 113066 131218 113302 131454
rect 112746 130898 112982 131134
rect 113066 130898 113302 131134
rect 112746 113218 112982 113454
rect 113066 113218 113302 113454
rect 112746 112898 112982 113134
rect 113066 112898 113302 113134
rect 112746 95218 112982 95454
rect 113066 95218 113302 95454
rect 112746 94898 112982 95134
rect 113066 94898 113302 95134
rect 112746 77218 112982 77454
rect 113066 77218 113302 77454
rect 112746 76898 112982 77134
rect 113066 76898 113302 77134
rect 112746 59218 112982 59454
rect 113066 59218 113302 59454
rect 112746 58898 112982 59134
rect 113066 58898 113302 59134
rect 116466 461816 116702 462052
rect 116786 461816 117022 462052
rect 116466 461496 116702 461732
rect 116786 461496 117022 461732
rect 116466 440938 116702 441174
rect 116786 440938 117022 441174
rect 116466 440618 116702 440854
rect 116786 440618 117022 440854
rect 116466 422938 116702 423174
rect 116786 422938 117022 423174
rect 116466 422618 116702 422854
rect 116786 422618 117022 422854
rect 116466 404938 116702 405174
rect 116786 404938 117022 405174
rect 116466 404618 116702 404854
rect 116786 404618 117022 404854
rect 116466 386938 116702 387174
rect 116786 386938 117022 387174
rect 116466 386618 116702 386854
rect 116786 386618 117022 386854
rect 116466 368938 116702 369174
rect 116786 368938 117022 369174
rect 116466 368618 116702 368854
rect 116786 368618 117022 368854
rect 116466 350938 116702 351174
rect 116786 350938 117022 351174
rect 116466 350618 116702 350854
rect 116786 350618 117022 350854
rect 116466 332938 116702 333174
rect 116786 332938 117022 333174
rect 116466 332618 116702 332854
rect 116786 332618 117022 332854
rect 116466 314938 116702 315174
rect 116786 314938 117022 315174
rect 116466 314618 116702 314854
rect 116786 314618 117022 314854
rect 116466 296938 116702 297174
rect 116786 296938 117022 297174
rect 116466 296618 116702 296854
rect 116786 296618 117022 296854
rect 116466 278938 116702 279174
rect 116786 278938 117022 279174
rect 116466 278618 116702 278854
rect 116786 278618 117022 278854
rect 116466 260938 116702 261174
rect 116786 260938 117022 261174
rect 116466 260618 116702 260854
rect 116786 260618 117022 260854
rect 116466 242938 116702 243174
rect 116786 242938 117022 243174
rect 116466 242618 116702 242854
rect 116786 242618 117022 242854
rect 116466 224938 116702 225174
rect 116786 224938 117022 225174
rect 116466 224618 116702 224854
rect 116786 224618 117022 224854
rect 116466 206938 116702 207174
rect 116786 206938 117022 207174
rect 116466 206618 116702 206854
rect 116786 206618 117022 206854
rect 116466 188938 116702 189174
rect 116786 188938 117022 189174
rect 116466 188618 116702 188854
rect 116786 188618 117022 188854
rect 116466 170938 116702 171174
rect 116786 170938 117022 171174
rect 116466 170618 116702 170854
rect 116786 170618 117022 170854
rect 116466 152938 116702 153174
rect 116786 152938 117022 153174
rect 116466 152618 116702 152854
rect 116786 152618 117022 152854
rect 116466 134938 116702 135174
rect 116786 134938 117022 135174
rect 116466 134618 116702 134854
rect 116786 134618 117022 134854
rect 116466 116938 116702 117174
rect 116786 116938 117022 117174
rect 116466 116618 116702 116854
rect 116786 116618 117022 116854
rect 116466 98938 116702 99174
rect 116786 98938 117022 99174
rect 116466 98618 116702 98854
rect 116786 98618 117022 98854
rect 116466 80938 116702 81174
rect 116786 80938 117022 81174
rect 116466 80618 116702 80854
rect 116786 80618 117022 80854
rect 116466 62938 116702 63174
rect 116786 62938 117022 63174
rect 116466 62618 116702 62854
rect 116786 62618 117022 62854
rect 120186 462776 120422 463012
rect 120506 462776 120742 463012
rect 120186 462456 120422 462692
rect 120506 462456 120742 462692
rect 120186 444658 120422 444894
rect 120506 444658 120742 444894
rect 120186 444338 120422 444574
rect 120506 444338 120742 444574
rect 120186 426658 120422 426894
rect 120506 426658 120742 426894
rect 120186 426338 120422 426574
rect 120506 426338 120742 426574
rect 120186 408658 120422 408894
rect 120506 408658 120742 408894
rect 120186 408338 120422 408574
rect 120506 408338 120742 408574
rect 120186 390658 120422 390894
rect 120506 390658 120742 390894
rect 120186 390338 120422 390574
rect 120506 390338 120742 390574
rect 120186 372658 120422 372894
rect 120506 372658 120742 372894
rect 120186 372338 120422 372574
rect 120506 372338 120742 372574
rect 120186 354658 120422 354894
rect 120506 354658 120742 354894
rect 120186 354338 120422 354574
rect 120506 354338 120742 354574
rect 120186 336658 120422 336894
rect 120506 336658 120742 336894
rect 120186 336338 120422 336574
rect 120506 336338 120742 336574
rect 120186 318658 120422 318894
rect 120506 318658 120742 318894
rect 120186 318338 120422 318574
rect 120506 318338 120742 318574
rect 120186 300658 120422 300894
rect 120506 300658 120742 300894
rect 120186 300338 120422 300574
rect 120506 300338 120742 300574
rect 120186 282658 120422 282894
rect 120506 282658 120742 282894
rect 120186 282338 120422 282574
rect 120506 282338 120742 282574
rect 120186 264658 120422 264894
rect 120506 264658 120742 264894
rect 120186 264338 120422 264574
rect 120506 264338 120742 264574
rect 120186 246658 120422 246894
rect 120506 246658 120742 246894
rect 120186 246338 120422 246574
rect 120506 246338 120742 246574
rect 120186 228658 120422 228894
rect 120506 228658 120742 228894
rect 120186 228338 120422 228574
rect 120506 228338 120742 228574
rect 120186 210658 120422 210894
rect 120506 210658 120742 210894
rect 120186 210338 120422 210574
rect 120506 210338 120742 210574
rect 120186 192658 120422 192894
rect 120506 192658 120742 192894
rect 120186 192338 120422 192574
rect 120506 192338 120742 192574
rect 120186 174658 120422 174894
rect 120506 174658 120742 174894
rect 120186 174338 120422 174574
rect 120506 174338 120742 174574
rect 120186 156658 120422 156894
rect 120506 156658 120742 156894
rect 120186 156338 120422 156574
rect 120506 156338 120742 156574
rect 120186 138658 120422 138894
rect 120506 138658 120742 138894
rect 120186 138338 120422 138574
rect 120506 138338 120742 138574
rect 120186 120658 120422 120894
rect 120506 120658 120742 120894
rect 120186 120338 120422 120574
rect 120506 120338 120742 120574
rect 120186 102658 120422 102894
rect 120506 102658 120742 102894
rect 120186 102338 120422 102574
rect 120506 102338 120742 102574
rect 120186 84658 120422 84894
rect 120506 84658 120742 84894
rect 120186 84338 120422 84574
rect 120506 84338 120742 84574
rect 120186 66658 120422 66894
rect 120506 66658 120742 66894
rect 120186 66338 120422 66574
rect 120506 66338 120742 66574
rect 117734 60212 117970 60298
rect 117734 60148 117820 60212
rect 117820 60148 117884 60212
rect 117884 60148 117970 60212
rect 117734 60062 117970 60148
rect 123906 463736 124142 463972
rect 124226 463736 124462 463972
rect 123906 463416 124142 463652
rect 124226 463416 124462 463652
rect 123906 448378 124142 448614
rect 124226 448378 124462 448614
rect 123906 448058 124142 448294
rect 124226 448058 124462 448294
rect 123906 430378 124142 430614
rect 124226 430378 124462 430614
rect 123906 430058 124142 430294
rect 124226 430058 124462 430294
rect 123906 412378 124142 412614
rect 124226 412378 124462 412614
rect 123906 412058 124142 412294
rect 124226 412058 124462 412294
rect 123906 394378 124142 394614
rect 124226 394378 124462 394614
rect 123906 394058 124142 394294
rect 124226 394058 124462 394294
rect 123906 376378 124142 376614
rect 124226 376378 124462 376614
rect 123906 376058 124142 376294
rect 124226 376058 124462 376294
rect 123906 358378 124142 358614
rect 124226 358378 124462 358614
rect 123906 358058 124142 358294
rect 124226 358058 124462 358294
rect 123906 340378 124142 340614
rect 124226 340378 124462 340614
rect 123906 340058 124142 340294
rect 124226 340058 124462 340294
rect 123906 322378 124142 322614
rect 124226 322378 124462 322614
rect 123906 322058 124142 322294
rect 124226 322058 124462 322294
rect 123906 304378 124142 304614
rect 124226 304378 124462 304614
rect 123906 304058 124142 304294
rect 124226 304058 124462 304294
rect 123906 286378 124142 286614
rect 124226 286378 124462 286614
rect 123906 286058 124142 286294
rect 124226 286058 124462 286294
rect 123906 268378 124142 268614
rect 124226 268378 124462 268614
rect 123906 268058 124142 268294
rect 124226 268058 124462 268294
rect 123906 250378 124142 250614
rect 124226 250378 124462 250614
rect 123906 250058 124142 250294
rect 124226 250058 124462 250294
rect 123906 232378 124142 232614
rect 124226 232378 124462 232614
rect 123906 232058 124142 232294
rect 124226 232058 124462 232294
rect 123906 214378 124142 214614
rect 124226 214378 124462 214614
rect 123906 214058 124142 214294
rect 124226 214058 124462 214294
rect 123906 196378 124142 196614
rect 124226 196378 124462 196614
rect 123906 196058 124142 196294
rect 124226 196058 124462 196294
rect 123906 178378 124142 178614
rect 124226 178378 124462 178614
rect 123906 178058 124142 178294
rect 124226 178058 124462 178294
rect 123906 160378 124142 160614
rect 124226 160378 124462 160614
rect 123906 160058 124142 160294
rect 124226 160058 124462 160294
rect 123906 142378 124142 142614
rect 124226 142378 124462 142614
rect 123906 142058 124142 142294
rect 124226 142058 124462 142294
rect 123906 124378 124142 124614
rect 124226 124378 124462 124614
rect 123906 124058 124142 124294
rect 124226 124058 124462 124294
rect 123906 106378 124142 106614
rect 124226 106378 124462 106614
rect 123906 106058 124142 106294
rect 124226 106058 124462 106294
rect 123906 88378 124142 88614
rect 124226 88378 124462 88614
rect 123906 88058 124142 88294
rect 124226 88058 124462 88294
rect 123906 70378 124142 70614
rect 124226 70378 124462 70614
rect 123906 70058 124142 70294
rect 124226 70058 124462 70294
rect 130746 460856 130982 461092
rect 131066 460856 131302 461092
rect 130746 460536 130982 460772
rect 131066 460536 131302 460772
rect 130746 455218 130982 455454
rect 131066 455218 131302 455454
rect 130746 454898 130982 455134
rect 131066 454898 131302 455134
rect 130746 437218 130982 437454
rect 131066 437218 131302 437454
rect 130746 436898 130982 437134
rect 131066 436898 131302 437134
rect 130746 419218 130982 419454
rect 131066 419218 131302 419454
rect 130746 418898 130982 419134
rect 131066 418898 131302 419134
rect 130746 401218 130982 401454
rect 131066 401218 131302 401454
rect 130746 400898 130982 401134
rect 131066 400898 131302 401134
rect 130746 383218 130982 383454
rect 131066 383218 131302 383454
rect 130746 382898 130982 383134
rect 131066 382898 131302 383134
rect 130746 365218 130982 365454
rect 131066 365218 131302 365454
rect 130746 364898 130982 365134
rect 131066 364898 131302 365134
rect 130746 347218 130982 347454
rect 131066 347218 131302 347454
rect 130746 346898 130982 347134
rect 131066 346898 131302 347134
rect 130746 329218 130982 329454
rect 131066 329218 131302 329454
rect 130746 328898 130982 329134
rect 131066 328898 131302 329134
rect 130746 311218 130982 311454
rect 131066 311218 131302 311454
rect 130746 310898 130982 311134
rect 131066 310898 131302 311134
rect 130746 293218 130982 293454
rect 131066 293218 131302 293454
rect 130746 292898 130982 293134
rect 131066 292898 131302 293134
rect 130746 275218 130982 275454
rect 131066 275218 131302 275454
rect 130746 274898 130982 275134
rect 131066 274898 131302 275134
rect 130746 257218 130982 257454
rect 131066 257218 131302 257454
rect 130746 256898 130982 257134
rect 131066 256898 131302 257134
rect 130746 239218 130982 239454
rect 131066 239218 131302 239454
rect 130746 238898 130982 239134
rect 131066 238898 131302 239134
rect 130746 221218 130982 221454
rect 131066 221218 131302 221454
rect 130746 220898 130982 221134
rect 131066 220898 131302 221134
rect 130746 203218 130982 203454
rect 131066 203218 131302 203454
rect 130746 202898 130982 203134
rect 131066 202898 131302 203134
rect 130746 185218 130982 185454
rect 131066 185218 131302 185454
rect 130746 184898 130982 185134
rect 131066 184898 131302 185134
rect 130746 167218 130982 167454
rect 131066 167218 131302 167454
rect 130746 166898 130982 167134
rect 131066 166898 131302 167134
rect 130746 149218 130982 149454
rect 131066 149218 131302 149454
rect 130746 148898 130982 149134
rect 131066 148898 131302 149134
rect 130746 131218 130982 131454
rect 131066 131218 131302 131454
rect 130746 130898 130982 131134
rect 131066 130898 131302 131134
rect 130746 113218 130982 113454
rect 131066 113218 131302 113454
rect 130746 112898 130982 113134
rect 131066 112898 131302 113134
rect 130746 95218 130982 95454
rect 131066 95218 131302 95454
rect 130746 94898 130982 95134
rect 131066 94898 131302 95134
rect 130746 77218 130982 77454
rect 131066 77218 131302 77454
rect 130746 76898 130982 77134
rect 131066 76898 131302 77134
rect 130746 59218 130982 59454
rect 131066 59218 131302 59454
rect 130746 58898 130982 59134
rect 131066 58898 131302 59134
rect 134466 461816 134702 462052
rect 134786 461816 135022 462052
rect 134466 461496 134702 461732
rect 134786 461496 135022 461732
rect 134466 440938 134702 441174
rect 134786 440938 135022 441174
rect 134466 440618 134702 440854
rect 134786 440618 135022 440854
rect 134466 422938 134702 423174
rect 134786 422938 135022 423174
rect 134466 422618 134702 422854
rect 134786 422618 135022 422854
rect 134466 404938 134702 405174
rect 134786 404938 135022 405174
rect 134466 404618 134702 404854
rect 134786 404618 135022 404854
rect 134466 386938 134702 387174
rect 134786 386938 135022 387174
rect 134466 386618 134702 386854
rect 134786 386618 135022 386854
rect 134466 368938 134702 369174
rect 134786 368938 135022 369174
rect 134466 368618 134702 368854
rect 134786 368618 135022 368854
rect 134466 350938 134702 351174
rect 134786 350938 135022 351174
rect 134466 350618 134702 350854
rect 134786 350618 135022 350854
rect 134466 332938 134702 333174
rect 134786 332938 135022 333174
rect 134466 332618 134702 332854
rect 134786 332618 135022 332854
rect 134466 314938 134702 315174
rect 134786 314938 135022 315174
rect 134466 314618 134702 314854
rect 134786 314618 135022 314854
rect 134466 296938 134702 297174
rect 134786 296938 135022 297174
rect 134466 296618 134702 296854
rect 134786 296618 135022 296854
rect 134466 278938 134702 279174
rect 134786 278938 135022 279174
rect 134466 278618 134702 278854
rect 134786 278618 135022 278854
rect 134466 260938 134702 261174
rect 134786 260938 135022 261174
rect 134466 260618 134702 260854
rect 134786 260618 135022 260854
rect 134466 242938 134702 243174
rect 134786 242938 135022 243174
rect 134466 242618 134702 242854
rect 134786 242618 135022 242854
rect 134466 224938 134702 225174
rect 134786 224938 135022 225174
rect 134466 224618 134702 224854
rect 134786 224618 135022 224854
rect 134466 206938 134702 207174
rect 134786 206938 135022 207174
rect 134466 206618 134702 206854
rect 134786 206618 135022 206854
rect 134466 188938 134702 189174
rect 134786 188938 135022 189174
rect 134466 188618 134702 188854
rect 134786 188618 135022 188854
rect 134466 170938 134702 171174
rect 134786 170938 135022 171174
rect 134466 170618 134702 170854
rect 134786 170618 135022 170854
rect 134466 152938 134702 153174
rect 134786 152938 135022 153174
rect 134466 152618 134702 152854
rect 134786 152618 135022 152854
rect 134466 134938 134702 135174
rect 134786 134938 135022 135174
rect 134466 134618 134702 134854
rect 134786 134618 135022 134854
rect 134466 116938 134702 117174
rect 134786 116938 135022 117174
rect 134466 116618 134702 116854
rect 134786 116618 135022 116854
rect 134466 98938 134702 99174
rect 134786 98938 135022 99174
rect 134466 98618 134702 98854
rect 134786 98618 135022 98854
rect 134466 80938 134702 81174
rect 134786 80938 135022 81174
rect 134466 80618 134702 80854
rect 134786 80618 135022 80854
rect 134466 62938 134702 63174
rect 134786 62938 135022 63174
rect 134466 62618 134702 62854
rect 134786 62618 135022 62854
rect 87906 52378 88142 52614
rect 88226 52378 88462 52614
rect 87906 52058 88142 52294
rect 88226 52058 88462 52294
rect 95830 44938 96066 45174
rect 95830 44618 96066 44854
rect 126550 44938 126786 45174
rect 126550 44618 126786 44854
rect 134466 44938 134702 45174
rect 134786 44938 135022 45174
rect 134466 44618 134702 44854
rect 134786 44618 135022 44854
rect 95170 41218 95406 41454
rect 95170 40898 95406 41134
rect 125890 41218 126126 41454
rect 125890 40898 126126 41134
rect 87906 34378 88142 34614
rect 88226 34378 88462 34614
rect 87906 34058 88142 34294
rect 88226 34058 88462 34294
rect 95830 26938 96066 27174
rect 95830 26618 96066 26854
rect 134466 26938 134702 27174
rect 134786 26938 135022 27174
rect 134466 26618 134702 26854
rect 134786 26618 135022 26854
rect 95170 23218 95406 23454
rect 95170 22898 95406 23134
rect 87906 16378 88142 16614
rect 88226 16378 88462 16614
rect 87906 16058 88142 16294
rect 88226 16058 88462 16294
rect 87906 -3972 88142 -3736
rect 88226 -3972 88462 -3736
rect 87906 -4292 88142 -4056
rect 88226 -4292 88462 -4056
rect 94746 5218 94982 5454
rect 95066 5218 95302 5454
rect 94746 4898 94982 5134
rect 95066 4898 95302 5134
rect 94746 -1092 94982 -856
rect 95066 -1092 95302 -856
rect 94746 -1412 94982 -1176
rect 95066 -1412 95302 -1176
rect 98466 8938 98702 9174
rect 98786 8938 99022 9174
rect 98466 8618 98702 8854
rect 98786 8618 99022 8854
rect 102186 12658 102422 12894
rect 102506 12658 102742 12894
rect 102186 12338 102422 12574
rect 102506 12338 102742 12574
rect 100254 902 100490 1138
rect 98466 -2052 98702 -1816
rect 98786 -2052 99022 -1816
rect 98466 -2372 98702 -2136
rect 98786 -2372 99022 -2136
rect 102186 -3012 102422 -2776
rect 102506 -3012 102742 -2776
rect 102186 -3332 102422 -3096
rect 102506 -3332 102742 -3096
rect 105906 16378 106142 16614
rect 106226 16378 106462 16614
rect 105906 16058 106142 16294
rect 106226 16058 106462 16294
rect 112746 5218 112982 5454
rect 113066 5218 113302 5454
rect 112746 4898 112982 5134
rect 113066 4898 113302 5134
rect 108166 1052 108402 1138
rect 108166 988 108252 1052
rect 108252 988 108316 1052
rect 108316 988 108402 1052
rect 108166 902 108402 988
rect 108902 902 109138 1138
rect 105906 -3972 106142 -3736
rect 106226 -3972 106462 -3736
rect 105906 -4292 106142 -4056
rect 106226 -4292 106462 -4056
rect 112746 -1092 112982 -856
rect 113066 -1092 113302 -856
rect 112746 -1412 112982 -1176
rect 113066 -1412 113302 -1176
rect 116466 8938 116702 9174
rect 116786 8938 117022 9174
rect 116466 8618 116702 8854
rect 116786 8618 117022 8854
rect 116466 -2052 116702 -1816
rect 116786 -2052 117022 -1816
rect 116466 -2372 116702 -2136
rect 116786 -2372 117022 -2136
rect 120186 12658 120422 12894
rect 120506 12658 120742 12894
rect 120186 12338 120422 12574
rect 120506 12338 120742 12574
rect 120186 -3012 120422 -2776
rect 120506 -3012 120742 -2776
rect 120186 -3332 120422 -3096
rect 120506 -3332 120742 -3096
rect 123906 16378 124142 16614
rect 124226 16378 124462 16614
rect 123906 16058 124142 16294
rect 124226 16058 124462 16294
rect 123906 -3972 124142 -3736
rect 124226 -3972 124462 -3736
rect 123906 -4292 124142 -4056
rect 124226 -4292 124462 -4056
rect 130746 5218 130982 5454
rect 131066 5218 131302 5454
rect 130746 4898 130982 5134
rect 131066 4898 131302 5134
rect 130746 -1092 130982 -856
rect 131066 -1092 131302 -856
rect 130746 -1412 130982 -1176
rect 131066 -1412 131302 -1176
rect 134466 8938 134702 9174
rect 134786 8938 135022 9174
rect 134466 8618 134702 8854
rect 134786 8618 135022 8854
rect 138186 462776 138422 463012
rect 138506 462776 138742 463012
rect 138186 462456 138422 462692
rect 138506 462456 138742 462692
rect 138186 444658 138422 444894
rect 138506 444658 138742 444894
rect 138186 444338 138422 444574
rect 138506 444338 138742 444574
rect 138186 426658 138422 426894
rect 138506 426658 138742 426894
rect 138186 426338 138422 426574
rect 138506 426338 138742 426574
rect 138186 408658 138422 408894
rect 138506 408658 138742 408894
rect 138186 408338 138422 408574
rect 138506 408338 138742 408574
rect 138186 390658 138422 390894
rect 138506 390658 138742 390894
rect 138186 390338 138422 390574
rect 138506 390338 138742 390574
rect 138186 372658 138422 372894
rect 138506 372658 138742 372894
rect 138186 372338 138422 372574
rect 138506 372338 138742 372574
rect 138186 354658 138422 354894
rect 138506 354658 138742 354894
rect 138186 354338 138422 354574
rect 138506 354338 138742 354574
rect 138186 336658 138422 336894
rect 138506 336658 138742 336894
rect 138186 336338 138422 336574
rect 138506 336338 138742 336574
rect 138186 318658 138422 318894
rect 138506 318658 138742 318894
rect 138186 318338 138422 318574
rect 138506 318338 138742 318574
rect 138186 300658 138422 300894
rect 138506 300658 138742 300894
rect 138186 300338 138422 300574
rect 138506 300338 138742 300574
rect 138186 282658 138422 282894
rect 138506 282658 138742 282894
rect 138186 282338 138422 282574
rect 138506 282338 138742 282574
rect 138186 264658 138422 264894
rect 138506 264658 138742 264894
rect 138186 264338 138422 264574
rect 138506 264338 138742 264574
rect 138186 246658 138422 246894
rect 138506 246658 138742 246894
rect 138186 246338 138422 246574
rect 138506 246338 138742 246574
rect 138186 228658 138422 228894
rect 138506 228658 138742 228894
rect 138186 228338 138422 228574
rect 138506 228338 138742 228574
rect 138186 210658 138422 210894
rect 138506 210658 138742 210894
rect 138186 210338 138422 210574
rect 138506 210338 138742 210574
rect 138186 192658 138422 192894
rect 138506 192658 138742 192894
rect 138186 192338 138422 192574
rect 138506 192338 138742 192574
rect 138186 174658 138422 174894
rect 138506 174658 138742 174894
rect 138186 174338 138422 174574
rect 138506 174338 138742 174574
rect 138186 156658 138422 156894
rect 138506 156658 138742 156894
rect 138186 156338 138422 156574
rect 138506 156338 138742 156574
rect 138186 138658 138422 138894
rect 138506 138658 138742 138894
rect 138186 138338 138422 138574
rect 138506 138338 138742 138574
rect 138186 120658 138422 120894
rect 138506 120658 138742 120894
rect 138186 120338 138422 120574
rect 138506 120338 138742 120574
rect 138186 102658 138422 102894
rect 138506 102658 138742 102894
rect 138186 102338 138422 102574
rect 138506 102338 138742 102574
rect 138186 84658 138422 84894
rect 138506 84658 138742 84894
rect 138186 84338 138422 84574
rect 138506 84338 138742 84574
rect 138186 66658 138422 66894
rect 138506 66658 138742 66894
rect 138186 66338 138422 66574
rect 138506 66338 138742 66574
rect 138186 48658 138422 48894
rect 138506 48658 138742 48894
rect 138186 48338 138422 48574
rect 138506 48338 138742 48574
rect 138186 30658 138422 30894
rect 138506 30658 138742 30894
rect 138186 30338 138422 30574
rect 138506 30338 138742 30574
rect 138186 12658 138422 12894
rect 138506 12658 138742 12894
rect 138186 12338 138422 12574
rect 138506 12338 138742 12574
rect 137422 1052 137658 1138
rect 137422 988 137508 1052
rect 137508 988 137572 1052
rect 137572 988 137658 1052
rect 137422 902 137658 988
rect 137790 222 138026 458
rect 134466 -2052 134702 -1816
rect 134786 -2052 135022 -1816
rect 134466 -2372 134702 -2136
rect 134786 -2372 135022 -2136
rect 138186 -3012 138422 -2776
rect 138506 -3012 138742 -2776
rect 138186 -3332 138422 -3096
rect 138506 -3332 138742 -3096
rect 141906 463736 142142 463972
rect 142226 463736 142462 463972
rect 141906 463416 142142 463652
rect 142226 463416 142462 463652
rect 141906 448378 142142 448614
rect 142226 448378 142462 448614
rect 141906 448058 142142 448294
rect 142226 448058 142462 448294
rect 141906 430378 142142 430614
rect 142226 430378 142462 430614
rect 141906 430058 142142 430294
rect 142226 430058 142462 430294
rect 141906 412378 142142 412614
rect 142226 412378 142462 412614
rect 141906 412058 142142 412294
rect 142226 412058 142462 412294
rect 141906 394378 142142 394614
rect 142226 394378 142462 394614
rect 141906 394058 142142 394294
rect 142226 394058 142462 394294
rect 141906 376378 142142 376614
rect 142226 376378 142462 376614
rect 141906 376058 142142 376294
rect 142226 376058 142462 376294
rect 141906 358378 142142 358614
rect 142226 358378 142462 358614
rect 141906 358058 142142 358294
rect 142226 358058 142462 358294
rect 141906 340378 142142 340614
rect 142226 340378 142462 340614
rect 141906 340058 142142 340294
rect 142226 340058 142462 340294
rect 141906 322378 142142 322614
rect 142226 322378 142462 322614
rect 141906 322058 142142 322294
rect 142226 322058 142462 322294
rect 141906 304378 142142 304614
rect 142226 304378 142462 304614
rect 141906 304058 142142 304294
rect 142226 304058 142462 304294
rect 141906 286378 142142 286614
rect 142226 286378 142462 286614
rect 141906 286058 142142 286294
rect 142226 286058 142462 286294
rect 141906 268378 142142 268614
rect 142226 268378 142462 268614
rect 141906 268058 142142 268294
rect 142226 268058 142462 268294
rect 141906 250378 142142 250614
rect 142226 250378 142462 250614
rect 141906 250058 142142 250294
rect 142226 250058 142462 250294
rect 141906 232378 142142 232614
rect 142226 232378 142462 232614
rect 141906 232058 142142 232294
rect 142226 232058 142462 232294
rect 141906 214378 142142 214614
rect 142226 214378 142462 214614
rect 141906 214058 142142 214294
rect 142226 214058 142462 214294
rect 141906 196378 142142 196614
rect 142226 196378 142462 196614
rect 141906 196058 142142 196294
rect 142226 196058 142462 196294
rect 141906 178378 142142 178614
rect 142226 178378 142462 178614
rect 141906 178058 142142 178294
rect 142226 178058 142462 178294
rect 141906 160378 142142 160614
rect 142226 160378 142462 160614
rect 141906 160058 142142 160294
rect 142226 160058 142462 160294
rect 141906 142378 142142 142614
rect 142226 142378 142462 142614
rect 141906 142058 142142 142294
rect 142226 142058 142462 142294
rect 141906 124378 142142 124614
rect 142226 124378 142462 124614
rect 141906 124058 142142 124294
rect 142226 124058 142462 124294
rect 141906 106378 142142 106614
rect 142226 106378 142462 106614
rect 141906 106058 142142 106294
rect 142226 106058 142462 106294
rect 141906 88378 142142 88614
rect 142226 88378 142462 88614
rect 141906 88058 142142 88294
rect 142226 88058 142462 88294
rect 141906 70378 142142 70614
rect 142226 70378 142462 70614
rect 141906 70058 142142 70294
rect 142226 70058 142462 70294
rect 141906 52378 142142 52614
rect 142226 52378 142462 52614
rect 141906 52058 142142 52294
rect 142226 52058 142462 52294
rect 141906 34378 142142 34614
rect 142226 34378 142462 34614
rect 141906 34058 142142 34294
rect 142226 34058 142462 34294
rect 141906 16378 142142 16614
rect 142226 16378 142462 16614
rect 141906 16058 142142 16294
rect 142226 16058 142462 16294
rect 141906 -3972 142142 -3736
rect 142226 -3972 142462 -3736
rect 141906 -4292 142142 -4056
rect 142226 -4292 142462 -4056
rect 148746 460856 148982 461092
rect 149066 460856 149302 461092
rect 148746 460536 148982 460772
rect 149066 460536 149302 460772
rect 148746 455218 148982 455454
rect 149066 455218 149302 455454
rect 148746 454898 148982 455134
rect 149066 454898 149302 455134
rect 148746 437218 148982 437454
rect 149066 437218 149302 437454
rect 148746 436898 148982 437134
rect 149066 436898 149302 437134
rect 148746 419218 148982 419454
rect 149066 419218 149302 419454
rect 148746 418898 148982 419134
rect 149066 418898 149302 419134
rect 148746 401218 148982 401454
rect 149066 401218 149302 401454
rect 148746 400898 148982 401134
rect 149066 400898 149302 401134
rect 148746 383218 148982 383454
rect 149066 383218 149302 383454
rect 148746 382898 148982 383134
rect 149066 382898 149302 383134
rect 148746 365218 148982 365454
rect 149066 365218 149302 365454
rect 148746 364898 148982 365134
rect 149066 364898 149302 365134
rect 148746 347218 148982 347454
rect 149066 347218 149302 347454
rect 148746 346898 148982 347134
rect 149066 346898 149302 347134
rect 148746 329218 148982 329454
rect 149066 329218 149302 329454
rect 148746 328898 148982 329134
rect 149066 328898 149302 329134
rect 148746 311218 148982 311454
rect 149066 311218 149302 311454
rect 148746 310898 148982 311134
rect 149066 310898 149302 311134
rect 148746 293218 148982 293454
rect 149066 293218 149302 293454
rect 148746 292898 148982 293134
rect 149066 292898 149302 293134
rect 148746 275218 148982 275454
rect 149066 275218 149302 275454
rect 148746 274898 148982 275134
rect 149066 274898 149302 275134
rect 148746 257218 148982 257454
rect 149066 257218 149302 257454
rect 148746 256898 148982 257134
rect 149066 256898 149302 257134
rect 148746 239218 148982 239454
rect 149066 239218 149302 239454
rect 148746 238898 148982 239134
rect 149066 238898 149302 239134
rect 148746 221218 148982 221454
rect 149066 221218 149302 221454
rect 148746 220898 148982 221134
rect 149066 220898 149302 221134
rect 148746 203218 148982 203454
rect 149066 203218 149302 203454
rect 148746 202898 148982 203134
rect 149066 202898 149302 203134
rect 148746 185218 148982 185454
rect 149066 185218 149302 185454
rect 148746 184898 148982 185134
rect 149066 184898 149302 185134
rect 148746 167218 148982 167454
rect 149066 167218 149302 167454
rect 148746 166898 148982 167134
rect 149066 166898 149302 167134
rect 148746 149218 148982 149454
rect 149066 149218 149302 149454
rect 148746 148898 148982 149134
rect 149066 148898 149302 149134
rect 148746 131218 148982 131454
rect 149066 131218 149302 131454
rect 148746 130898 148982 131134
rect 149066 130898 149302 131134
rect 148746 113218 148982 113454
rect 149066 113218 149302 113454
rect 148746 112898 148982 113134
rect 149066 112898 149302 113134
rect 148746 95218 148982 95454
rect 149066 95218 149302 95454
rect 148746 94898 148982 95134
rect 149066 94898 149302 95134
rect 148746 77218 148982 77454
rect 149066 77218 149302 77454
rect 148746 76898 148982 77134
rect 149066 76898 149302 77134
rect 148746 59218 148982 59454
rect 149066 59218 149302 59454
rect 148746 58898 148982 59134
rect 149066 58898 149302 59134
rect 148746 41218 148982 41454
rect 149066 41218 149302 41454
rect 148746 40898 148982 41134
rect 149066 40898 149302 41134
rect 148746 23218 148982 23454
rect 149066 23218 149302 23454
rect 148746 22898 148982 23134
rect 149066 22898 149302 23134
rect 152466 461816 152702 462052
rect 152786 461816 153022 462052
rect 152466 461496 152702 461732
rect 152786 461496 153022 461732
rect 152466 440938 152702 441174
rect 152786 440938 153022 441174
rect 152466 440618 152702 440854
rect 152786 440618 153022 440854
rect 152466 422938 152702 423174
rect 152786 422938 153022 423174
rect 152466 422618 152702 422854
rect 152786 422618 153022 422854
rect 152466 404938 152702 405174
rect 152786 404938 153022 405174
rect 152466 404618 152702 404854
rect 152786 404618 153022 404854
rect 152466 386938 152702 387174
rect 152786 386938 153022 387174
rect 152466 386618 152702 386854
rect 152786 386618 153022 386854
rect 152466 368938 152702 369174
rect 152786 368938 153022 369174
rect 152466 368618 152702 368854
rect 152786 368618 153022 368854
rect 152466 350938 152702 351174
rect 152786 350938 153022 351174
rect 152466 350618 152702 350854
rect 152786 350618 153022 350854
rect 152466 332938 152702 333174
rect 152786 332938 153022 333174
rect 152466 332618 152702 332854
rect 152786 332618 153022 332854
rect 152466 314938 152702 315174
rect 152786 314938 153022 315174
rect 152466 314618 152702 314854
rect 152786 314618 153022 314854
rect 152466 296938 152702 297174
rect 152786 296938 153022 297174
rect 152466 296618 152702 296854
rect 152786 296618 153022 296854
rect 152466 278938 152702 279174
rect 152786 278938 153022 279174
rect 152466 278618 152702 278854
rect 152786 278618 153022 278854
rect 152466 260938 152702 261174
rect 152786 260938 153022 261174
rect 152466 260618 152702 260854
rect 152786 260618 153022 260854
rect 152466 242938 152702 243174
rect 152786 242938 153022 243174
rect 152466 242618 152702 242854
rect 152786 242618 153022 242854
rect 152466 224938 152702 225174
rect 152786 224938 153022 225174
rect 152466 224618 152702 224854
rect 152786 224618 153022 224854
rect 152466 206938 152702 207174
rect 152786 206938 153022 207174
rect 152466 206618 152702 206854
rect 152786 206618 153022 206854
rect 152466 188938 152702 189174
rect 152786 188938 153022 189174
rect 152466 188618 152702 188854
rect 152786 188618 153022 188854
rect 152466 170938 152702 171174
rect 152786 170938 153022 171174
rect 152466 170618 152702 170854
rect 152786 170618 153022 170854
rect 152466 152938 152702 153174
rect 152786 152938 153022 153174
rect 152466 152618 152702 152854
rect 152786 152618 153022 152854
rect 152466 134938 152702 135174
rect 152786 134938 153022 135174
rect 152466 134618 152702 134854
rect 152786 134618 153022 134854
rect 152466 116938 152702 117174
rect 152786 116938 153022 117174
rect 152466 116618 152702 116854
rect 152786 116618 153022 116854
rect 152466 98938 152702 99174
rect 152786 98938 153022 99174
rect 152466 98618 152702 98854
rect 152786 98618 153022 98854
rect 152466 80938 152702 81174
rect 152786 80938 153022 81174
rect 152466 80618 152702 80854
rect 152786 80618 153022 80854
rect 152466 62938 152702 63174
rect 152786 62938 153022 63174
rect 152466 62618 152702 62854
rect 152786 62618 153022 62854
rect 156186 462776 156422 463012
rect 156506 462776 156742 463012
rect 156186 462456 156422 462692
rect 156506 462456 156742 462692
rect 156186 444658 156422 444894
rect 156506 444658 156742 444894
rect 156186 444338 156422 444574
rect 156506 444338 156742 444574
rect 156186 426658 156422 426894
rect 156506 426658 156742 426894
rect 156186 426338 156422 426574
rect 156506 426338 156742 426574
rect 156186 408658 156422 408894
rect 156506 408658 156742 408894
rect 156186 408338 156422 408574
rect 156506 408338 156742 408574
rect 156186 390658 156422 390894
rect 156506 390658 156742 390894
rect 156186 390338 156422 390574
rect 156506 390338 156742 390574
rect 156186 372658 156422 372894
rect 156506 372658 156742 372894
rect 156186 372338 156422 372574
rect 156506 372338 156742 372574
rect 156186 354658 156422 354894
rect 156506 354658 156742 354894
rect 156186 354338 156422 354574
rect 156506 354338 156742 354574
rect 156186 336658 156422 336894
rect 156506 336658 156742 336894
rect 156186 336338 156422 336574
rect 156506 336338 156742 336574
rect 156186 318658 156422 318894
rect 156506 318658 156742 318894
rect 156186 318338 156422 318574
rect 156506 318338 156742 318574
rect 156186 300658 156422 300894
rect 156506 300658 156742 300894
rect 156186 300338 156422 300574
rect 156506 300338 156742 300574
rect 156186 282658 156422 282894
rect 156506 282658 156742 282894
rect 156186 282338 156422 282574
rect 156506 282338 156742 282574
rect 156186 264658 156422 264894
rect 156506 264658 156742 264894
rect 156186 264338 156422 264574
rect 156506 264338 156742 264574
rect 156186 246658 156422 246894
rect 156506 246658 156742 246894
rect 156186 246338 156422 246574
rect 156506 246338 156742 246574
rect 156186 228658 156422 228894
rect 156506 228658 156742 228894
rect 156186 228338 156422 228574
rect 156506 228338 156742 228574
rect 156186 210658 156422 210894
rect 156506 210658 156742 210894
rect 156186 210338 156422 210574
rect 156506 210338 156742 210574
rect 156186 192658 156422 192894
rect 156506 192658 156742 192894
rect 156186 192338 156422 192574
rect 156506 192338 156742 192574
rect 156186 174658 156422 174894
rect 156506 174658 156742 174894
rect 156186 174338 156422 174574
rect 156506 174338 156742 174574
rect 156186 156658 156422 156894
rect 156506 156658 156742 156894
rect 156186 156338 156422 156574
rect 156506 156338 156742 156574
rect 156186 138658 156422 138894
rect 156506 138658 156742 138894
rect 156186 138338 156422 138574
rect 156506 138338 156742 138574
rect 156186 120658 156422 120894
rect 156506 120658 156742 120894
rect 156186 120338 156422 120574
rect 156506 120338 156742 120574
rect 156186 102658 156422 102894
rect 156506 102658 156742 102894
rect 156186 102338 156422 102574
rect 156506 102338 156742 102574
rect 156186 84658 156422 84894
rect 156506 84658 156742 84894
rect 156186 84338 156422 84574
rect 156506 84338 156742 84574
rect 156186 66658 156422 66894
rect 156506 66658 156742 66894
rect 156186 66338 156422 66574
rect 156506 66338 156742 66574
rect 159906 463736 160142 463972
rect 160226 463736 160462 463972
rect 159906 463416 160142 463652
rect 160226 463416 160462 463652
rect 159906 448378 160142 448614
rect 160226 448378 160462 448614
rect 159906 448058 160142 448294
rect 160226 448058 160462 448294
rect 159906 430378 160142 430614
rect 160226 430378 160462 430614
rect 159906 430058 160142 430294
rect 160226 430058 160462 430294
rect 159906 412378 160142 412614
rect 160226 412378 160462 412614
rect 159906 412058 160142 412294
rect 160226 412058 160462 412294
rect 159906 394378 160142 394614
rect 160226 394378 160462 394614
rect 159906 394058 160142 394294
rect 160226 394058 160462 394294
rect 159906 376378 160142 376614
rect 160226 376378 160462 376614
rect 159906 376058 160142 376294
rect 160226 376058 160462 376294
rect 159906 358378 160142 358614
rect 160226 358378 160462 358614
rect 159906 358058 160142 358294
rect 160226 358058 160462 358294
rect 159906 340378 160142 340614
rect 160226 340378 160462 340614
rect 159906 340058 160142 340294
rect 160226 340058 160462 340294
rect 159906 322378 160142 322614
rect 160226 322378 160462 322614
rect 159906 322058 160142 322294
rect 160226 322058 160462 322294
rect 159906 304378 160142 304614
rect 160226 304378 160462 304614
rect 159906 304058 160142 304294
rect 160226 304058 160462 304294
rect 159906 286378 160142 286614
rect 160226 286378 160462 286614
rect 159906 286058 160142 286294
rect 160226 286058 160462 286294
rect 159906 268378 160142 268614
rect 160226 268378 160462 268614
rect 159906 268058 160142 268294
rect 160226 268058 160462 268294
rect 159906 250378 160142 250614
rect 160226 250378 160462 250614
rect 159906 250058 160142 250294
rect 160226 250058 160462 250294
rect 159906 232378 160142 232614
rect 160226 232378 160462 232614
rect 159906 232058 160142 232294
rect 160226 232058 160462 232294
rect 159906 214378 160142 214614
rect 160226 214378 160462 214614
rect 159906 214058 160142 214294
rect 160226 214058 160462 214294
rect 159906 196378 160142 196614
rect 160226 196378 160462 196614
rect 159906 196058 160142 196294
rect 160226 196058 160462 196294
rect 159906 178378 160142 178614
rect 160226 178378 160462 178614
rect 159906 178058 160142 178294
rect 160226 178058 160462 178294
rect 159906 160378 160142 160614
rect 160226 160378 160462 160614
rect 159906 160058 160142 160294
rect 160226 160058 160462 160294
rect 159906 142378 160142 142614
rect 160226 142378 160462 142614
rect 159906 142058 160142 142294
rect 160226 142058 160462 142294
rect 159906 124378 160142 124614
rect 160226 124378 160462 124614
rect 159906 124058 160142 124294
rect 160226 124058 160462 124294
rect 159906 106378 160142 106614
rect 160226 106378 160462 106614
rect 159906 106058 160142 106294
rect 160226 106058 160462 106294
rect 159906 88378 160142 88614
rect 160226 88378 160462 88614
rect 159906 88058 160142 88294
rect 160226 88058 160462 88294
rect 159906 70378 160142 70614
rect 160226 70378 160462 70614
rect 159906 70058 160142 70294
rect 160226 70058 160462 70294
rect 159906 52378 160142 52614
rect 160226 52378 160462 52614
rect 159906 52058 160142 52294
rect 160226 52058 160462 52294
rect 152466 44938 152702 45174
rect 152786 44938 153022 45174
rect 152466 44618 152702 44854
rect 152786 44618 153022 44854
rect 157270 44938 157506 45174
rect 157270 44618 157506 44854
rect 156610 41218 156846 41454
rect 156610 40898 156846 41134
rect 159906 34378 160142 34614
rect 160226 34378 160462 34614
rect 159906 34058 160142 34294
rect 160226 34058 160462 34294
rect 152466 26938 152702 27174
rect 152786 26938 153022 27174
rect 152466 26618 152702 26854
rect 152786 26618 153022 26854
rect 148746 5218 148982 5454
rect 149066 5218 149302 5454
rect 148746 4898 148982 5134
rect 149066 4898 149302 5134
rect 157270 26938 157506 27174
rect 157270 26618 157506 26854
rect 156610 23218 156846 23454
rect 156610 22898 156846 23134
rect 152466 8938 152702 9174
rect 152786 8938 153022 9174
rect 152466 8618 152702 8854
rect 152786 8618 153022 8854
rect 151774 222 152010 458
rect 148746 -1092 148982 -856
rect 149066 -1092 149302 -856
rect 148746 -1412 148982 -1176
rect 149066 -1412 149302 -1176
rect 152466 -2052 152702 -1816
rect 152786 -2052 153022 -1816
rect 152466 -2372 152702 -2136
rect 152786 -2372 153022 -2136
rect 156186 12658 156422 12894
rect 156506 12658 156742 12894
rect 156186 12338 156422 12574
rect 156506 12338 156742 12574
rect 156186 -3012 156422 -2776
rect 156506 -3012 156742 -2776
rect 156186 -3332 156422 -3096
rect 156506 -3332 156742 -3096
rect 159906 16378 160142 16614
rect 160226 16378 160462 16614
rect 159906 16058 160142 16294
rect 160226 16058 160462 16294
rect 159906 -3972 160142 -3736
rect 160226 -3972 160462 -3736
rect 159906 -4292 160142 -4056
rect 160226 -4292 160462 -4056
rect 166746 460856 166982 461092
rect 167066 460856 167302 461092
rect 166746 460536 166982 460772
rect 167066 460536 167302 460772
rect 166746 455218 166982 455454
rect 167066 455218 167302 455454
rect 166746 454898 166982 455134
rect 167066 454898 167302 455134
rect 166746 437218 166982 437454
rect 167066 437218 167302 437454
rect 166746 436898 166982 437134
rect 167066 436898 167302 437134
rect 166746 419218 166982 419454
rect 167066 419218 167302 419454
rect 166746 418898 166982 419134
rect 167066 418898 167302 419134
rect 166746 401218 166982 401454
rect 167066 401218 167302 401454
rect 166746 400898 166982 401134
rect 167066 400898 167302 401134
rect 166746 383218 166982 383454
rect 167066 383218 167302 383454
rect 166746 382898 166982 383134
rect 167066 382898 167302 383134
rect 166746 365218 166982 365454
rect 167066 365218 167302 365454
rect 166746 364898 166982 365134
rect 167066 364898 167302 365134
rect 166746 347218 166982 347454
rect 167066 347218 167302 347454
rect 166746 346898 166982 347134
rect 167066 346898 167302 347134
rect 166746 329218 166982 329454
rect 167066 329218 167302 329454
rect 166746 328898 166982 329134
rect 167066 328898 167302 329134
rect 166746 311218 166982 311454
rect 167066 311218 167302 311454
rect 166746 310898 166982 311134
rect 167066 310898 167302 311134
rect 166746 293218 166982 293454
rect 167066 293218 167302 293454
rect 166746 292898 166982 293134
rect 167066 292898 167302 293134
rect 166746 275218 166982 275454
rect 167066 275218 167302 275454
rect 166746 274898 166982 275134
rect 167066 274898 167302 275134
rect 166746 257218 166982 257454
rect 167066 257218 167302 257454
rect 166746 256898 166982 257134
rect 167066 256898 167302 257134
rect 166746 239218 166982 239454
rect 167066 239218 167302 239454
rect 166746 238898 166982 239134
rect 167066 238898 167302 239134
rect 166746 221218 166982 221454
rect 167066 221218 167302 221454
rect 166746 220898 166982 221134
rect 167066 220898 167302 221134
rect 166746 203218 166982 203454
rect 167066 203218 167302 203454
rect 166746 202898 166982 203134
rect 167066 202898 167302 203134
rect 166746 185218 166982 185454
rect 167066 185218 167302 185454
rect 166746 184898 166982 185134
rect 167066 184898 167302 185134
rect 166746 167218 166982 167454
rect 167066 167218 167302 167454
rect 166746 166898 166982 167134
rect 167066 166898 167302 167134
rect 166746 149218 166982 149454
rect 167066 149218 167302 149454
rect 166746 148898 166982 149134
rect 167066 148898 167302 149134
rect 166746 131218 166982 131454
rect 167066 131218 167302 131454
rect 166746 130898 166982 131134
rect 167066 130898 167302 131134
rect 166746 113218 166982 113454
rect 167066 113218 167302 113454
rect 166746 112898 166982 113134
rect 167066 112898 167302 113134
rect 166746 95218 166982 95454
rect 167066 95218 167302 95454
rect 166746 94898 166982 95134
rect 167066 94898 167302 95134
rect 166746 77218 166982 77454
rect 167066 77218 167302 77454
rect 166746 76898 166982 77134
rect 167066 76898 167302 77134
rect 166746 59218 166982 59454
rect 167066 59218 167302 59454
rect 166746 58898 166982 59134
rect 167066 58898 167302 59134
rect 166746 41218 166982 41454
rect 167066 41218 167302 41454
rect 166746 40898 166982 41134
rect 167066 40898 167302 41134
rect 166746 23218 166982 23454
rect 167066 23218 167302 23454
rect 166746 22898 166982 23134
rect 167066 22898 167302 23134
rect 166746 5218 166982 5454
rect 167066 5218 167302 5454
rect 166746 4898 166982 5134
rect 167066 4898 167302 5134
rect 166746 -1092 166982 -856
rect 167066 -1092 167302 -856
rect 166746 -1412 166982 -1176
rect 167066 -1412 167302 -1176
rect 170466 461816 170702 462052
rect 170786 461816 171022 462052
rect 170466 461496 170702 461732
rect 170786 461496 171022 461732
rect 170466 440938 170702 441174
rect 170786 440938 171022 441174
rect 170466 440618 170702 440854
rect 170786 440618 171022 440854
rect 170466 422938 170702 423174
rect 170786 422938 171022 423174
rect 170466 422618 170702 422854
rect 170786 422618 171022 422854
rect 170466 404938 170702 405174
rect 170786 404938 171022 405174
rect 170466 404618 170702 404854
rect 170786 404618 171022 404854
rect 170466 386938 170702 387174
rect 170786 386938 171022 387174
rect 170466 386618 170702 386854
rect 170786 386618 171022 386854
rect 170466 368938 170702 369174
rect 170786 368938 171022 369174
rect 170466 368618 170702 368854
rect 170786 368618 171022 368854
rect 170466 350938 170702 351174
rect 170786 350938 171022 351174
rect 170466 350618 170702 350854
rect 170786 350618 171022 350854
rect 170466 332938 170702 333174
rect 170786 332938 171022 333174
rect 170466 332618 170702 332854
rect 170786 332618 171022 332854
rect 170466 314938 170702 315174
rect 170786 314938 171022 315174
rect 170466 314618 170702 314854
rect 170786 314618 171022 314854
rect 170466 296938 170702 297174
rect 170786 296938 171022 297174
rect 170466 296618 170702 296854
rect 170786 296618 171022 296854
rect 170466 278938 170702 279174
rect 170786 278938 171022 279174
rect 170466 278618 170702 278854
rect 170786 278618 171022 278854
rect 170466 260938 170702 261174
rect 170786 260938 171022 261174
rect 170466 260618 170702 260854
rect 170786 260618 171022 260854
rect 170466 242938 170702 243174
rect 170786 242938 171022 243174
rect 170466 242618 170702 242854
rect 170786 242618 171022 242854
rect 170466 224938 170702 225174
rect 170786 224938 171022 225174
rect 170466 224618 170702 224854
rect 170786 224618 171022 224854
rect 170466 206938 170702 207174
rect 170786 206938 171022 207174
rect 170466 206618 170702 206854
rect 170786 206618 171022 206854
rect 170466 188938 170702 189174
rect 170786 188938 171022 189174
rect 170466 188618 170702 188854
rect 170786 188618 171022 188854
rect 170466 170938 170702 171174
rect 170786 170938 171022 171174
rect 170466 170618 170702 170854
rect 170786 170618 171022 170854
rect 170466 152938 170702 153174
rect 170786 152938 171022 153174
rect 170466 152618 170702 152854
rect 170786 152618 171022 152854
rect 170466 134938 170702 135174
rect 170786 134938 171022 135174
rect 170466 134618 170702 134854
rect 170786 134618 171022 134854
rect 170466 116938 170702 117174
rect 170786 116938 171022 117174
rect 170466 116618 170702 116854
rect 170786 116618 171022 116854
rect 170466 98938 170702 99174
rect 170786 98938 171022 99174
rect 170466 98618 170702 98854
rect 170786 98618 171022 98854
rect 170466 80938 170702 81174
rect 170786 80938 171022 81174
rect 170466 80618 170702 80854
rect 170786 80618 171022 80854
rect 170466 62938 170702 63174
rect 170786 62938 171022 63174
rect 170466 62618 170702 62854
rect 170786 62618 171022 62854
rect 170466 44938 170702 45174
rect 170786 44938 171022 45174
rect 170466 44618 170702 44854
rect 170786 44618 171022 44854
rect 170466 26938 170702 27174
rect 170786 26938 171022 27174
rect 170466 26618 170702 26854
rect 170786 26618 171022 26854
rect 170466 8938 170702 9174
rect 170786 8938 171022 9174
rect 170466 8618 170702 8854
rect 170786 8618 171022 8854
rect 170466 -2052 170702 -1816
rect 170786 -2052 171022 -1816
rect 170466 -2372 170702 -2136
rect 170786 -2372 171022 -2136
rect 174186 462776 174422 463012
rect 174506 462776 174742 463012
rect 174186 462456 174422 462692
rect 174506 462456 174742 462692
rect 174186 444658 174422 444894
rect 174506 444658 174742 444894
rect 174186 444338 174422 444574
rect 174506 444338 174742 444574
rect 174186 426658 174422 426894
rect 174506 426658 174742 426894
rect 174186 426338 174422 426574
rect 174506 426338 174742 426574
rect 174186 408658 174422 408894
rect 174506 408658 174742 408894
rect 174186 408338 174422 408574
rect 174506 408338 174742 408574
rect 174186 390658 174422 390894
rect 174506 390658 174742 390894
rect 174186 390338 174422 390574
rect 174506 390338 174742 390574
rect 174186 372658 174422 372894
rect 174506 372658 174742 372894
rect 174186 372338 174422 372574
rect 174506 372338 174742 372574
rect 174186 354658 174422 354894
rect 174506 354658 174742 354894
rect 174186 354338 174422 354574
rect 174506 354338 174742 354574
rect 174186 336658 174422 336894
rect 174506 336658 174742 336894
rect 174186 336338 174422 336574
rect 174506 336338 174742 336574
rect 174186 318658 174422 318894
rect 174506 318658 174742 318894
rect 174186 318338 174422 318574
rect 174506 318338 174742 318574
rect 174186 300658 174422 300894
rect 174506 300658 174742 300894
rect 174186 300338 174422 300574
rect 174506 300338 174742 300574
rect 174186 282658 174422 282894
rect 174506 282658 174742 282894
rect 174186 282338 174422 282574
rect 174506 282338 174742 282574
rect 174186 264658 174422 264894
rect 174506 264658 174742 264894
rect 174186 264338 174422 264574
rect 174506 264338 174742 264574
rect 174186 246658 174422 246894
rect 174506 246658 174742 246894
rect 174186 246338 174422 246574
rect 174506 246338 174742 246574
rect 174186 228658 174422 228894
rect 174506 228658 174742 228894
rect 174186 228338 174422 228574
rect 174506 228338 174742 228574
rect 174186 210658 174422 210894
rect 174506 210658 174742 210894
rect 174186 210338 174422 210574
rect 174506 210338 174742 210574
rect 174186 192658 174422 192894
rect 174506 192658 174742 192894
rect 174186 192338 174422 192574
rect 174506 192338 174742 192574
rect 174186 174658 174422 174894
rect 174506 174658 174742 174894
rect 174186 174338 174422 174574
rect 174506 174338 174742 174574
rect 174186 156658 174422 156894
rect 174506 156658 174742 156894
rect 174186 156338 174422 156574
rect 174506 156338 174742 156574
rect 174186 138658 174422 138894
rect 174506 138658 174742 138894
rect 174186 138338 174422 138574
rect 174506 138338 174742 138574
rect 174186 120658 174422 120894
rect 174506 120658 174742 120894
rect 174186 120338 174422 120574
rect 174506 120338 174742 120574
rect 174186 102658 174422 102894
rect 174506 102658 174742 102894
rect 174186 102338 174422 102574
rect 174506 102338 174742 102574
rect 174186 84658 174422 84894
rect 174506 84658 174742 84894
rect 174186 84338 174422 84574
rect 174506 84338 174742 84574
rect 174186 66658 174422 66894
rect 174506 66658 174742 66894
rect 174186 66338 174422 66574
rect 174506 66338 174742 66574
rect 174186 48658 174422 48894
rect 174506 48658 174742 48894
rect 174186 48338 174422 48574
rect 174506 48338 174742 48574
rect 174186 30658 174422 30894
rect 174506 30658 174742 30894
rect 174186 30338 174422 30574
rect 174506 30338 174742 30574
rect 174186 12658 174422 12894
rect 174506 12658 174742 12894
rect 174186 12338 174422 12574
rect 174506 12338 174742 12574
rect 174186 -3012 174422 -2776
rect 174506 -3012 174742 -2776
rect 174186 -3332 174422 -3096
rect 174506 -3332 174742 -3096
rect 177906 463736 178142 463972
rect 178226 463736 178462 463972
rect 177906 463416 178142 463652
rect 178226 463416 178462 463652
rect 177906 448378 178142 448614
rect 178226 448378 178462 448614
rect 177906 448058 178142 448294
rect 178226 448058 178462 448294
rect 177906 430378 178142 430614
rect 178226 430378 178462 430614
rect 177906 430058 178142 430294
rect 178226 430058 178462 430294
rect 177906 412378 178142 412614
rect 178226 412378 178462 412614
rect 177906 412058 178142 412294
rect 178226 412058 178462 412294
rect 177906 394378 178142 394614
rect 178226 394378 178462 394614
rect 177906 394058 178142 394294
rect 178226 394058 178462 394294
rect 177906 376378 178142 376614
rect 178226 376378 178462 376614
rect 177906 376058 178142 376294
rect 178226 376058 178462 376294
rect 177906 358378 178142 358614
rect 178226 358378 178462 358614
rect 177906 358058 178142 358294
rect 178226 358058 178462 358294
rect 177906 340378 178142 340614
rect 178226 340378 178462 340614
rect 177906 340058 178142 340294
rect 178226 340058 178462 340294
rect 177906 322378 178142 322614
rect 178226 322378 178462 322614
rect 177906 322058 178142 322294
rect 178226 322058 178462 322294
rect 177906 304378 178142 304614
rect 178226 304378 178462 304614
rect 177906 304058 178142 304294
rect 178226 304058 178462 304294
rect 177906 286378 178142 286614
rect 178226 286378 178462 286614
rect 177906 286058 178142 286294
rect 178226 286058 178462 286294
rect 177906 268378 178142 268614
rect 178226 268378 178462 268614
rect 177906 268058 178142 268294
rect 178226 268058 178462 268294
rect 177906 250378 178142 250614
rect 178226 250378 178462 250614
rect 177906 250058 178142 250294
rect 178226 250058 178462 250294
rect 177906 232378 178142 232614
rect 178226 232378 178462 232614
rect 177906 232058 178142 232294
rect 178226 232058 178462 232294
rect 177906 214378 178142 214614
rect 178226 214378 178462 214614
rect 177906 214058 178142 214294
rect 178226 214058 178462 214294
rect 177906 196378 178142 196614
rect 178226 196378 178462 196614
rect 177906 196058 178142 196294
rect 178226 196058 178462 196294
rect 177906 178378 178142 178614
rect 178226 178378 178462 178614
rect 177906 178058 178142 178294
rect 178226 178058 178462 178294
rect 177906 160378 178142 160614
rect 178226 160378 178462 160614
rect 177906 160058 178142 160294
rect 178226 160058 178462 160294
rect 177906 142378 178142 142614
rect 178226 142378 178462 142614
rect 177906 142058 178142 142294
rect 178226 142058 178462 142294
rect 177906 124378 178142 124614
rect 178226 124378 178462 124614
rect 177906 124058 178142 124294
rect 178226 124058 178462 124294
rect 177906 106378 178142 106614
rect 178226 106378 178462 106614
rect 177906 106058 178142 106294
rect 178226 106058 178462 106294
rect 177906 88378 178142 88614
rect 178226 88378 178462 88614
rect 177906 88058 178142 88294
rect 178226 88058 178462 88294
rect 177906 70378 178142 70614
rect 178226 70378 178462 70614
rect 177906 70058 178142 70294
rect 178226 70058 178462 70294
rect 177906 52378 178142 52614
rect 178226 52378 178462 52614
rect 177906 52058 178142 52294
rect 178226 52058 178462 52294
rect 177906 34378 178142 34614
rect 178226 34378 178462 34614
rect 177906 34058 178142 34294
rect 178226 34058 178462 34294
rect 177906 16378 178142 16614
rect 178226 16378 178462 16614
rect 177906 16058 178142 16294
rect 178226 16058 178462 16294
rect 177906 -3972 178142 -3736
rect 178226 -3972 178462 -3736
rect 177906 -4292 178142 -4056
rect 178226 -4292 178462 -4056
rect 184746 460856 184982 461092
rect 185066 460856 185302 461092
rect 184746 460536 184982 460772
rect 185066 460536 185302 460772
rect 184746 455218 184982 455454
rect 185066 455218 185302 455454
rect 184746 454898 184982 455134
rect 185066 454898 185302 455134
rect 184746 437218 184982 437454
rect 185066 437218 185302 437454
rect 184746 436898 184982 437134
rect 185066 436898 185302 437134
rect 184746 419218 184982 419454
rect 185066 419218 185302 419454
rect 184746 418898 184982 419134
rect 185066 418898 185302 419134
rect 184746 401218 184982 401454
rect 185066 401218 185302 401454
rect 184746 400898 184982 401134
rect 185066 400898 185302 401134
rect 184746 383218 184982 383454
rect 185066 383218 185302 383454
rect 184746 382898 184982 383134
rect 185066 382898 185302 383134
rect 184746 365218 184982 365454
rect 185066 365218 185302 365454
rect 184746 364898 184982 365134
rect 185066 364898 185302 365134
rect 184746 347218 184982 347454
rect 185066 347218 185302 347454
rect 184746 346898 184982 347134
rect 185066 346898 185302 347134
rect 184746 329218 184982 329454
rect 185066 329218 185302 329454
rect 184746 328898 184982 329134
rect 185066 328898 185302 329134
rect 184746 311218 184982 311454
rect 185066 311218 185302 311454
rect 184746 310898 184982 311134
rect 185066 310898 185302 311134
rect 184746 293218 184982 293454
rect 185066 293218 185302 293454
rect 184746 292898 184982 293134
rect 185066 292898 185302 293134
rect 184746 275218 184982 275454
rect 185066 275218 185302 275454
rect 184746 274898 184982 275134
rect 185066 274898 185302 275134
rect 184746 257218 184982 257454
rect 185066 257218 185302 257454
rect 184746 256898 184982 257134
rect 185066 256898 185302 257134
rect 184746 239218 184982 239454
rect 185066 239218 185302 239454
rect 184746 238898 184982 239134
rect 185066 238898 185302 239134
rect 184746 221218 184982 221454
rect 185066 221218 185302 221454
rect 184746 220898 184982 221134
rect 185066 220898 185302 221134
rect 184746 203218 184982 203454
rect 185066 203218 185302 203454
rect 184746 202898 184982 203134
rect 185066 202898 185302 203134
rect 184746 185218 184982 185454
rect 185066 185218 185302 185454
rect 184746 184898 184982 185134
rect 185066 184898 185302 185134
rect 184746 167218 184982 167454
rect 185066 167218 185302 167454
rect 184746 166898 184982 167134
rect 185066 166898 185302 167134
rect 184746 149218 184982 149454
rect 185066 149218 185302 149454
rect 184746 148898 184982 149134
rect 185066 148898 185302 149134
rect 184746 131218 184982 131454
rect 185066 131218 185302 131454
rect 184746 130898 184982 131134
rect 185066 130898 185302 131134
rect 184746 113218 184982 113454
rect 185066 113218 185302 113454
rect 184746 112898 184982 113134
rect 185066 112898 185302 113134
rect 184746 95218 184982 95454
rect 185066 95218 185302 95454
rect 184746 94898 184982 95134
rect 185066 94898 185302 95134
rect 184746 77218 184982 77454
rect 185066 77218 185302 77454
rect 184746 76898 184982 77134
rect 185066 76898 185302 77134
rect 184746 59218 184982 59454
rect 185066 59218 185302 59454
rect 184746 58898 184982 59134
rect 185066 58898 185302 59134
rect 184746 41218 184982 41454
rect 185066 41218 185302 41454
rect 184746 40898 184982 41134
rect 185066 40898 185302 41134
rect 184746 23218 184982 23454
rect 185066 23218 185302 23454
rect 184746 22898 184982 23134
rect 185066 22898 185302 23134
rect 184746 5218 184982 5454
rect 185066 5218 185302 5454
rect 184746 4898 184982 5134
rect 185066 4898 185302 5134
rect 184746 -1092 184982 -856
rect 185066 -1092 185302 -856
rect 184746 -1412 184982 -1176
rect 185066 -1412 185302 -1176
rect 188466 461816 188702 462052
rect 188786 461816 189022 462052
rect 188466 461496 188702 461732
rect 188786 461496 189022 461732
rect 188466 440938 188702 441174
rect 188786 440938 189022 441174
rect 188466 440618 188702 440854
rect 188786 440618 189022 440854
rect 188466 422938 188702 423174
rect 188786 422938 189022 423174
rect 188466 422618 188702 422854
rect 188786 422618 189022 422854
rect 188466 404938 188702 405174
rect 188786 404938 189022 405174
rect 188466 404618 188702 404854
rect 188786 404618 189022 404854
rect 188466 386938 188702 387174
rect 188786 386938 189022 387174
rect 188466 386618 188702 386854
rect 188786 386618 189022 386854
rect 188466 368938 188702 369174
rect 188786 368938 189022 369174
rect 188466 368618 188702 368854
rect 188786 368618 189022 368854
rect 188466 350938 188702 351174
rect 188786 350938 189022 351174
rect 188466 350618 188702 350854
rect 188786 350618 189022 350854
rect 188466 332938 188702 333174
rect 188786 332938 189022 333174
rect 188466 332618 188702 332854
rect 188786 332618 189022 332854
rect 188466 314938 188702 315174
rect 188786 314938 189022 315174
rect 188466 314618 188702 314854
rect 188786 314618 189022 314854
rect 188466 296938 188702 297174
rect 188786 296938 189022 297174
rect 188466 296618 188702 296854
rect 188786 296618 189022 296854
rect 188466 278938 188702 279174
rect 188786 278938 189022 279174
rect 188466 278618 188702 278854
rect 188786 278618 189022 278854
rect 188466 260938 188702 261174
rect 188786 260938 189022 261174
rect 188466 260618 188702 260854
rect 188786 260618 189022 260854
rect 188466 242938 188702 243174
rect 188786 242938 189022 243174
rect 188466 242618 188702 242854
rect 188786 242618 189022 242854
rect 188466 224938 188702 225174
rect 188786 224938 189022 225174
rect 188466 224618 188702 224854
rect 188786 224618 189022 224854
rect 188466 206938 188702 207174
rect 188786 206938 189022 207174
rect 188466 206618 188702 206854
rect 188786 206618 189022 206854
rect 188466 188938 188702 189174
rect 188786 188938 189022 189174
rect 188466 188618 188702 188854
rect 188786 188618 189022 188854
rect 188466 170938 188702 171174
rect 188786 170938 189022 171174
rect 188466 170618 188702 170854
rect 188786 170618 189022 170854
rect 188466 152938 188702 153174
rect 188786 152938 189022 153174
rect 188466 152618 188702 152854
rect 188786 152618 189022 152854
rect 188466 134938 188702 135174
rect 188786 134938 189022 135174
rect 188466 134618 188702 134854
rect 188786 134618 189022 134854
rect 188466 116938 188702 117174
rect 188786 116938 189022 117174
rect 188466 116618 188702 116854
rect 188786 116618 189022 116854
rect 188466 98938 188702 99174
rect 188786 98938 189022 99174
rect 188466 98618 188702 98854
rect 188786 98618 189022 98854
rect 188466 80938 188702 81174
rect 188786 80938 189022 81174
rect 188466 80618 188702 80854
rect 188786 80618 189022 80854
rect 188466 62938 188702 63174
rect 188786 62938 189022 63174
rect 188466 62618 188702 62854
rect 188786 62618 189022 62854
rect 188466 44938 188702 45174
rect 188786 44938 189022 45174
rect 188466 44618 188702 44854
rect 188786 44618 189022 44854
rect 188466 26938 188702 27174
rect 188786 26938 189022 27174
rect 188466 26618 188702 26854
rect 188786 26618 189022 26854
rect 188466 8938 188702 9174
rect 188786 8938 189022 9174
rect 188466 8618 188702 8854
rect 188786 8618 189022 8854
rect 188466 -2052 188702 -1816
rect 188786 -2052 189022 -1816
rect 188466 -2372 188702 -2136
rect 188786 -2372 189022 -2136
rect 192186 462776 192422 463012
rect 192506 462776 192742 463012
rect 192186 462456 192422 462692
rect 192506 462456 192742 462692
rect 192186 444658 192422 444894
rect 192506 444658 192742 444894
rect 192186 444338 192422 444574
rect 192506 444338 192742 444574
rect 192186 426658 192422 426894
rect 192506 426658 192742 426894
rect 192186 426338 192422 426574
rect 192506 426338 192742 426574
rect 192186 408658 192422 408894
rect 192506 408658 192742 408894
rect 192186 408338 192422 408574
rect 192506 408338 192742 408574
rect 192186 390658 192422 390894
rect 192506 390658 192742 390894
rect 192186 390338 192422 390574
rect 192506 390338 192742 390574
rect 192186 372658 192422 372894
rect 192506 372658 192742 372894
rect 192186 372338 192422 372574
rect 192506 372338 192742 372574
rect 192186 354658 192422 354894
rect 192506 354658 192742 354894
rect 192186 354338 192422 354574
rect 192506 354338 192742 354574
rect 192186 336658 192422 336894
rect 192506 336658 192742 336894
rect 192186 336338 192422 336574
rect 192506 336338 192742 336574
rect 192186 318658 192422 318894
rect 192506 318658 192742 318894
rect 192186 318338 192422 318574
rect 192506 318338 192742 318574
rect 192186 300658 192422 300894
rect 192506 300658 192742 300894
rect 192186 300338 192422 300574
rect 192506 300338 192742 300574
rect 192186 282658 192422 282894
rect 192506 282658 192742 282894
rect 192186 282338 192422 282574
rect 192506 282338 192742 282574
rect 192186 264658 192422 264894
rect 192506 264658 192742 264894
rect 192186 264338 192422 264574
rect 192506 264338 192742 264574
rect 192186 246658 192422 246894
rect 192506 246658 192742 246894
rect 192186 246338 192422 246574
rect 192506 246338 192742 246574
rect 192186 228658 192422 228894
rect 192506 228658 192742 228894
rect 192186 228338 192422 228574
rect 192506 228338 192742 228574
rect 192186 210658 192422 210894
rect 192506 210658 192742 210894
rect 192186 210338 192422 210574
rect 192506 210338 192742 210574
rect 192186 192658 192422 192894
rect 192506 192658 192742 192894
rect 192186 192338 192422 192574
rect 192506 192338 192742 192574
rect 192186 174658 192422 174894
rect 192506 174658 192742 174894
rect 192186 174338 192422 174574
rect 192506 174338 192742 174574
rect 192186 156658 192422 156894
rect 192506 156658 192742 156894
rect 192186 156338 192422 156574
rect 192506 156338 192742 156574
rect 192186 138658 192422 138894
rect 192506 138658 192742 138894
rect 192186 138338 192422 138574
rect 192506 138338 192742 138574
rect 192186 120658 192422 120894
rect 192506 120658 192742 120894
rect 192186 120338 192422 120574
rect 192506 120338 192742 120574
rect 192186 102658 192422 102894
rect 192506 102658 192742 102894
rect 192186 102338 192422 102574
rect 192506 102338 192742 102574
rect 192186 84658 192422 84894
rect 192506 84658 192742 84894
rect 192186 84338 192422 84574
rect 192506 84338 192742 84574
rect 192186 66658 192422 66894
rect 192506 66658 192742 66894
rect 192186 66338 192422 66574
rect 192506 66338 192742 66574
rect 192186 48658 192422 48894
rect 192506 48658 192742 48894
rect 192186 48338 192422 48574
rect 192506 48338 192742 48574
rect 192186 30658 192422 30894
rect 192506 30658 192742 30894
rect 192186 30338 192422 30574
rect 192506 30338 192742 30574
rect 192186 12658 192422 12894
rect 192506 12658 192742 12894
rect 192186 12338 192422 12574
rect 192506 12338 192742 12574
rect 192186 -3012 192422 -2776
rect 192506 -3012 192742 -2776
rect 192186 -3332 192422 -3096
rect 192506 -3332 192742 -3096
rect 195906 463736 196142 463972
rect 196226 463736 196462 463972
rect 195906 463416 196142 463652
rect 196226 463416 196462 463652
rect 195906 448378 196142 448614
rect 196226 448378 196462 448614
rect 195906 448058 196142 448294
rect 196226 448058 196462 448294
rect 195906 430378 196142 430614
rect 196226 430378 196462 430614
rect 195906 430058 196142 430294
rect 196226 430058 196462 430294
rect 195906 412378 196142 412614
rect 196226 412378 196462 412614
rect 195906 412058 196142 412294
rect 196226 412058 196462 412294
rect 195906 394378 196142 394614
rect 196226 394378 196462 394614
rect 195906 394058 196142 394294
rect 196226 394058 196462 394294
rect 195906 376378 196142 376614
rect 196226 376378 196462 376614
rect 195906 376058 196142 376294
rect 196226 376058 196462 376294
rect 195906 358378 196142 358614
rect 196226 358378 196462 358614
rect 195906 358058 196142 358294
rect 196226 358058 196462 358294
rect 195906 340378 196142 340614
rect 196226 340378 196462 340614
rect 195906 340058 196142 340294
rect 196226 340058 196462 340294
rect 195906 322378 196142 322614
rect 196226 322378 196462 322614
rect 195906 322058 196142 322294
rect 196226 322058 196462 322294
rect 195906 304378 196142 304614
rect 196226 304378 196462 304614
rect 195906 304058 196142 304294
rect 196226 304058 196462 304294
rect 195906 286378 196142 286614
rect 196226 286378 196462 286614
rect 195906 286058 196142 286294
rect 196226 286058 196462 286294
rect 195906 268378 196142 268614
rect 196226 268378 196462 268614
rect 195906 268058 196142 268294
rect 196226 268058 196462 268294
rect 195906 250378 196142 250614
rect 196226 250378 196462 250614
rect 195906 250058 196142 250294
rect 196226 250058 196462 250294
rect 195906 232378 196142 232614
rect 196226 232378 196462 232614
rect 195906 232058 196142 232294
rect 196226 232058 196462 232294
rect 195906 214378 196142 214614
rect 196226 214378 196462 214614
rect 195906 214058 196142 214294
rect 196226 214058 196462 214294
rect 195906 196378 196142 196614
rect 196226 196378 196462 196614
rect 195906 196058 196142 196294
rect 196226 196058 196462 196294
rect 195906 178378 196142 178614
rect 196226 178378 196462 178614
rect 195906 178058 196142 178294
rect 196226 178058 196462 178294
rect 195906 160378 196142 160614
rect 196226 160378 196462 160614
rect 195906 160058 196142 160294
rect 196226 160058 196462 160294
rect 195906 142378 196142 142614
rect 196226 142378 196462 142614
rect 195906 142058 196142 142294
rect 196226 142058 196462 142294
rect 195906 124378 196142 124614
rect 196226 124378 196462 124614
rect 195906 124058 196142 124294
rect 196226 124058 196462 124294
rect 195906 106378 196142 106614
rect 196226 106378 196462 106614
rect 195906 106058 196142 106294
rect 196226 106058 196462 106294
rect 195906 88378 196142 88614
rect 196226 88378 196462 88614
rect 195906 88058 196142 88294
rect 196226 88058 196462 88294
rect 195906 70378 196142 70614
rect 196226 70378 196462 70614
rect 195906 70058 196142 70294
rect 196226 70058 196462 70294
rect 195906 52378 196142 52614
rect 196226 52378 196462 52614
rect 195906 52058 196142 52294
rect 196226 52058 196462 52294
rect 195906 34378 196142 34614
rect 196226 34378 196462 34614
rect 195906 34058 196142 34294
rect 196226 34058 196462 34294
rect 195906 16378 196142 16614
rect 196226 16378 196462 16614
rect 195906 16058 196142 16294
rect 196226 16058 196462 16294
rect 195906 -3972 196142 -3736
rect 196226 -3972 196462 -3736
rect 195906 -4292 196142 -4056
rect 196226 -4292 196462 -4056
rect 202746 460856 202982 461092
rect 203066 460856 203302 461092
rect 202746 460536 202982 460772
rect 203066 460536 203302 460772
rect 202746 455218 202982 455454
rect 203066 455218 203302 455454
rect 202746 454898 202982 455134
rect 203066 454898 203302 455134
rect 202746 437218 202982 437454
rect 203066 437218 203302 437454
rect 202746 436898 202982 437134
rect 203066 436898 203302 437134
rect 202746 419218 202982 419454
rect 203066 419218 203302 419454
rect 202746 418898 202982 419134
rect 203066 418898 203302 419134
rect 202746 401218 202982 401454
rect 203066 401218 203302 401454
rect 202746 400898 202982 401134
rect 203066 400898 203302 401134
rect 202746 383218 202982 383454
rect 203066 383218 203302 383454
rect 202746 382898 202982 383134
rect 203066 382898 203302 383134
rect 202746 365218 202982 365454
rect 203066 365218 203302 365454
rect 202746 364898 202982 365134
rect 203066 364898 203302 365134
rect 202746 347218 202982 347454
rect 203066 347218 203302 347454
rect 202746 346898 202982 347134
rect 203066 346898 203302 347134
rect 202746 329218 202982 329454
rect 203066 329218 203302 329454
rect 202746 328898 202982 329134
rect 203066 328898 203302 329134
rect 202746 311218 202982 311454
rect 203066 311218 203302 311454
rect 202746 310898 202982 311134
rect 203066 310898 203302 311134
rect 202746 293218 202982 293454
rect 203066 293218 203302 293454
rect 202746 292898 202982 293134
rect 203066 292898 203302 293134
rect 202746 275218 202982 275454
rect 203066 275218 203302 275454
rect 202746 274898 202982 275134
rect 203066 274898 203302 275134
rect 202746 257218 202982 257454
rect 203066 257218 203302 257454
rect 202746 256898 202982 257134
rect 203066 256898 203302 257134
rect 202746 239218 202982 239454
rect 203066 239218 203302 239454
rect 202746 238898 202982 239134
rect 203066 238898 203302 239134
rect 202746 221218 202982 221454
rect 203066 221218 203302 221454
rect 202746 220898 202982 221134
rect 203066 220898 203302 221134
rect 202746 203218 202982 203454
rect 203066 203218 203302 203454
rect 202746 202898 202982 203134
rect 203066 202898 203302 203134
rect 202746 185218 202982 185454
rect 203066 185218 203302 185454
rect 202746 184898 202982 185134
rect 203066 184898 203302 185134
rect 202746 167218 202982 167454
rect 203066 167218 203302 167454
rect 202746 166898 202982 167134
rect 203066 166898 203302 167134
rect 202746 149218 202982 149454
rect 203066 149218 203302 149454
rect 202746 148898 202982 149134
rect 203066 148898 203302 149134
rect 202746 131218 202982 131454
rect 203066 131218 203302 131454
rect 202746 130898 202982 131134
rect 203066 130898 203302 131134
rect 202746 113218 202982 113454
rect 203066 113218 203302 113454
rect 202746 112898 202982 113134
rect 203066 112898 203302 113134
rect 202746 95218 202982 95454
rect 203066 95218 203302 95454
rect 202746 94898 202982 95134
rect 203066 94898 203302 95134
rect 202746 77218 202982 77454
rect 203066 77218 203302 77454
rect 202746 76898 202982 77134
rect 203066 76898 203302 77134
rect 202746 59218 202982 59454
rect 203066 59218 203302 59454
rect 202746 58898 202982 59134
rect 203066 58898 203302 59134
rect 202746 41218 202982 41454
rect 203066 41218 203302 41454
rect 202746 40898 202982 41134
rect 203066 40898 203302 41134
rect 202746 23218 202982 23454
rect 203066 23218 203302 23454
rect 202746 22898 202982 23134
rect 203066 22898 203302 23134
rect 202746 5218 202982 5454
rect 203066 5218 203302 5454
rect 202746 4898 202982 5134
rect 203066 4898 203302 5134
rect 202746 -1092 202982 -856
rect 203066 -1092 203302 -856
rect 202746 -1412 202982 -1176
rect 203066 -1412 203302 -1176
rect 206466 461816 206702 462052
rect 206786 461816 207022 462052
rect 206466 461496 206702 461732
rect 206786 461496 207022 461732
rect 206466 440938 206702 441174
rect 206786 440938 207022 441174
rect 206466 440618 206702 440854
rect 206786 440618 207022 440854
rect 206466 422938 206702 423174
rect 206786 422938 207022 423174
rect 206466 422618 206702 422854
rect 206786 422618 207022 422854
rect 206466 404938 206702 405174
rect 206786 404938 207022 405174
rect 206466 404618 206702 404854
rect 206786 404618 207022 404854
rect 206466 386938 206702 387174
rect 206786 386938 207022 387174
rect 206466 386618 206702 386854
rect 206786 386618 207022 386854
rect 206466 368938 206702 369174
rect 206786 368938 207022 369174
rect 206466 368618 206702 368854
rect 206786 368618 207022 368854
rect 206466 350938 206702 351174
rect 206786 350938 207022 351174
rect 206466 350618 206702 350854
rect 206786 350618 207022 350854
rect 206466 332938 206702 333174
rect 206786 332938 207022 333174
rect 206466 332618 206702 332854
rect 206786 332618 207022 332854
rect 206466 314938 206702 315174
rect 206786 314938 207022 315174
rect 206466 314618 206702 314854
rect 206786 314618 207022 314854
rect 206466 296938 206702 297174
rect 206786 296938 207022 297174
rect 206466 296618 206702 296854
rect 206786 296618 207022 296854
rect 206466 278938 206702 279174
rect 206786 278938 207022 279174
rect 206466 278618 206702 278854
rect 206786 278618 207022 278854
rect 206466 260938 206702 261174
rect 206786 260938 207022 261174
rect 206466 260618 206702 260854
rect 206786 260618 207022 260854
rect 206466 242938 206702 243174
rect 206786 242938 207022 243174
rect 206466 242618 206702 242854
rect 206786 242618 207022 242854
rect 206466 224938 206702 225174
rect 206786 224938 207022 225174
rect 206466 224618 206702 224854
rect 206786 224618 207022 224854
rect 206466 206938 206702 207174
rect 206786 206938 207022 207174
rect 206466 206618 206702 206854
rect 206786 206618 207022 206854
rect 206466 188938 206702 189174
rect 206786 188938 207022 189174
rect 206466 188618 206702 188854
rect 206786 188618 207022 188854
rect 206466 170938 206702 171174
rect 206786 170938 207022 171174
rect 206466 170618 206702 170854
rect 206786 170618 207022 170854
rect 206466 152938 206702 153174
rect 206786 152938 207022 153174
rect 206466 152618 206702 152854
rect 206786 152618 207022 152854
rect 206466 134938 206702 135174
rect 206786 134938 207022 135174
rect 206466 134618 206702 134854
rect 206786 134618 207022 134854
rect 206466 116938 206702 117174
rect 206786 116938 207022 117174
rect 206466 116618 206702 116854
rect 206786 116618 207022 116854
rect 206466 98938 206702 99174
rect 206786 98938 207022 99174
rect 206466 98618 206702 98854
rect 206786 98618 207022 98854
rect 206466 80938 206702 81174
rect 206786 80938 207022 81174
rect 206466 80618 206702 80854
rect 206786 80618 207022 80854
rect 206466 62938 206702 63174
rect 206786 62938 207022 63174
rect 206466 62618 206702 62854
rect 206786 62618 207022 62854
rect 206466 44938 206702 45174
rect 206786 44938 207022 45174
rect 206466 44618 206702 44854
rect 206786 44618 207022 44854
rect 206466 26938 206702 27174
rect 206786 26938 207022 27174
rect 206466 26618 206702 26854
rect 206786 26618 207022 26854
rect 206466 8938 206702 9174
rect 206786 8938 207022 9174
rect 206466 8618 206702 8854
rect 206786 8618 207022 8854
rect 206466 -2052 206702 -1816
rect 206786 -2052 207022 -1816
rect 206466 -2372 206702 -2136
rect 206786 -2372 207022 -2136
rect 210186 462776 210422 463012
rect 210506 462776 210742 463012
rect 210186 462456 210422 462692
rect 210506 462456 210742 462692
rect 210186 444658 210422 444894
rect 210506 444658 210742 444894
rect 210186 444338 210422 444574
rect 210506 444338 210742 444574
rect 210186 426658 210422 426894
rect 210506 426658 210742 426894
rect 210186 426338 210422 426574
rect 210506 426338 210742 426574
rect 210186 408658 210422 408894
rect 210506 408658 210742 408894
rect 210186 408338 210422 408574
rect 210506 408338 210742 408574
rect 210186 390658 210422 390894
rect 210506 390658 210742 390894
rect 210186 390338 210422 390574
rect 210506 390338 210742 390574
rect 210186 372658 210422 372894
rect 210506 372658 210742 372894
rect 210186 372338 210422 372574
rect 210506 372338 210742 372574
rect 210186 354658 210422 354894
rect 210506 354658 210742 354894
rect 210186 354338 210422 354574
rect 210506 354338 210742 354574
rect 210186 336658 210422 336894
rect 210506 336658 210742 336894
rect 210186 336338 210422 336574
rect 210506 336338 210742 336574
rect 210186 318658 210422 318894
rect 210506 318658 210742 318894
rect 210186 318338 210422 318574
rect 210506 318338 210742 318574
rect 210186 300658 210422 300894
rect 210506 300658 210742 300894
rect 210186 300338 210422 300574
rect 210506 300338 210742 300574
rect 210186 282658 210422 282894
rect 210506 282658 210742 282894
rect 210186 282338 210422 282574
rect 210506 282338 210742 282574
rect 210186 264658 210422 264894
rect 210506 264658 210742 264894
rect 210186 264338 210422 264574
rect 210506 264338 210742 264574
rect 210186 246658 210422 246894
rect 210506 246658 210742 246894
rect 210186 246338 210422 246574
rect 210506 246338 210742 246574
rect 210186 228658 210422 228894
rect 210506 228658 210742 228894
rect 210186 228338 210422 228574
rect 210506 228338 210742 228574
rect 210186 210658 210422 210894
rect 210506 210658 210742 210894
rect 210186 210338 210422 210574
rect 210506 210338 210742 210574
rect 210186 192658 210422 192894
rect 210506 192658 210742 192894
rect 210186 192338 210422 192574
rect 210506 192338 210742 192574
rect 210186 174658 210422 174894
rect 210506 174658 210742 174894
rect 210186 174338 210422 174574
rect 210506 174338 210742 174574
rect 210186 156658 210422 156894
rect 210506 156658 210742 156894
rect 210186 156338 210422 156574
rect 210506 156338 210742 156574
rect 210186 138658 210422 138894
rect 210506 138658 210742 138894
rect 210186 138338 210422 138574
rect 210506 138338 210742 138574
rect 210186 120658 210422 120894
rect 210506 120658 210742 120894
rect 210186 120338 210422 120574
rect 210506 120338 210742 120574
rect 210186 102658 210422 102894
rect 210506 102658 210742 102894
rect 210186 102338 210422 102574
rect 210506 102338 210742 102574
rect 210186 84658 210422 84894
rect 210506 84658 210742 84894
rect 210186 84338 210422 84574
rect 210506 84338 210742 84574
rect 210186 66658 210422 66894
rect 210506 66658 210742 66894
rect 210186 66338 210422 66574
rect 210506 66338 210742 66574
rect 210186 48658 210422 48894
rect 210506 48658 210742 48894
rect 210186 48338 210422 48574
rect 210506 48338 210742 48574
rect 210186 30658 210422 30894
rect 210506 30658 210742 30894
rect 210186 30338 210422 30574
rect 210506 30338 210742 30574
rect 210186 12658 210422 12894
rect 210506 12658 210742 12894
rect 210186 12338 210422 12574
rect 210506 12338 210742 12574
rect 210186 -3012 210422 -2776
rect 210506 -3012 210742 -2776
rect 210186 -3332 210422 -3096
rect 210506 -3332 210742 -3096
rect 213906 463736 214142 463972
rect 214226 463736 214462 463972
rect 213906 463416 214142 463652
rect 214226 463416 214462 463652
rect 213906 448378 214142 448614
rect 214226 448378 214462 448614
rect 213906 448058 214142 448294
rect 214226 448058 214462 448294
rect 213906 430378 214142 430614
rect 214226 430378 214462 430614
rect 213906 430058 214142 430294
rect 214226 430058 214462 430294
rect 213906 412378 214142 412614
rect 214226 412378 214462 412614
rect 213906 412058 214142 412294
rect 214226 412058 214462 412294
rect 213906 394378 214142 394614
rect 214226 394378 214462 394614
rect 213906 394058 214142 394294
rect 214226 394058 214462 394294
rect 213906 376378 214142 376614
rect 214226 376378 214462 376614
rect 213906 376058 214142 376294
rect 214226 376058 214462 376294
rect 213906 358378 214142 358614
rect 214226 358378 214462 358614
rect 213906 358058 214142 358294
rect 214226 358058 214462 358294
rect 213906 340378 214142 340614
rect 214226 340378 214462 340614
rect 213906 340058 214142 340294
rect 214226 340058 214462 340294
rect 213906 322378 214142 322614
rect 214226 322378 214462 322614
rect 213906 322058 214142 322294
rect 214226 322058 214462 322294
rect 213906 304378 214142 304614
rect 214226 304378 214462 304614
rect 213906 304058 214142 304294
rect 214226 304058 214462 304294
rect 213906 286378 214142 286614
rect 214226 286378 214462 286614
rect 213906 286058 214142 286294
rect 214226 286058 214462 286294
rect 213906 268378 214142 268614
rect 214226 268378 214462 268614
rect 213906 268058 214142 268294
rect 214226 268058 214462 268294
rect 213906 250378 214142 250614
rect 214226 250378 214462 250614
rect 213906 250058 214142 250294
rect 214226 250058 214462 250294
rect 213906 232378 214142 232614
rect 214226 232378 214462 232614
rect 213906 232058 214142 232294
rect 214226 232058 214462 232294
rect 213906 214378 214142 214614
rect 214226 214378 214462 214614
rect 213906 214058 214142 214294
rect 214226 214058 214462 214294
rect 213906 196378 214142 196614
rect 214226 196378 214462 196614
rect 213906 196058 214142 196294
rect 214226 196058 214462 196294
rect 213906 178378 214142 178614
rect 214226 178378 214462 178614
rect 213906 178058 214142 178294
rect 214226 178058 214462 178294
rect 213906 160378 214142 160614
rect 214226 160378 214462 160614
rect 213906 160058 214142 160294
rect 214226 160058 214462 160294
rect 213906 142378 214142 142614
rect 214226 142378 214462 142614
rect 213906 142058 214142 142294
rect 214226 142058 214462 142294
rect 213906 124378 214142 124614
rect 214226 124378 214462 124614
rect 213906 124058 214142 124294
rect 214226 124058 214462 124294
rect 213906 106378 214142 106614
rect 214226 106378 214462 106614
rect 213906 106058 214142 106294
rect 214226 106058 214462 106294
rect 213906 88378 214142 88614
rect 214226 88378 214462 88614
rect 213906 88058 214142 88294
rect 214226 88058 214462 88294
rect 213906 70378 214142 70614
rect 214226 70378 214462 70614
rect 213906 70058 214142 70294
rect 214226 70058 214462 70294
rect 213906 52378 214142 52614
rect 214226 52378 214462 52614
rect 213906 52058 214142 52294
rect 214226 52058 214462 52294
rect 213906 34378 214142 34614
rect 214226 34378 214462 34614
rect 213906 34058 214142 34294
rect 214226 34058 214462 34294
rect 213906 16378 214142 16614
rect 214226 16378 214462 16614
rect 213906 16058 214142 16294
rect 214226 16058 214462 16294
rect 213906 -3972 214142 -3736
rect 214226 -3972 214462 -3736
rect 213906 -4292 214142 -4056
rect 214226 -4292 214462 -4056
rect 220746 460856 220982 461092
rect 221066 460856 221302 461092
rect 220746 460536 220982 460772
rect 221066 460536 221302 460772
rect 220746 455218 220982 455454
rect 221066 455218 221302 455454
rect 220746 454898 220982 455134
rect 221066 454898 221302 455134
rect 220746 437218 220982 437454
rect 221066 437218 221302 437454
rect 220746 436898 220982 437134
rect 221066 436898 221302 437134
rect 220746 419218 220982 419454
rect 221066 419218 221302 419454
rect 220746 418898 220982 419134
rect 221066 418898 221302 419134
rect 220746 401218 220982 401454
rect 221066 401218 221302 401454
rect 220746 400898 220982 401134
rect 221066 400898 221302 401134
rect 220746 383218 220982 383454
rect 221066 383218 221302 383454
rect 220746 382898 220982 383134
rect 221066 382898 221302 383134
rect 220746 365218 220982 365454
rect 221066 365218 221302 365454
rect 220746 364898 220982 365134
rect 221066 364898 221302 365134
rect 220746 347218 220982 347454
rect 221066 347218 221302 347454
rect 220746 346898 220982 347134
rect 221066 346898 221302 347134
rect 220746 329218 220982 329454
rect 221066 329218 221302 329454
rect 220746 328898 220982 329134
rect 221066 328898 221302 329134
rect 220746 311218 220982 311454
rect 221066 311218 221302 311454
rect 220746 310898 220982 311134
rect 221066 310898 221302 311134
rect 220746 293218 220982 293454
rect 221066 293218 221302 293454
rect 220746 292898 220982 293134
rect 221066 292898 221302 293134
rect 220746 275218 220982 275454
rect 221066 275218 221302 275454
rect 220746 274898 220982 275134
rect 221066 274898 221302 275134
rect 220746 257218 220982 257454
rect 221066 257218 221302 257454
rect 220746 256898 220982 257134
rect 221066 256898 221302 257134
rect 220746 239218 220982 239454
rect 221066 239218 221302 239454
rect 220746 238898 220982 239134
rect 221066 238898 221302 239134
rect 220746 221218 220982 221454
rect 221066 221218 221302 221454
rect 220746 220898 220982 221134
rect 221066 220898 221302 221134
rect 220746 203218 220982 203454
rect 221066 203218 221302 203454
rect 220746 202898 220982 203134
rect 221066 202898 221302 203134
rect 220746 185218 220982 185454
rect 221066 185218 221302 185454
rect 220746 184898 220982 185134
rect 221066 184898 221302 185134
rect 220746 167218 220982 167454
rect 221066 167218 221302 167454
rect 220746 166898 220982 167134
rect 221066 166898 221302 167134
rect 220746 149218 220982 149454
rect 221066 149218 221302 149454
rect 220746 148898 220982 149134
rect 221066 148898 221302 149134
rect 220746 131218 220982 131454
rect 221066 131218 221302 131454
rect 220746 130898 220982 131134
rect 221066 130898 221302 131134
rect 220746 113218 220982 113454
rect 221066 113218 221302 113454
rect 220746 112898 220982 113134
rect 221066 112898 221302 113134
rect 220746 95218 220982 95454
rect 221066 95218 221302 95454
rect 220746 94898 220982 95134
rect 221066 94898 221302 95134
rect 220746 77218 220982 77454
rect 221066 77218 221302 77454
rect 220746 76898 220982 77134
rect 221066 76898 221302 77134
rect 220746 59218 220982 59454
rect 221066 59218 221302 59454
rect 220746 58898 220982 59134
rect 221066 58898 221302 59134
rect 220746 41218 220982 41454
rect 221066 41218 221302 41454
rect 220746 40898 220982 41134
rect 221066 40898 221302 41134
rect 220746 23218 220982 23454
rect 221066 23218 221302 23454
rect 220746 22898 220982 23134
rect 221066 22898 221302 23134
rect 220746 5218 220982 5454
rect 221066 5218 221302 5454
rect 220746 4898 220982 5134
rect 221066 4898 221302 5134
rect 220746 -1092 220982 -856
rect 221066 -1092 221302 -856
rect 220746 -1412 220982 -1176
rect 221066 -1412 221302 -1176
rect 224466 461816 224702 462052
rect 224786 461816 225022 462052
rect 224466 461496 224702 461732
rect 224786 461496 225022 461732
rect 224466 440938 224702 441174
rect 224786 440938 225022 441174
rect 224466 440618 224702 440854
rect 224786 440618 225022 440854
rect 224466 422938 224702 423174
rect 224786 422938 225022 423174
rect 224466 422618 224702 422854
rect 224786 422618 225022 422854
rect 224466 404938 224702 405174
rect 224786 404938 225022 405174
rect 224466 404618 224702 404854
rect 224786 404618 225022 404854
rect 224466 386938 224702 387174
rect 224786 386938 225022 387174
rect 224466 386618 224702 386854
rect 224786 386618 225022 386854
rect 224466 368938 224702 369174
rect 224786 368938 225022 369174
rect 224466 368618 224702 368854
rect 224786 368618 225022 368854
rect 224466 350938 224702 351174
rect 224786 350938 225022 351174
rect 224466 350618 224702 350854
rect 224786 350618 225022 350854
rect 224466 332938 224702 333174
rect 224786 332938 225022 333174
rect 224466 332618 224702 332854
rect 224786 332618 225022 332854
rect 224466 314938 224702 315174
rect 224786 314938 225022 315174
rect 224466 314618 224702 314854
rect 224786 314618 225022 314854
rect 224466 296938 224702 297174
rect 224786 296938 225022 297174
rect 224466 296618 224702 296854
rect 224786 296618 225022 296854
rect 224466 278938 224702 279174
rect 224786 278938 225022 279174
rect 224466 278618 224702 278854
rect 224786 278618 225022 278854
rect 224466 260938 224702 261174
rect 224786 260938 225022 261174
rect 224466 260618 224702 260854
rect 224786 260618 225022 260854
rect 224466 242938 224702 243174
rect 224786 242938 225022 243174
rect 224466 242618 224702 242854
rect 224786 242618 225022 242854
rect 224466 224938 224702 225174
rect 224786 224938 225022 225174
rect 224466 224618 224702 224854
rect 224786 224618 225022 224854
rect 224466 206938 224702 207174
rect 224786 206938 225022 207174
rect 224466 206618 224702 206854
rect 224786 206618 225022 206854
rect 224466 188938 224702 189174
rect 224786 188938 225022 189174
rect 224466 188618 224702 188854
rect 224786 188618 225022 188854
rect 224466 170938 224702 171174
rect 224786 170938 225022 171174
rect 224466 170618 224702 170854
rect 224786 170618 225022 170854
rect 224466 152938 224702 153174
rect 224786 152938 225022 153174
rect 224466 152618 224702 152854
rect 224786 152618 225022 152854
rect 224466 134938 224702 135174
rect 224786 134938 225022 135174
rect 224466 134618 224702 134854
rect 224786 134618 225022 134854
rect 224466 116938 224702 117174
rect 224786 116938 225022 117174
rect 224466 116618 224702 116854
rect 224786 116618 225022 116854
rect 224466 98938 224702 99174
rect 224786 98938 225022 99174
rect 224466 98618 224702 98854
rect 224786 98618 225022 98854
rect 224466 80938 224702 81174
rect 224786 80938 225022 81174
rect 224466 80618 224702 80854
rect 224786 80618 225022 80854
rect 224466 62938 224702 63174
rect 224786 62938 225022 63174
rect 224466 62618 224702 62854
rect 224786 62618 225022 62854
rect 224466 44938 224702 45174
rect 224786 44938 225022 45174
rect 224466 44618 224702 44854
rect 224786 44618 225022 44854
rect 224466 26938 224702 27174
rect 224786 26938 225022 27174
rect 224466 26618 224702 26854
rect 224786 26618 225022 26854
rect 224466 8938 224702 9174
rect 224786 8938 225022 9174
rect 224466 8618 224702 8854
rect 224786 8618 225022 8854
rect 224466 -2052 224702 -1816
rect 224786 -2052 225022 -1816
rect 224466 -2372 224702 -2136
rect 224786 -2372 225022 -2136
rect 228186 462776 228422 463012
rect 228506 462776 228742 463012
rect 228186 462456 228422 462692
rect 228506 462456 228742 462692
rect 228186 444658 228422 444894
rect 228506 444658 228742 444894
rect 228186 444338 228422 444574
rect 228506 444338 228742 444574
rect 228186 426658 228422 426894
rect 228506 426658 228742 426894
rect 228186 426338 228422 426574
rect 228506 426338 228742 426574
rect 228186 408658 228422 408894
rect 228506 408658 228742 408894
rect 228186 408338 228422 408574
rect 228506 408338 228742 408574
rect 228186 390658 228422 390894
rect 228506 390658 228742 390894
rect 228186 390338 228422 390574
rect 228506 390338 228742 390574
rect 228186 372658 228422 372894
rect 228506 372658 228742 372894
rect 228186 372338 228422 372574
rect 228506 372338 228742 372574
rect 228186 354658 228422 354894
rect 228506 354658 228742 354894
rect 228186 354338 228422 354574
rect 228506 354338 228742 354574
rect 228186 336658 228422 336894
rect 228506 336658 228742 336894
rect 228186 336338 228422 336574
rect 228506 336338 228742 336574
rect 228186 318658 228422 318894
rect 228506 318658 228742 318894
rect 228186 318338 228422 318574
rect 228506 318338 228742 318574
rect 228186 300658 228422 300894
rect 228506 300658 228742 300894
rect 228186 300338 228422 300574
rect 228506 300338 228742 300574
rect 228186 282658 228422 282894
rect 228506 282658 228742 282894
rect 228186 282338 228422 282574
rect 228506 282338 228742 282574
rect 228186 264658 228422 264894
rect 228506 264658 228742 264894
rect 228186 264338 228422 264574
rect 228506 264338 228742 264574
rect 228186 246658 228422 246894
rect 228506 246658 228742 246894
rect 228186 246338 228422 246574
rect 228506 246338 228742 246574
rect 228186 228658 228422 228894
rect 228506 228658 228742 228894
rect 228186 228338 228422 228574
rect 228506 228338 228742 228574
rect 228186 210658 228422 210894
rect 228506 210658 228742 210894
rect 228186 210338 228422 210574
rect 228506 210338 228742 210574
rect 228186 192658 228422 192894
rect 228506 192658 228742 192894
rect 228186 192338 228422 192574
rect 228506 192338 228742 192574
rect 228186 174658 228422 174894
rect 228506 174658 228742 174894
rect 228186 174338 228422 174574
rect 228506 174338 228742 174574
rect 228186 156658 228422 156894
rect 228506 156658 228742 156894
rect 228186 156338 228422 156574
rect 228506 156338 228742 156574
rect 228186 138658 228422 138894
rect 228506 138658 228742 138894
rect 228186 138338 228422 138574
rect 228506 138338 228742 138574
rect 228186 120658 228422 120894
rect 228506 120658 228742 120894
rect 228186 120338 228422 120574
rect 228506 120338 228742 120574
rect 228186 102658 228422 102894
rect 228506 102658 228742 102894
rect 228186 102338 228422 102574
rect 228506 102338 228742 102574
rect 228186 84658 228422 84894
rect 228506 84658 228742 84894
rect 228186 84338 228422 84574
rect 228506 84338 228742 84574
rect 228186 66658 228422 66894
rect 228506 66658 228742 66894
rect 228186 66338 228422 66574
rect 228506 66338 228742 66574
rect 228186 48658 228422 48894
rect 228506 48658 228742 48894
rect 228186 48338 228422 48574
rect 228506 48338 228742 48574
rect 228186 30658 228422 30894
rect 228506 30658 228742 30894
rect 228186 30338 228422 30574
rect 228506 30338 228742 30574
rect 228186 12658 228422 12894
rect 228506 12658 228742 12894
rect 228186 12338 228422 12574
rect 228506 12338 228742 12574
rect 228186 -3012 228422 -2776
rect 228506 -3012 228742 -2776
rect 228186 -3332 228422 -3096
rect 228506 -3332 228742 -3096
rect 231906 463736 232142 463972
rect 232226 463736 232462 463972
rect 231906 463416 232142 463652
rect 232226 463416 232462 463652
rect 231906 448378 232142 448614
rect 232226 448378 232462 448614
rect 231906 448058 232142 448294
rect 232226 448058 232462 448294
rect 231906 430378 232142 430614
rect 232226 430378 232462 430614
rect 231906 430058 232142 430294
rect 232226 430058 232462 430294
rect 231906 412378 232142 412614
rect 232226 412378 232462 412614
rect 231906 412058 232142 412294
rect 232226 412058 232462 412294
rect 231906 394378 232142 394614
rect 232226 394378 232462 394614
rect 231906 394058 232142 394294
rect 232226 394058 232462 394294
rect 231906 376378 232142 376614
rect 232226 376378 232462 376614
rect 231906 376058 232142 376294
rect 232226 376058 232462 376294
rect 231906 358378 232142 358614
rect 232226 358378 232462 358614
rect 231906 358058 232142 358294
rect 232226 358058 232462 358294
rect 231906 340378 232142 340614
rect 232226 340378 232462 340614
rect 231906 340058 232142 340294
rect 232226 340058 232462 340294
rect 231906 322378 232142 322614
rect 232226 322378 232462 322614
rect 231906 322058 232142 322294
rect 232226 322058 232462 322294
rect 231906 304378 232142 304614
rect 232226 304378 232462 304614
rect 231906 304058 232142 304294
rect 232226 304058 232462 304294
rect 231906 286378 232142 286614
rect 232226 286378 232462 286614
rect 231906 286058 232142 286294
rect 232226 286058 232462 286294
rect 231906 268378 232142 268614
rect 232226 268378 232462 268614
rect 231906 268058 232142 268294
rect 232226 268058 232462 268294
rect 231906 250378 232142 250614
rect 232226 250378 232462 250614
rect 231906 250058 232142 250294
rect 232226 250058 232462 250294
rect 231906 232378 232142 232614
rect 232226 232378 232462 232614
rect 231906 232058 232142 232294
rect 232226 232058 232462 232294
rect 231906 214378 232142 214614
rect 232226 214378 232462 214614
rect 231906 214058 232142 214294
rect 232226 214058 232462 214294
rect 231906 196378 232142 196614
rect 232226 196378 232462 196614
rect 231906 196058 232142 196294
rect 232226 196058 232462 196294
rect 231906 178378 232142 178614
rect 232226 178378 232462 178614
rect 231906 178058 232142 178294
rect 232226 178058 232462 178294
rect 231906 160378 232142 160614
rect 232226 160378 232462 160614
rect 231906 160058 232142 160294
rect 232226 160058 232462 160294
rect 231906 142378 232142 142614
rect 232226 142378 232462 142614
rect 231906 142058 232142 142294
rect 232226 142058 232462 142294
rect 231906 124378 232142 124614
rect 232226 124378 232462 124614
rect 231906 124058 232142 124294
rect 232226 124058 232462 124294
rect 231906 106378 232142 106614
rect 232226 106378 232462 106614
rect 231906 106058 232142 106294
rect 232226 106058 232462 106294
rect 231906 88378 232142 88614
rect 232226 88378 232462 88614
rect 231906 88058 232142 88294
rect 232226 88058 232462 88294
rect 231906 70378 232142 70614
rect 232226 70378 232462 70614
rect 231906 70058 232142 70294
rect 232226 70058 232462 70294
rect 231906 52378 232142 52614
rect 232226 52378 232462 52614
rect 231906 52058 232142 52294
rect 232226 52058 232462 52294
rect 231906 34378 232142 34614
rect 232226 34378 232462 34614
rect 231906 34058 232142 34294
rect 232226 34058 232462 34294
rect 231906 16378 232142 16614
rect 232226 16378 232462 16614
rect 231906 16058 232142 16294
rect 232226 16058 232462 16294
rect 231906 -3972 232142 -3736
rect 232226 -3972 232462 -3736
rect 231906 -4292 232142 -4056
rect 232226 -4292 232462 -4056
rect 238746 460856 238982 461092
rect 239066 460856 239302 461092
rect 238746 460536 238982 460772
rect 239066 460536 239302 460772
rect 238746 455218 238982 455454
rect 239066 455218 239302 455454
rect 238746 454898 238982 455134
rect 239066 454898 239302 455134
rect 238746 437218 238982 437454
rect 239066 437218 239302 437454
rect 238746 436898 238982 437134
rect 239066 436898 239302 437134
rect 238746 419218 238982 419454
rect 239066 419218 239302 419454
rect 238746 418898 238982 419134
rect 239066 418898 239302 419134
rect 238746 401218 238982 401454
rect 239066 401218 239302 401454
rect 238746 400898 238982 401134
rect 239066 400898 239302 401134
rect 238746 383218 238982 383454
rect 239066 383218 239302 383454
rect 238746 382898 238982 383134
rect 239066 382898 239302 383134
rect 238746 365218 238982 365454
rect 239066 365218 239302 365454
rect 238746 364898 238982 365134
rect 239066 364898 239302 365134
rect 238746 347218 238982 347454
rect 239066 347218 239302 347454
rect 238746 346898 238982 347134
rect 239066 346898 239302 347134
rect 238746 329218 238982 329454
rect 239066 329218 239302 329454
rect 238746 328898 238982 329134
rect 239066 328898 239302 329134
rect 238746 311218 238982 311454
rect 239066 311218 239302 311454
rect 238746 310898 238982 311134
rect 239066 310898 239302 311134
rect 238746 293218 238982 293454
rect 239066 293218 239302 293454
rect 238746 292898 238982 293134
rect 239066 292898 239302 293134
rect 238746 275218 238982 275454
rect 239066 275218 239302 275454
rect 238746 274898 238982 275134
rect 239066 274898 239302 275134
rect 238746 257218 238982 257454
rect 239066 257218 239302 257454
rect 238746 256898 238982 257134
rect 239066 256898 239302 257134
rect 238746 239218 238982 239454
rect 239066 239218 239302 239454
rect 238746 238898 238982 239134
rect 239066 238898 239302 239134
rect 238746 221218 238982 221454
rect 239066 221218 239302 221454
rect 238746 220898 238982 221134
rect 239066 220898 239302 221134
rect 238746 203218 238982 203454
rect 239066 203218 239302 203454
rect 238746 202898 238982 203134
rect 239066 202898 239302 203134
rect 238746 185218 238982 185454
rect 239066 185218 239302 185454
rect 238746 184898 238982 185134
rect 239066 184898 239302 185134
rect 238746 167218 238982 167454
rect 239066 167218 239302 167454
rect 238746 166898 238982 167134
rect 239066 166898 239302 167134
rect 238746 149218 238982 149454
rect 239066 149218 239302 149454
rect 238746 148898 238982 149134
rect 239066 148898 239302 149134
rect 238746 131218 238982 131454
rect 239066 131218 239302 131454
rect 238746 130898 238982 131134
rect 239066 130898 239302 131134
rect 238746 113218 238982 113454
rect 239066 113218 239302 113454
rect 238746 112898 238982 113134
rect 239066 112898 239302 113134
rect 238746 95218 238982 95454
rect 239066 95218 239302 95454
rect 238746 94898 238982 95134
rect 239066 94898 239302 95134
rect 238746 77218 238982 77454
rect 239066 77218 239302 77454
rect 238746 76898 238982 77134
rect 239066 76898 239302 77134
rect 238746 59218 238982 59454
rect 239066 59218 239302 59454
rect 238746 58898 238982 59134
rect 239066 58898 239302 59134
rect 238746 41218 238982 41454
rect 239066 41218 239302 41454
rect 238746 40898 238982 41134
rect 239066 40898 239302 41134
rect 238746 23218 238982 23454
rect 239066 23218 239302 23454
rect 238746 22898 238982 23134
rect 239066 22898 239302 23134
rect 238746 5218 238982 5454
rect 239066 5218 239302 5454
rect 238746 4898 238982 5134
rect 239066 4898 239302 5134
rect 238746 -1092 238982 -856
rect 239066 -1092 239302 -856
rect 238746 -1412 238982 -1176
rect 239066 -1412 239302 -1176
rect 242466 461816 242702 462052
rect 242786 461816 243022 462052
rect 242466 461496 242702 461732
rect 242786 461496 243022 461732
rect 242466 440938 242702 441174
rect 242786 440938 243022 441174
rect 242466 440618 242702 440854
rect 242786 440618 243022 440854
rect 242466 422938 242702 423174
rect 242786 422938 243022 423174
rect 242466 422618 242702 422854
rect 242786 422618 243022 422854
rect 242466 404938 242702 405174
rect 242786 404938 243022 405174
rect 242466 404618 242702 404854
rect 242786 404618 243022 404854
rect 242466 386938 242702 387174
rect 242786 386938 243022 387174
rect 242466 386618 242702 386854
rect 242786 386618 243022 386854
rect 242466 368938 242702 369174
rect 242786 368938 243022 369174
rect 242466 368618 242702 368854
rect 242786 368618 243022 368854
rect 242466 350938 242702 351174
rect 242786 350938 243022 351174
rect 242466 350618 242702 350854
rect 242786 350618 243022 350854
rect 242466 332938 242702 333174
rect 242786 332938 243022 333174
rect 242466 332618 242702 332854
rect 242786 332618 243022 332854
rect 242466 314938 242702 315174
rect 242786 314938 243022 315174
rect 242466 314618 242702 314854
rect 242786 314618 243022 314854
rect 242466 296938 242702 297174
rect 242786 296938 243022 297174
rect 242466 296618 242702 296854
rect 242786 296618 243022 296854
rect 242466 278938 242702 279174
rect 242786 278938 243022 279174
rect 242466 278618 242702 278854
rect 242786 278618 243022 278854
rect 242466 260938 242702 261174
rect 242786 260938 243022 261174
rect 242466 260618 242702 260854
rect 242786 260618 243022 260854
rect 242466 242938 242702 243174
rect 242786 242938 243022 243174
rect 242466 242618 242702 242854
rect 242786 242618 243022 242854
rect 242466 224938 242702 225174
rect 242786 224938 243022 225174
rect 242466 224618 242702 224854
rect 242786 224618 243022 224854
rect 242466 206938 242702 207174
rect 242786 206938 243022 207174
rect 242466 206618 242702 206854
rect 242786 206618 243022 206854
rect 242466 188938 242702 189174
rect 242786 188938 243022 189174
rect 242466 188618 242702 188854
rect 242786 188618 243022 188854
rect 242466 170938 242702 171174
rect 242786 170938 243022 171174
rect 242466 170618 242702 170854
rect 242786 170618 243022 170854
rect 242466 152938 242702 153174
rect 242786 152938 243022 153174
rect 242466 152618 242702 152854
rect 242786 152618 243022 152854
rect 242466 134938 242702 135174
rect 242786 134938 243022 135174
rect 242466 134618 242702 134854
rect 242786 134618 243022 134854
rect 242466 116938 242702 117174
rect 242786 116938 243022 117174
rect 242466 116618 242702 116854
rect 242786 116618 243022 116854
rect 242466 98938 242702 99174
rect 242786 98938 243022 99174
rect 242466 98618 242702 98854
rect 242786 98618 243022 98854
rect 242466 80938 242702 81174
rect 242786 80938 243022 81174
rect 242466 80618 242702 80854
rect 242786 80618 243022 80854
rect 242466 62938 242702 63174
rect 242786 62938 243022 63174
rect 242466 62618 242702 62854
rect 242786 62618 243022 62854
rect 242466 44938 242702 45174
rect 242786 44938 243022 45174
rect 242466 44618 242702 44854
rect 242786 44618 243022 44854
rect 242466 26938 242702 27174
rect 242786 26938 243022 27174
rect 242466 26618 242702 26854
rect 242786 26618 243022 26854
rect 242466 8938 242702 9174
rect 242786 8938 243022 9174
rect 242466 8618 242702 8854
rect 242786 8618 243022 8854
rect 242466 -2052 242702 -1816
rect 242786 -2052 243022 -1816
rect 242466 -2372 242702 -2136
rect 242786 -2372 243022 -2136
rect 246186 462776 246422 463012
rect 246506 462776 246742 463012
rect 246186 462456 246422 462692
rect 246506 462456 246742 462692
rect 246186 444658 246422 444894
rect 246506 444658 246742 444894
rect 246186 444338 246422 444574
rect 246506 444338 246742 444574
rect 246186 426658 246422 426894
rect 246506 426658 246742 426894
rect 246186 426338 246422 426574
rect 246506 426338 246742 426574
rect 246186 408658 246422 408894
rect 246506 408658 246742 408894
rect 246186 408338 246422 408574
rect 246506 408338 246742 408574
rect 246186 390658 246422 390894
rect 246506 390658 246742 390894
rect 246186 390338 246422 390574
rect 246506 390338 246742 390574
rect 246186 372658 246422 372894
rect 246506 372658 246742 372894
rect 246186 372338 246422 372574
rect 246506 372338 246742 372574
rect 246186 354658 246422 354894
rect 246506 354658 246742 354894
rect 246186 354338 246422 354574
rect 246506 354338 246742 354574
rect 246186 336658 246422 336894
rect 246506 336658 246742 336894
rect 246186 336338 246422 336574
rect 246506 336338 246742 336574
rect 246186 318658 246422 318894
rect 246506 318658 246742 318894
rect 246186 318338 246422 318574
rect 246506 318338 246742 318574
rect 246186 300658 246422 300894
rect 246506 300658 246742 300894
rect 246186 300338 246422 300574
rect 246506 300338 246742 300574
rect 246186 282658 246422 282894
rect 246506 282658 246742 282894
rect 246186 282338 246422 282574
rect 246506 282338 246742 282574
rect 246186 264658 246422 264894
rect 246506 264658 246742 264894
rect 246186 264338 246422 264574
rect 246506 264338 246742 264574
rect 246186 246658 246422 246894
rect 246506 246658 246742 246894
rect 246186 246338 246422 246574
rect 246506 246338 246742 246574
rect 246186 228658 246422 228894
rect 246506 228658 246742 228894
rect 246186 228338 246422 228574
rect 246506 228338 246742 228574
rect 246186 210658 246422 210894
rect 246506 210658 246742 210894
rect 246186 210338 246422 210574
rect 246506 210338 246742 210574
rect 246186 192658 246422 192894
rect 246506 192658 246742 192894
rect 246186 192338 246422 192574
rect 246506 192338 246742 192574
rect 246186 174658 246422 174894
rect 246506 174658 246742 174894
rect 246186 174338 246422 174574
rect 246506 174338 246742 174574
rect 246186 156658 246422 156894
rect 246506 156658 246742 156894
rect 246186 156338 246422 156574
rect 246506 156338 246742 156574
rect 246186 138658 246422 138894
rect 246506 138658 246742 138894
rect 246186 138338 246422 138574
rect 246506 138338 246742 138574
rect 246186 120658 246422 120894
rect 246506 120658 246742 120894
rect 246186 120338 246422 120574
rect 246506 120338 246742 120574
rect 246186 102658 246422 102894
rect 246506 102658 246742 102894
rect 246186 102338 246422 102574
rect 246506 102338 246742 102574
rect 246186 84658 246422 84894
rect 246506 84658 246742 84894
rect 246186 84338 246422 84574
rect 246506 84338 246742 84574
rect 246186 66658 246422 66894
rect 246506 66658 246742 66894
rect 246186 66338 246422 66574
rect 246506 66338 246742 66574
rect 246186 48658 246422 48894
rect 246506 48658 246742 48894
rect 246186 48338 246422 48574
rect 246506 48338 246742 48574
rect 246186 30658 246422 30894
rect 246506 30658 246742 30894
rect 246186 30338 246422 30574
rect 246506 30338 246742 30574
rect 246186 12658 246422 12894
rect 246506 12658 246742 12894
rect 246186 12338 246422 12574
rect 246506 12338 246742 12574
rect 246186 -3012 246422 -2776
rect 246506 -3012 246742 -2776
rect 246186 -3332 246422 -3096
rect 246506 -3332 246742 -3096
rect 249906 463736 250142 463972
rect 250226 463736 250462 463972
rect 249906 463416 250142 463652
rect 250226 463416 250462 463652
rect 249906 448378 250142 448614
rect 250226 448378 250462 448614
rect 249906 448058 250142 448294
rect 250226 448058 250462 448294
rect 249906 430378 250142 430614
rect 250226 430378 250462 430614
rect 249906 430058 250142 430294
rect 250226 430058 250462 430294
rect 249906 412378 250142 412614
rect 250226 412378 250462 412614
rect 249906 412058 250142 412294
rect 250226 412058 250462 412294
rect 249906 394378 250142 394614
rect 250226 394378 250462 394614
rect 249906 394058 250142 394294
rect 250226 394058 250462 394294
rect 249906 376378 250142 376614
rect 250226 376378 250462 376614
rect 249906 376058 250142 376294
rect 250226 376058 250462 376294
rect 249906 358378 250142 358614
rect 250226 358378 250462 358614
rect 249906 358058 250142 358294
rect 250226 358058 250462 358294
rect 249906 340378 250142 340614
rect 250226 340378 250462 340614
rect 249906 340058 250142 340294
rect 250226 340058 250462 340294
rect 249906 322378 250142 322614
rect 250226 322378 250462 322614
rect 249906 322058 250142 322294
rect 250226 322058 250462 322294
rect 249906 304378 250142 304614
rect 250226 304378 250462 304614
rect 249906 304058 250142 304294
rect 250226 304058 250462 304294
rect 249906 286378 250142 286614
rect 250226 286378 250462 286614
rect 249906 286058 250142 286294
rect 250226 286058 250462 286294
rect 249906 268378 250142 268614
rect 250226 268378 250462 268614
rect 249906 268058 250142 268294
rect 250226 268058 250462 268294
rect 249906 250378 250142 250614
rect 250226 250378 250462 250614
rect 249906 250058 250142 250294
rect 250226 250058 250462 250294
rect 249906 232378 250142 232614
rect 250226 232378 250462 232614
rect 249906 232058 250142 232294
rect 250226 232058 250462 232294
rect 249906 214378 250142 214614
rect 250226 214378 250462 214614
rect 249906 214058 250142 214294
rect 250226 214058 250462 214294
rect 249906 196378 250142 196614
rect 250226 196378 250462 196614
rect 249906 196058 250142 196294
rect 250226 196058 250462 196294
rect 249906 178378 250142 178614
rect 250226 178378 250462 178614
rect 249906 178058 250142 178294
rect 250226 178058 250462 178294
rect 249906 160378 250142 160614
rect 250226 160378 250462 160614
rect 249906 160058 250142 160294
rect 250226 160058 250462 160294
rect 249906 142378 250142 142614
rect 250226 142378 250462 142614
rect 249906 142058 250142 142294
rect 250226 142058 250462 142294
rect 249906 124378 250142 124614
rect 250226 124378 250462 124614
rect 249906 124058 250142 124294
rect 250226 124058 250462 124294
rect 249906 106378 250142 106614
rect 250226 106378 250462 106614
rect 249906 106058 250142 106294
rect 250226 106058 250462 106294
rect 249906 88378 250142 88614
rect 250226 88378 250462 88614
rect 249906 88058 250142 88294
rect 250226 88058 250462 88294
rect 249906 70378 250142 70614
rect 250226 70378 250462 70614
rect 249906 70058 250142 70294
rect 250226 70058 250462 70294
rect 249906 52378 250142 52614
rect 250226 52378 250462 52614
rect 249906 52058 250142 52294
rect 250226 52058 250462 52294
rect 249906 34378 250142 34614
rect 250226 34378 250462 34614
rect 249906 34058 250142 34294
rect 250226 34058 250462 34294
rect 249906 16378 250142 16614
rect 250226 16378 250462 16614
rect 249906 16058 250142 16294
rect 250226 16058 250462 16294
rect 249906 -3972 250142 -3736
rect 250226 -3972 250462 -3736
rect 249906 -4292 250142 -4056
rect 250226 -4292 250462 -4056
rect 256746 460856 256982 461092
rect 257066 460856 257302 461092
rect 256746 460536 256982 460772
rect 257066 460536 257302 460772
rect 256746 455218 256982 455454
rect 257066 455218 257302 455454
rect 256746 454898 256982 455134
rect 257066 454898 257302 455134
rect 256746 437218 256982 437454
rect 257066 437218 257302 437454
rect 256746 436898 256982 437134
rect 257066 436898 257302 437134
rect 256746 419218 256982 419454
rect 257066 419218 257302 419454
rect 256746 418898 256982 419134
rect 257066 418898 257302 419134
rect 256746 401218 256982 401454
rect 257066 401218 257302 401454
rect 256746 400898 256982 401134
rect 257066 400898 257302 401134
rect 256746 383218 256982 383454
rect 257066 383218 257302 383454
rect 256746 382898 256982 383134
rect 257066 382898 257302 383134
rect 256746 365218 256982 365454
rect 257066 365218 257302 365454
rect 256746 364898 256982 365134
rect 257066 364898 257302 365134
rect 256746 347218 256982 347454
rect 257066 347218 257302 347454
rect 256746 346898 256982 347134
rect 257066 346898 257302 347134
rect 256746 329218 256982 329454
rect 257066 329218 257302 329454
rect 256746 328898 256982 329134
rect 257066 328898 257302 329134
rect 256746 311218 256982 311454
rect 257066 311218 257302 311454
rect 256746 310898 256982 311134
rect 257066 310898 257302 311134
rect 256746 293218 256982 293454
rect 257066 293218 257302 293454
rect 256746 292898 256982 293134
rect 257066 292898 257302 293134
rect 256746 275218 256982 275454
rect 257066 275218 257302 275454
rect 256746 274898 256982 275134
rect 257066 274898 257302 275134
rect 256746 257218 256982 257454
rect 257066 257218 257302 257454
rect 256746 256898 256982 257134
rect 257066 256898 257302 257134
rect 256746 239218 256982 239454
rect 257066 239218 257302 239454
rect 256746 238898 256982 239134
rect 257066 238898 257302 239134
rect 256746 221218 256982 221454
rect 257066 221218 257302 221454
rect 256746 220898 256982 221134
rect 257066 220898 257302 221134
rect 256746 203218 256982 203454
rect 257066 203218 257302 203454
rect 256746 202898 256982 203134
rect 257066 202898 257302 203134
rect 256746 185218 256982 185454
rect 257066 185218 257302 185454
rect 256746 184898 256982 185134
rect 257066 184898 257302 185134
rect 256746 167218 256982 167454
rect 257066 167218 257302 167454
rect 256746 166898 256982 167134
rect 257066 166898 257302 167134
rect 256746 149218 256982 149454
rect 257066 149218 257302 149454
rect 256746 148898 256982 149134
rect 257066 148898 257302 149134
rect 256746 131218 256982 131454
rect 257066 131218 257302 131454
rect 256746 130898 256982 131134
rect 257066 130898 257302 131134
rect 256746 113218 256982 113454
rect 257066 113218 257302 113454
rect 256746 112898 256982 113134
rect 257066 112898 257302 113134
rect 256746 95218 256982 95454
rect 257066 95218 257302 95454
rect 256746 94898 256982 95134
rect 257066 94898 257302 95134
rect 256746 77218 256982 77454
rect 257066 77218 257302 77454
rect 256746 76898 256982 77134
rect 257066 76898 257302 77134
rect 256746 59218 256982 59454
rect 257066 59218 257302 59454
rect 256746 58898 256982 59134
rect 257066 58898 257302 59134
rect 256746 41218 256982 41454
rect 257066 41218 257302 41454
rect 256746 40898 256982 41134
rect 257066 40898 257302 41134
rect 256746 23218 256982 23454
rect 257066 23218 257302 23454
rect 256746 22898 256982 23134
rect 257066 22898 257302 23134
rect 256746 5218 256982 5454
rect 257066 5218 257302 5454
rect 256746 4898 256982 5134
rect 257066 4898 257302 5134
rect 256746 -1092 256982 -856
rect 257066 -1092 257302 -856
rect 256746 -1412 256982 -1176
rect 257066 -1412 257302 -1176
rect 260466 461816 260702 462052
rect 260786 461816 261022 462052
rect 260466 461496 260702 461732
rect 260786 461496 261022 461732
rect 260466 440938 260702 441174
rect 260786 440938 261022 441174
rect 260466 440618 260702 440854
rect 260786 440618 261022 440854
rect 260466 422938 260702 423174
rect 260786 422938 261022 423174
rect 260466 422618 260702 422854
rect 260786 422618 261022 422854
rect 260466 404938 260702 405174
rect 260786 404938 261022 405174
rect 260466 404618 260702 404854
rect 260786 404618 261022 404854
rect 260466 386938 260702 387174
rect 260786 386938 261022 387174
rect 260466 386618 260702 386854
rect 260786 386618 261022 386854
rect 260466 368938 260702 369174
rect 260786 368938 261022 369174
rect 260466 368618 260702 368854
rect 260786 368618 261022 368854
rect 260466 350938 260702 351174
rect 260786 350938 261022 351174
rect 260466 350618 260702 350854
rect 260786 350618 261022 350854
rect 260466 332938 260702 333174
rect 260786 332938 261022 333174
rect 260466 332618 260702 332854
rect 260786 332618 261022 332854
rect 260466 314938 260702 315174
rect 260786 314938 261022 315174
rect 260466 314618 260702 314854
rect 260786 314618 261022 314854
rect 260466 296938 260702 297174
rect 260786 296938 261022 297174
rect 260466 296618 260702 296854
rect 260786 296618 261022 296854
rect 260466 278938 260702 279174
rect 260786 278938 261022 279174
rect 260466 278618 260702 278854
rect 260786 278618 261022 278854
rect 260466 260938 260702 261174
rect 260786 260938 261022 261174
rect 260466 260618 260702 260854
rect 260786 260618 261022 260854
rect 260466 242938 260702 243174
rect 260786 242938 261022 243174
rect 260466 242618 260702 242854
rect 260786 242618 261022 242854
rect 260466 224938 260702 225174
rect 260786 224938 261022 225174
rect 260466 224618 260702 224854
rect 260786 224618 261022 224854
rect 260466 206938 260702 207174
rect 260786 206938 261022 207174
rect 260466 206618 260702 206854
rect 260786 206618 261022 206854
rect 260466 188938 260702 189174
rect 260786 188938 261022 189174
rect 260466 188618 260702 188854
rect 260786 188618 261022 188854
rect 260466 170938 260702 171174
rect 260786 170938 261022 171174
rect 260466 170618 260702 170854
rect 260786 170618 261022 170854
rect 260466 152938 260702 153174
rect 260786 152938 261022 153174
rect 260466 152618 260702 152854
rect 260786 152618 261022 152854
rect 260466 134938 260702 135174
rect 260786 134938 261022 135174
rect 260466 134618 260702 134854
rect 260786 134618 261022 134854
rect 260466 116938 260702 117174
rect 260786 116938 261022 117174
rect 260466 116618 260702 116854
rect 260786 116618 261022 116854
rect 260466 98938 260702 99174
rect 260786 98938 261022 99174
rect 260466 98618 260702 98854
rect 260786 98618 261022 98854
rect 260466 80938 260702 81174
rect 260786 80938 261022 81174
rect 260466 80618 260702 80854
rect 260786 80618 261022 80854
rect 260466 62938 260702 63174
rect 260786 62938 261022 63174
rect 260466 62618 260702 62854
rect 260786 62618 261022 62854
rect 260466 44938 260702 45174
rect 260786 44938 261022 45174
rect 260466 44618 260702 44854
rect 260786 44618 261022 44854
rect 260466 26938 260702 27174
rect 260786 26938 261022 27174
rect 260466 26618 260702 26854
rect 260786 26618 261022 26854
rect 260466 8938 260702 9174
rect 260786 8938 261022 9174
rect 260466 8618 260702 8854
rect 260786 8618 261022 8854
rect 260466 -2052 260702 -1816
rect 260786 -2052 261022 -1816
rect 260466 -2372 260702 -2136
rect 260786 -2372 261022 -2136
rect 264186 462776 264422 463012
rect 264506 462776 264742 463012
rect 264186 462456 264422 462692
rect 264506 462456 264742 462692
rect 264186 444658 264422 444894
rect 264506 444658 264742 444894
rect 264186 444338 264422 444574
rect 264506 444338 264742 444574
rect 264186 426658 264422 426894
rect 264506 426658 264742 426894
rect 264186 426338 264422 426574
rect 264506 426338 264742 426574
rect 264186 408658 264422 408894
rect 264506 408658 264742 408894
rect 264186 408338 264422 408574
rect 264506 408338 264742 408574
rect 264186 390658 264422 390894
rect 264506 390658 264742 390894
rect 264186 390338 264422 390574
rect 264506 390338 264742 390574
rect 264186 372658 264422 372894
rect 264506 372658 264742 372894
rect 264186 372338 264422 372574
rect 264506 372338 264742 372574
rect 264186 354658 264422 354894
rect 264506 354658 264742 354894
rect 264186 354338 264422 354574
rect 264506 354338 264742 354574
rect 264186 336658 264422 336894
rect 264506 336658 264742 336894
rect 264186 336338 264422 336574
rect 264506 336338 264742 336574
rect 264186 318658 264422 318894
rect 264506 318658 264742 318894
rect 264186 318338 264422 318574
rect 264506 318338 264742 318574
rect 264186 300658 264422 300894
rect 264506 300658 264742 300894
rect 264186 300338 264422 300574
rect 264506 300338 264742 300574
rect 264186 282658 264422 282894
rect 264506 282658 264742 282894
rect 264186 282338 264422 282574
rect 264506 282338 264742 282574
rect 264186 264658 264422 264894
rect 264506 264658 264742 264894
rect 264186 264338 264422 264574
rect 264506 264338 264742 264574
rect 264186 246658 264422 246894
rect 264506 246658 264742 246894
rect 264186 246338 264422 246574
rect 264506 246338 264742 246574
rect 264186 228658 264422 228894
rect 264506 228658 264742 228894
rect 264186 228338 264422 228574
rect 264506 228338 264742 228574
rect 264186 210658 264422 210894
rect 264506 210658 264742 210894
rect 264186 210338 264422 210574
rect 264506 210338 264742 210574
rect 264186 192658 264422 192894
rect 264506 192658 264742 192894
rect 264186 192338 264422 192574
rect 264506 192338 264742 192574
rect 264186 174658 264422 174894
rect 264506 174658 264742 174894
rect 264186 174338 264422 174574
rect 264506 174338 264742 174574
rect 264186 156658 264422 156894
rect 264506 156658 264742 156894
rect 264186 156338 264422 156574
rect 264506 156338 264742 156574
rect 264186 138658 264422 138894
rect 264506 138658 264742 138894
rect 264186 138338 264422 138574
rect 264506 138338 264742 138574
rect 264186 120658 264422 120894
rect 264506 120658 264742 120894
rect 264186 120338 264422 120574
rect 264506 120338 264742 120574
rect 264186 102658 264422 102894
rect 264506 102658 264742 102894
rect 264186 102338 264422 102574
rect 264506 102338 264742 102574
rect 264186 84658 264422 84894
rect 264506 84658 264742 84894
rect 264186 84338 264422 84574
rect 264506 84338 264742 84574
rect 264186 66658 264422 66894
rect 264506 66658 264742 66894
rect 264186 66338 264422 66574
rect 264506 66338 264742 66574
rect 264186 48658 264422 48894
rect 264506 48658 264742 48894
rect 264186 48338 264422 48574
rect 264506 48338 264742 48574
rect 264186 30658 264422 30894
rect 264506 30658 264742 30894
rect 264186 30338 264422 30574
rect 264506 30338 264742 30574
rect 264186 12658 264422 12894
rect 264506 12658 264742 12894
rect 264186 12338 264422 12574
rect 264506 12338 264742 12574
rect 264186 -3012 264422 -2776
rect 264506 -3012 264742 -2776
rect 264186 -3332 264422 -3096
rect 264506 -3332 264742 -3096
rect 267906 463736 268142 463972
rect 268226 463736 268462 463972
rect 267906 463416 268142 463652
rect 268226 463416 268462 463652
rect 267906 448378 268142 448614
rect 268226 448378 268462 448614
rect 267906 448058 268142 448294
rect 268226 448058 268462 448294
rect 267906 430378 268142 430614
rect 268226 430378 268462 430614
rect 267906 430058 268142 430294
rect 268226 430058 268462 430294
rect 267906 412378 268142 412614
rect 268226 412378 268462 412614
rect 267906 412058 268142 412294
rect 268226 412058 268462 412294
rect 267906 394378 268142 394614
rect 268226 394378 268462 394614
rect 267906 394058 268142 394294
rect 268226 394058 268462 394294
rect 267906 376378 268142 376614
rect 268226 376378 268462 376614
rect 267906 376058 268142 376294
rect 268226 376058 268462 376294
rect 267906 358378 268142 358614
rect 268226 358378 268462 358614
rect 267906 358058 268142 358294
rect 268226 358058 268462 358294
rect 267906 340378 268142 340614
rect 268226 340378 268462 340614
rect 267906 340058 268142 340294
rect 268226 340058 268462 340294
rect 267906 322378 268142 322614
rect 268226 322378 268462 322614
rect 267906 322058 268142 322294
rect 268226 322058 268462 322294
rect 267906 304378 268142 304614
rect 268226 304378 268462 304614
rect 267906 304058 268142 304294
rect 268226 304058 268462 304294
rect 267906 286378 268142 286614
rect 268226 286378 268462 286614
rect 267906 286058 268142 286294
rect 268226 286058 268462 286294
rect 267906 268378 268142 268614
rect 268226 268378 268462 268614
rect 267906 268058 268142 268294
rect 268226 268058 268462 268294
rect 267906 250378 268142 250614
rect 268226 250378 268462 250614
rect 267906 250058 268142 250294
rect 268226 250058 268462 250294
rect 267906 232378 268142 232614
rect 268226 232378 268462 232614
rect 267906 232058 268142 232294
rect 268226 232058 268462 232294
rect 267906 214378 268142 214614
rect 268226 214378 268462 214614
rect 267906 214058 268142 214294
rect 268226 214058 268462 214294
rect 267906 196378 268142 196614
rect 268226 196378 268462 196614
rect 267906 196058 268142 196294
rect 268226 196058 268462 196294
rect 267906 178378 268142 178614
rect 268226 178378 268462 178614
rect 267906 178058 268142 178294
rect 268226 178058 268462 178294
rect 267906 160378 268142 160614
rect 268226 160378 268462 160614
rect 267906 160058 268142 160294
rect 268226 160058 268462 160294
rect 267906 142378 268142 142614
rect 268226 142378 268462 142614
rect 267906 142058 268142 142294
rect 268226 142058 268462 142294
rect 267906 124378 268142 124614
rect 268226 124378 268462 124614
rect 267906 124058 268142 124294
rect 268226 124058 268462 124294
rect 267906 106378 268142 106614
rect 268226 106378 268462 106614
rect 267906 106058 268142 106294
rect 268226 106058 268462 106294
rect 267906 88378 268142 88614
rect 268226 88378 268462 88614
rect 267906 88058 268142 88294
rect 268226 88058 268462 88294
rect 267906 70378 268142 70614
rect 268226 70378 268462 70614
rect 267906 70058 268142 70294
rect 268226 70058 268462 70294
rect 267906 52378 268142 52614
rect 268226 52378 268462 52614
rect 267906 52058 268142 52294
rect 268226 52058 268462 52294
rect 267906 34378 268142 34614
rect 268226 34378 268462 34614
rect 267906 34058 268142 34294
rect 268226 34058 268462 34294
rect 267906 16378 268142 16614
rect 268226 16378 268462 16614
rect 267906 16058 268142 16294
rect 268226 16058 268462 16294
rect 267906 -3972 268142 -3736
rect 268226 -3972 268462 -3736
rect 267906 -4292 268142 -4056
rect 268226 -4292 268462 -4056
rect 274746 460856 274982 461092
rect 275066 460856 275302 461092
rect 274746 460536 274982 460772
rect 275066 460536 275302 460772
rect 274746 455218 274982 455454
rect 275066 455218 275302 455454
rect 274746 454898 274982 455134
rect 275066 454898 275302 455134
rect 274746 437218 274982 437454
rect 275066 437218 275302 437454
rect 274746 436898 274982 437134
rect 275066 436898 275302 437134
rect 274746 419218 274982 419454
rect 275066 419218 275302 419454
rect 274746 418898 274982 419134
rect 275066 418898 275302 419134
rect 274746 401218 274982 401454
rect 275066 401218 275302 401454
rect 274746 400898 274982 401134
rect 275066 400898 275302 401134
rect 274746 383218 274982 383454
rect 275066 383218 275302 383454
rect 274746 382898 274982 383134
rect 275066 382898 275302 383134
rect 274746 365218 274982 365454
rect 275066 365218 275302 365454
rect 274746 364898 274982 365134
rect 275066 364898 275302 365134
rect 274746 347218 274982 347454
rect 275066 347218 275302 347454
rect 274746 346898 274982 347134
rect 275066 346898 275302 347134
rect 274746 329218 274982 329454
rect 275066 329218 275302 329454
rect 274746 328898 274982 329134
rect 275066 328898 275302 329134
rect 274746 311218 274982 311454
rect 275066 311218 275302 311454
rect 274746 310898 274982 311134
rect 275066 310898 275302 311134
rect 274746 293218 274982 293454
rect 275066 293218 275302 293454
rect 274746 292898 274982 293134
rect 275066 292898 275302 293134
rect 274746 275218 274982 275454
rect 275066 275218 275302 275454
rect 274746 274898 274982 275134
rect 275066 274898 275302 275134
rect 274746 257218 274982 257454
rect 275066 257218 275302 257454
rect 274746 256898 274982 257134
rect 275066 256898 275302 257134
rect 274746 239218 274982 239454
rect 275066 239218 275302 239454
rect 274746 238898 274982 239134
rect 275066 238898 275302 239134
rect 274746 221218 274982 221454
rect 275066 221218 275302 221454
rect 274746 220898 274982 221134
rect 275066 220898 275302 221134
rect 274746 203218 274982 203454
rect 275066 203218 275302 203454
rect 274746 202898 274982 203134
rect 275066 202898 275302 203134
rect 274746 185218 274982 185454
rect 275066 185218 275302 185454
rect 274746 184898 274982 185134
rect 275066 184898 275302 185134
rect 274746 167218 274982 167454
rect 275066 167218 275302 167454
rect 274746 166898 274982 167134
rect 275066 166898 275302 167134
rect 274746 149218 274982 149454
rect 275066 149218 275302 149454
rect 274746 148898 274982 149134
rect 275066 148898 275302 149134
rect 274746 131218 274982 131454
rect 275066 131218 275302 131454
rect 274746 130898 274982 131134
rect 275066 130898 275302 131134
rect 274746 113218 274982 113454
rect 275066 113218 275302 113454
rect 274746 112898 274982 113134
rect 275066 112898 275302 113134
rect 274746 95218 274982 95454
rect 275066 95218 275302 95454
rect 274746 94898 274982 95134
rect 275066 94898 275302 95134
rect 274746 77218 274982 77454
rect 275066 77218 275302 77454
rect 274746 76898 274982 77134
rect 275066 76898 275302 77134
rect 274746 59218 274982 59454
rect 275066 59218 275302 59454
rect 274746 58898 274982 59134
rect 275066 58898 275302 59134
rect 274746 41218 274982 41454
rect 275066 41218 275302 41454
rect 274746 40898 274982 41134
rect 275066 40898 275302 41134
rect 274746 23218 274982 23454
rect 275066 23218 275302 23454
rect 274746 22898 274982 23134
rect 275066 22898 275302 23134
rect 274746 5218 274982 5454
rect 275066 5218 275302 5454
rect 274746 4898 274982 5134
rect 275066 4898 275302 5134
rect 274746 -1092 274982 -856
rect 275066 -1092 275302 -856
rect 274746 -1412 274982 -1176
rect 275066 -1412 275302 -1176
rect 278466 461816 278702 462052
rect 278786 461816 279022 462052
rect 278466 461496 278702 461732
rect 278786 461496 279022 461732
rect 278466 440938 278702 441174
rect 278786 440938 279022 441174
rect 278466 440618 278702 440854
rect 278786 440618 279022 440854
rect 278466 422938 278702 423174
rect 278786 422938 279022 423174
rect 278466 422618 278702 422854
rect 278786 422618 279022 422854
rect 278466 404938 278702 405174
rect 278786 404938 279022 405174
rect 278466 404618 278702 404854
rect 278786 404618 279022 404854
rect 278466 386938 278702 387174
rect 278786 386938 279022 387174
rect 278466 386618 278702 386854
rect 278786 386618 279022 386854
rect 278466 368938 278702 369174
rect 278786 368938 279022 369174
rect 278466 368618 278702 368854
rect 278786 368618 279022 368854
rect 278466 350938 278702 351174
rect 278786 350938 279022 351174
rect 278466 350618 278702 350854
rect 278786 350618 279022 350854
rect 278466 332938 278702 333174
rect 278786 332938 279022 333174
rect 278466 332618 278702 332854
rect 278786 332618 279022 332854
rect 278466 314938 278702 315174
rect 278786 314938 279022 315174
rect 278466 314618 278702 314854
rect 278786 314618 279022 314854
rect 278466 296938 278702 297174
rect 278786 296938 279022 297174
rect 278466 296618 278702 296854
rect 278786 296618 279022 296854
rect 278466 278938 278702 279174
rect 278786 278938 279022 279174
rect 278466 278618 278702 278854
rect 278786 278618 279022 278854
rect 278466 260938 278702 261174
rect 278786 260938 279022 261174
rect 278466 260618 278702 260854
rect 278786 260618 279022 260854
rect 278466 242938 278702 243174
rect 278786 242938 279022 243174
rect 278466 242618 278702 242854
rect 278786 242618 279022 242854
rect 278466 224938 278702 225174
rect 278786 224938 279022 225174
rect 278466 224618 278702 224854
rect 278786 224618 279022 224854
rect 278466 206938 278702 207174
rect 278786 206938 279022 207174
rect 278466 206618 278702 206854
rect 278786 206618 279022 206854
rect 278466 188938 278702 189174
rect 278786 188938 279022 189174
rect 278466 188618 278702 188854
rect 278786 188618 279022 188854
rect 278466 170938 278702 171174
rect 278786 170938 279022 171174
rect 278466 170618 278702 170854
rect 278786 170618 279022 170854
rect 278466 152938 278702 153174
rect 278786 152938 279022 153174
rect 278466 152618 278702 152854
rect 278786 152618 279022 152854
rect 278466 134938 278702 135174
rect 278786 134938 279022 135174
rect 278466 134618 278702 134854
rect 278786 134618 279022 134854
rect 278466 116938 278702 117174
rect 278786 116938 279022 117174
rect 278466 116618 278702 116854
rect 278786 116618 279022 116854
rect 278466 98938 278702 99174
rect 278786 98938 279022 99174
rect 278466 98618 278702 98854
rect 278786 98618 279022 98854
rect 278466 80938 278702 81174
rect 278786 80938 279022 81174
rect 278466 80618 278702 80854
rect 278786 80618 279022 80854
rect 278466 62938 278702 63174
rect 278786 62938 279022 63174
rect 278466 62618 278702 62854
rect 278786 62618 279022 62854
rect 278466 44938 278702 45174
rect 278786 44938 279022 45174
rect 278466 44618 278702 44854
rect 278786 44618 279022 44854
rect 278466 26938 278702 27174
rect 278786 26938 279022 27174
rect 278466 26618 278702 26854
rect 278786 26618 279022 26854
rect 278466 8938 278702 9174
rect 278786 8938 279022 9174
rect 278466 8618 278702 8854
rect 278786 8618 279022 8854
rect 278466 -2052 278702 -1816
rect 278786 -2052 279022 -1816
rect 278466 -2372 278702 -2136
rect 278786 -2372 279022 -2136
rect 282186 462776 282422 463012
rect 282506 462776 282742 463012
rect 282186 462456 282422 462692
rect 282506 462456 282742 462692
rect 282186 444658 282422 444894
rect 282506 444658 282742 444894
rect 282186 444338 282422 444574
rect 282506 444338 282742 444574
rect 282186 426658 282422 426894
rect 282506 426658 282742 426894
rect 282186 426338 282422 426574
rect 282506 426338 282742 426574
rect 282186 408658 282422 408894
rect 282506 408658 282742 408894
rect 282186 408338 282422 408574
rect 282506 408338 282742 408574
rect 282186 390658 282422 390894
rect 282506 390658 282742 390894
rect 282186 390338 282422 390574
rect 282506 390338 282742 390574
rect 282186 372658 282422 372894
rect 282506 372658 282742 372894
rect 282186 372338 282422 372574
rect 282506 372338 282742 372574
rect 282186 354658 282422 354894
rect 282506 354658 282742 354894
rect 282186 354338 282422 354574
rect 282506 354338 282742 354574
rect 282186 336658 282422 336894
rect 282506 336658 282742 336894
rect 282186 336338 282422 336574
rect 282506 336338 282742 336574
rect 282186 318658 282422 318894
rect 282506 318658 282742 318894
rect 282186 318338 282422 318574
rect 282506 318338 282742 318574
rect 282186 300658 282422 300894
rect 282506 300658 282742 300894
rect 282186 300338 282422 300574
rect 282506 300338 282742 300574
rect 282186 282658 282422 282894
rect 282506 282658 282742 282894
rect 282186 282338 282422 282574
rect 282506 282338 282742 282574
rect 282186 264658 282422 264894
rect 282506 264658 282742 264894
rect 282186 264338 282422 264574
rect 282506 264338 282742 264574
rect 282186 246658 282422 246894
rect 282506 246658 282742 246894
rect 282186 246338 282422 246574
rect 282506 246338 282742 246574
rect 282186 228658 282422 228894
rect 282506 228658 282742 228894
rect 282186 228338 282422 228574
rect 282506 228338 282742 228574
rect 282186 210658 282422 210894
rect 282506 210658 282742 210894
rect 282186 210338 282422 210574
rect 282506 210338 282742 210574
rect 282186 192658 282422 192894
rect 282506 192658 282742 192894
rect 282186 192338 282422 192574
rect 282506 192338 282742 192574
rect 282186 174658 282422 174894
rect 282506 174658 282742 174894
rect 282186 174338 282422 174574
rect 282506 174338 282742 174574
rect 282186 156658 282422 156894
rect 282506 156658 282742 156894
rect 282186 156338 282422 156574
rect 282506 156338 282742 156574
rect 282186 138658 282422 138894
rect 282506 138658 282742 138894
rect 282186 138338 282422 138574
rect 282506 138338 282742 138574
rect 282186 120658 282422 120894
rect 282506 120658 282742 120894
rect 282186 120338 282422 120574
rect 282506 120338 282742 120574
rect 282186 102658 282422 102894
rect 282506 102658 282742 102894
rect 282186 102338 282422 102574
rect 282506 102338 282742 102574
rect 282186 84658 282422 84894
rect 282506 84658 282742 84894
rect 282186 84338 282422 84574
rect 282506 84338 282742 84574
rect 282186 66658 282422 66894
rect 282506 66658 282742 66894
rect 282186 66338 282422 66574
rect 282506 66338 282742 66574
rect 282186 48658 282422 48894
rect 282506 48658 282742 48894
rect 282186 48338 282422 48574
rect 282506 48338 282742 48574
rect 282186 30658 282422 30894
rect 282506 30658 282742 30894
rect 282186 30338 282422 30574
rect 282506 30338 282742 30574
rect 282186 12658 282422 12894
rect 282506 12658 282742 12894
rect 282186 12338 282422 12574
rect 282506 12338 282742 12574
rect 282186 -3012 282422 -2776
rect 282506 -3012 282742 -2776
rect 282186 -3332 282422 -3096
rect 282506 -3332 282742 -3096
rect 285906 463736 286142 463972
rect 286226 463736 286462 463972
rect 285906 463416 286142 463652
rect 286226 463416 286462 463652
rect 285906 448378 286142 448614
rect 286226 448378 286462 448614
rect 285906 448058 286142 448294
rect 286226 448058 286462 448294
rect 285906 430378 286142 430614
rect 286226 430378 286462 430614
rect 285906 430058 286142 430294
rect 286226 430058 286462 430294
rect 285906 412378 286142 412614
rect 286226 412378 286462 412614
rect 285906 412058 286142 412294
rect 286226 412058 286462 412294
rect 285906 394378 286142 394614
rect 286226 394378 286462 394614
rect 285906 394058 286142 394294
rect 286226 394058 286462 394294
rect 285906 376378 286142 376614
rect 286226 376378 286462 376614
rect 285906 376058 286142 376294
rect 286226 376058 286462 376294
rect 285906 358378 286142 358614
rect 286226 358378 286462 358614
rect 285906 358058 286142 358294
rect 286226 358058 286462 358294
rect 285906 340378 286142 340614
rect 286226 340378 286462 340614
rect 285906 340058 286142 340294
rect 286226 340058 286462 340294
rect 285906 322378 286142 322614
rect 286226 322378 286462 322614
rect 285906 322058 286142 322294
rect 286226 322058 286462 322294
rect 285906 304378 286142 304614
rect 286226 304378 286462 304614
rect 285906 304058 286142 304294
rect 286226 304058 286462 304294
rect 285906 286378 286142 286614
rect 286226 286378 286462 286614
rect 285906 286058 286142 286294
rect 286226 286058 286462 286294
rect 285906 268378 286142 268614
rect 286226 268378 286462 268614
rect 285906 268058 286142 268294
rect 286226 268058 286462 268294
rect 285906 250378 286142 250614
rect 286226 250378 286462 250614
rect 285906 250058 286142 250294
rect 286226 250058 286462 250294
rect 285906 232378 286142 232614
rect 286226 232378 286462 232614
rect 285906 232058 286142 232294
rect 286226 232058 286462 232294
rect 285906 214378 286142 214614
rect 286226 214378 286462 214614
rect 285906 214058 286142 214294
rect 286226 214058 286462 214294
rect 285906 196378 286142 196614
rect 286226 196378 286462 196614
rect 285906 196058 286142 196294
rect 286226 196058 286462 196294
rect 285906 178378 286142 178614
rect 286226 178378 286462 178614
rect 285906 178058 286142 178294
rect 286226 178058 286462 178294
rect 285906 160378 286142 160614
rect 286226 160378 286462 160614
rect 285906 160058 286142 160294
rect 286226 160058 286462 160294
rect 285906 142378 286142 142614
rect 286226 142378 286462 142614
rect 285906 142058 286142 142294
rect 286226 142058 286462 142294
rect 285906 124378 286142 124614
rect 286226 124378 286462 124614
rect 285906 124058 286142 124294
rect 286226 124058 286462 124294
rect 285906 106378 286142 106614
rect 286226 106378 286462 106614
rect 285906 106058 286142 106294
rect 286226 106058 286462 106294
rect 285906 88378 286142 88614
rect 286226 88378 286462 88614
rect 285906 88058 286142 88294
rect 286226 88058 286462 88294
rect 285906 70378 286142 70614
rect 286226 70378 286462 70614
rect 285906 70058 286142 70294
rect 286226 70058 286462 70294
rect 285906 52378 286142 52614
rect 286226 52378 286462 52614
rect 285906 52058 286142 52294
rect 286226 52058 286462 52294
rect 285906 34378 286142 34614
rect 286226 34378 286462 34614
rect 285906 34058 286142 34294
rect 286226 34058 286462 34294
rect 285906 16378 286142 16614
rect 286226 16378 286462 16614
rect 285906 16058 286142 16294
rect 286226 16058 286462 16294
rect 285906 -3972 286142 -3736
rect 286226 -3972 286462 -3736
rect 285906 -4292 286142 -4056
rect 286226 -4292 286462 -4056
rect 292746 460856 292982 461092
rect 293066 460856 293302 461092
rect 292746 460536 292982 460772
rect 293066 460536 293302 460772
rect 292746 455218 292982 455454
rect 293066 455218 293302 455454
rect 292746 454898 292982 455134
rect 293066 454898 293302 455134
rect 292746 437218 292982 437454
rect 293066 437218 293302 437454
rect 292746 436898 292982 437134
rect 293066 436898 293302 437134
rect 292746 419218 292982 419454
rect 293066 419218 293302 419454
rect 292746 418898 292982 419134
rect 293066 418898 293302 419134
rect 292746 401218 292982 401454
rect 293066 401218 293302 401454
rect 292746 400898 292982 401134
rect 293066 400898 293302 401134
rect 292746 383218 292982 383454
rect 293066 383218 293302 383454
rect 292746 382898 292982 383134
rect 293066 382898 293302 383134
rect 292746 365218 292982 365454
rect 293066 365218 293302 365454
rect 292746 364898 292982 365134
rect 293066 364898 293302 365134
rect 292746 347218 292982 347454
rect 293066 347218 293302 347454
rect 292746 346898 292982 347134
rect 293066 346898 293302 347134
rect 292746 329218 292982 329454
rect 293066 329218 293302 329454
rect 292746 328898 292982 329134
rect 293066 328898 293302 329134
rect 292746 311218 292982 311454
rect 293066 311218 293302 311454
rect 292746 310898 292982 311134
rect 293066 310898 293302 311134
rect 292746 293218 292982 293454
rect 293066 293218 293302 293454
rect 292746 292898 292982 293134
rect 293066 292898 293302 293134
rect 292746 275218 292982 275454
rect 293066 275218 293302 275454
rect 292746 274898 292982 275134
rect 293066 274898 293302 275134
rect 292746 257218 292982 257454
rect 293066 257218 293302 257454
rect 292746 256898 292982 257134
rect 293066 256898 293302 257134
rect 292746 239218 292982 239454
rect 293066 239218 293302 239454
rect 292746 238898 292982 239134
rect 293066 238898 293302 239134
rect 292746 221218 292982 221454
rect 293066 221218 293302 221454
rect 292746 220898 292982 221134
rect 293066 220898 293302 221134
rect 292746 203218 292982 203454
rect 293066 203218 293302 203454
rect 292746 202898 292982 203134
rect 293066 202898 293302 203134
rect 292746 185218 292982 185454
rect 293066 185218 293302 185454
rect 292746 184898 292982 185134
rect 293066 184898 293302 185134
rect 292746 167218 292982 167454
rect 293066 167218 293302 167454
rect 292746 166898 292982 167134
rect 293066 166898 293302 167134
rect 292746 149218 292982 149454
rect 293066 149218 293302 149454
rect 292746 148898 292982 149134
rect 293066 148898 293302 149134
rect 292746 131218 292982 131454
rect 293066 131218 293302 131454
rect 292746 130898 292982 131134
rect 293066 130898 293302 131134
rect 292746 113218 292982 113454
rect 293066 113218 293302 113454
rect 292746 112898 292982 113134
rect 293066 112898 293302 113134
rect 292746 95218 292982 95454
rect 293066 95218 293302 95454
rect 292746 94898 292982 95134
rect 293066 94898 293302 95134
rect 292746 77218 292982 77454
rect 293066 77218 293302 77454
rect 292746 76898 292982 77134
rect 293066 76898 293302 77134
rect 292746 59218 292982 59454
rect 293066 59218 293302 59454
rect 292746 58898 292982 59134
rect 293066 58898 293302 59134
rect 292746 41218 292982 41454
rect 293066 41218 293302 41454
rect 292746 40898 292982 41134
rect 293066 40898 293302 41134
rect 292746 23218 292982 23454
rect 293066 23218 293302 23454
rect 292746 22898 292982 23134
rect 293066 22898 293302 23134
rect 292746 5218 292982 5454
rect 293066 5218 293302 5454
rect 292746 4898 292982 5134
rect 293066 4898 293302 5134
rect 292746 -1092 292982 -856
rect 293066 -1092 293302 -856
rect 292746 -1412 292982 -1176
rect 293066 -1412 293302 -1176
rect 296466 461816 296702 462052
rect 296786 461816 297022 462052
rect 296466 461496 296702 461732
rect 296786 461496 297022 461732
rect 296466 440938 296702 441174
rect 296786 440938 297022 441174
rect 296466 440618 296702 440854
rect 296786 440618 297022 440854
rect 296466 422938 296702 423174
rect 296786 422938 297022 423174
rect 296466 422618 296702 422854
rect 296786 422618 297022 422854
rect 296466 404938 296702 405174
rect 296786 404938 297022 405174
rect 296466 404618 296702 404854
rect 296786 404618 297022 404854
rect 296466 386938 296702 387174
rect 296786 386938 297022 387174
rect 296466 386618 296702 386854
rect 296786 386618 297022 386854
rect 296466 368938 296702 369174
rect 296786 368938 297022 369174
rect 296466 368618 296702 368854
rect 296786 368618 297022 368854
rect 296466 350938 296702 351174
rect 296786 350938 297022 351174
rect 296466 350618 296702 350854
rect 296786 350618 297022 350854
rect 296466 332938 296702 333174
rect 296786 332938 297022 333174
rect 296466 332618 296702 332854
rect 296786 332618 297022 332854
rect 296466 314938 296702 315174
rect 296786 314938 297022 315174
rect 296466 314618 296702 314854
rect 296786 314618 297022 314854
rect 296466 296938 296702 297174
rect 296786 296938 297022 297174
rect 296466 296618 296702 296854
rect 296786 296618 297022 296854
rect 296466 278938 296702 279174
rect 296786 278938 297022 279174
rect 296466 278618 296702 278854
rect 296786 278618 297022 278854
rect 296466 260938 296702 261174
rect 296786 260938 297022 261174
rect 296466 260618 296702 260854
rect 296786 260618 297022 260854
rect 296466 242938 296702 243174
rect 296786 242938 297022 243174
rect 296466 242618 296702 242854
rect 296786 242618 297022 242854
rect 296466 224938 296702 225174
rect 296786 224938 297022 225174
rect 296466 224618 296702 224854
rect 296786 224618 297022 224854
rect 296466 206938 296702 207174
rect 296786 206938 297022 207174
rect 296466 206618 296702 206854
rect 296786 206618 297022 206854
rect 296466 188938 296702 189174
rect 296786 188938 297022 189174
rect 296466 188618 296702 188854
rect 296786 188618 297022 188854
rect 296466 170938 296702 171174
rect 296786 170938 297022 171174
rect 296466 170618 296702 170854
rect 296786 170618 297022 170854
rect 296466 152938 296702 153174
rect 296786 152938 297022 153174
rect 296466 152618 296702 152854
rect 296786 152618 297022 152854
rect 296466 134938 296702 135174
rect 296786 134938 297022 135174
rect 296466 134618 296702 134854
rect 296786 134618 297022 134854
rect 296466 116938 296702 117174
rect 296786 116938 297022 117174
rect 296466 116618 296702 116854
rect 296786 116618 297022 116854
rect 296466 98938 296702 99174
rect 296786 98938 297022 99174
rect 296466 98618 296702 98854
rect 296786 98618 297022 98854
rect 296466 80938 296702 81174
rect 296786 80938 297022 81174
rect 296466 80618 296702 80854
rect 296786 80618 297022 80854
rect 296466 62938 296702 63174
rect 296786 62938 297022 63174
rect 296466 62618 296702 62854
rect 296786 62618 297022 62854
rect 296466 44938 296702 45174
rect 296786 44938 297022 45174
rect 296466 44618 296702 44854
rect 296786 44618 297022 44854
rect 296466 26938 296702 27174
rect 296786 26938 297022 27174
rect 296466 26618 296702 26854
rect 296786 26618 297022 26854
rect 296466 8938 296702 9174
rect 296786 8938 297022 9174
rect 296466 8618 296702 8854
rect 296786 8618 297022 8854
rect 296466 -2052 296702 -1816
rect 296786 -2052 297022 -1816
rect 296466 -2372 296702 -2136
rect 296786 -2372 297022 -2136
rect 300186 462776 300422 463012
rect 300506 462776 300742 463012
rect 300186 462456 300422 462692
rect 300506 462456 300742 462692
rect 300186 444658 300422 444894
rect 300506 444658 300742 444894
rect 300186 444338 300422 444574
rect 300506 444338 300742 444574
rect 300186 426658 300422 426894
rect 300506 426658 300742 426894
rect 300186 426338 300422 426574
rect 300506 426338 300742 426574
rect 300186 408658 300422 408894
rect 300506 408658 300742 408894
rect 300186 408338 300422 408574
rect 300506 408338 300742 408574
rect 300186 390658 300422 390894
rect 300506 390658 300742 390894
rect 300186 390338 300422 390574
rect 300506 390338 300742 390574
rect 300186 372658 300422 372894
rect 300506 372658 300742 372894
rect 300186 372338 300422 372574
rect 300506 372338 300742 372574
rect 300186 354658 300422 354894
rect 300506 354658 300742 354894
rect 300186 354338 300422 354574
rect 300506 354338 300742 354574
rect 300186 336658 300422 336894
rect 300506 336658 300742 336894
rect 300186 336338 300422 336574
rect 300506 336338 300742 336574
rect 300186 318658 300422 318894
rect 300506 318658 300742 318894
rect 300186 318338 300422 318574
rect 300506 318338 300742 318574
rect 300186 300658 300422 300894
rect 300506 300658 300742 300894
rect 300186 300338 300422 300574
rect 300506 300338 300742 300574
rect 300186 282658 300422 282894
rect 300506 282658 300742 282894
rect 300186 282338 300422 282574
rect 300506 282338 300742 282574
rect 300186 264658 300422 264894
rect 300506 264658 300742 264894
rect 300186 264338 300422 264574
rect 300506 264338 300742 264574
rect 300186 246658 300422 246894
rect 300506 246658 300742 246894
rect 300186 246338 300422 246574
rect 300506 246338 300742 246574
rect 300186 228658 300422 228894
rect 300506 228658 300742 228894
rect 300186 228338 300422 228574
rect 300506 228338 300742 228574
rect 300186 210658 300422 210894
rect 300506 210658 300742 210894
rect 300186 210338 300422 210574
rect 300506 210338 300742 210574
rect 300186 192658 300422 192894
rect 300506 192658 300742 192894
rect 300186 192338 300422 192574
rect 300506 192338 300742 192574
rect 300186 174658 300422 174894
rect 300506 174658 300742 174894
rect 300186 174338 300422 174574
rect 300506 174338 300742 174574
rect 300186 156658 300422 156894
rect 300506 156658 300742 156894
rect 300186 156338 300422 156574
rect 300506 156338 300742 156574
rect 300186 138658 300422 138894
rect 300506 138658 300742 138894
rect 300186 138338 300422 138574
rect 300506 138338 300742 138574
rect 300186 120658 300422 120894
rect 300506 120658 300742 120894
rect 300186 120338 300422 120574
rect 300506 120338 300742 120574
rect 300186 102658 300422 102894
rect 300506 102658 300742 102894
rect 300186 102338 300422 102574
rect 300506 102338 300742 102574
rect 300186 84658 300422 84894
rect 300506 84658 300742 84894
rect 300186 84338 300422 84574
rect 300506 84338 300742 84574
rect 300186 66658 300422 66894
rect 300506 66658 300742 66894
rect 300186 66338 300422 66574
rect 300506 66338 300742 66574
rect 300186 48658 300422 48894
rect 300506 48658 300742 48894
rect 300186 48338 300422 48574
rect 300506 48338 300742 48574
rect 300186 30658 300422 30894
rect 300506 30658 300742 30894
rect 300186 30338 300422 30574
rect 300506 30338 300742 30574
rect 300186 12658 300422 12894
rect 300506 12658 300742 12894
rect 300186 12338 300422 12574
rect 300506 12338 300742 12574
rect 300186 -3012 300422 -2776
rect 300506 -3012 300742 -2776
rect 300186 -3332 300422 -3096
rect 300506 -3332 300742 -3096
rect 303906 463736 304142 463972
rect 304226 463736 304462 463972
rect 303906 463416 304142 463652
rect 304226 463416 304462 463652
rect 303906 448378 304142 448614
rect 304226 448378 304462 448614
rect 303906 448058 304142 448294
rect 304226 448058 304462 448294
rect 303906 430378 304142 430614
rect 304226 430378 304462 430614
rect 303906 430058 304142 430294
rect 304226 430058 304462 430294
rect 303906 412378 304142 412614
rect 304226 412378 304462 412614
rect 303906 412058 304142 412294
rect 304226 412058 304462 412294
rect 303906 394378 304142 394614
rect 304226 394378 304462 394614
rect 303906 394058 304142 394294
rect 304226 394058 304462 394294
rect 303906 376378 304142 376614
rect 304226 376378 304462 376614
rect 303906 376058 304142 376294
rect 304226 376058 304462 376294
rect 303906 358378 304142 358614
rect 304226 358378 304462 358614
rect 303906 358058 304142 358294
rect 304226 358058 304462 358294
rect 303906 340378 304142 340614
rect 304226 340378 304462 340614
rect 303906 340058 304142 340294
rect 304226 340058 304462 340294
rect 303906 322378 304142 322614
rect 304226 322378 304462 322614
rect 303906 322058 304142 322294
rect 304226 322058 304462 322294
rect 303906 304378 304142 304614
rect 304226 304378 304462 304614
rect 303906 304058 304142 304294
rect 304226 304058 304462 304294
rect 303906 286378 304142 286614
rect 304226 286378 304462 286614
rect 303906 286058 304142 286294
rect 304226 286058 304462 286294
rect 303906 268378 304142 268614
rect 304226 268378 304462 268614
rect 303906 268058 304142 268294
rect 304226 268058 304462 268294
rect 303906 250378 304142 250614
rect 304226 250378 304462 250614
rect 303906 250058 304142 250294
rect 304226 250058 304462 250294
rect 303906 232378 304142 232614
rect 304226 232378 304462 232614
rect 303906 232058 304142 232294
rect 304226 232058 304462 232294
rect 303906 214378 304142 214614
rect 304226 214378 304462 214614
rect 303906 214058 304142 214294
rect 304226 214058 304462 214294
rect 303906 196378 304142 196614
rect 304226 196378 304462 196614
rect 303906 196058 304142 196294
rect 304226 196058 304462 196294
rect 303906 178378 304142 178614
rect 304226 178378 304462 178614
rect 303906 178058 304142 178294
rect 304226 178058 304462 178294
rect 303906 160378 304142 160614
rect 304226 160378 304462 160614
rect 303906 160058 304142 160294
rect 304226 160058 304462 160294
rect 303906 142378 304142 142614
rect 304226 142378 304462 142614
rect 303906 142058 304142 142294
rect 304226 142058 304462 142294
rect 303906 124378 304142 124614
rect 304226 124378 304462 124614
rect 303906 124058 304142 124294
rect 304226 124058 304462 124294
rect 303906 106378 304142 106614
rect 304226 106378 304462 106614
rect 303906 106058 304142 106294
rect 304226 106058 304462 106294
rect 303906 88378 304142 88614
rect 304226 88378 304462 88614
rect 303906 88058 304142 88294
rect 304226 88058 304462 88294
rect 303906 70378 304142 70614
rect 304226 70378 304462 70614
rect 303906 70058 304142 70294
rect 304226 70058 304462 70294
rect 303906 52378 304142 52614
rect 304226 52378 304462 52614
rect 303906 52058 304142 52294
rect 304226 52058 304462 52294
rect 303906 34378 304142 34614
rect 304226 34378 304462 34614
rect 303906 34058 304142 34294
rect 304226 34058 304462 34294
rect 303906 16378 304142 16614
rect 304226 16378 304462 16614
rect 303906 16058 304142 16294
rect 304226 16058 304462 16294
rect 303906 -3972 304142 -3736
rect 304226 -3972 304462 -3736
rect 303906 -4292 304142 -4056
rect 304226 -4292 304462 -4056
rect 310746 460856 310982 461092
rect 311066 460856 311302 461092
rect 310746 460536 310982 460772
rect 311066 460536 311302 460772
rect 310746 455218 310982 455454
rect 311066 455218 311302 455454
rect 310746 454898 310982 455134
rect 311066 454898 311302 455134
rect 310746 437218 310982 437454
rect 311066 437218 311302 437454
rect 310746 436898 310982 437134
rect 311066 436898 311302 437134
rect 310746 419218 310982 419454
rect 311066 419218 311302 419454
rect 310746 418898 310982 419134
rect 311066 418898 311302 419134
rect 310746 401218 310982 401454
rect 311066 401218 311302 401454
rect 310746 400898 310982 401134
rect 311066 400898 311302 401134
rect 310746 383218 310982 383454
rect 311066 383218 311302 383454
rect 310746 382898 310982 383134
rect 311066 382898 311302 383134
rect 310746 365218 310982 365454
rect 311066 365218 311302 365454
rect 310746 364898 310982 365134
rect 311066 364898 311302 365134
rect 310746 347218 310982 347454
rect 311066 347218 311302 347454
rect 310746 346898 310982 347134
rect 311066 346898 311302 347134
rect 310746 329218 310982 329454
rect 311066 329218 311302 329454
rect 310746 328898 310982 329134
rect 311066 328898 311302 329134
rect 310746 311218 310982 311454
rect 311066 311218 311302 311454
rect 310746 310898 310982 311134
rect 311066 310898 311302 311134
rect 310746 293218 310982 293454
rect 311066 293218 311302 293454
rect 310746 292898 310982 293134
rect 311066 292898 311302 293134
rect 310746 275218 310982 275454
rect 311066 275218 311302 275454
rect 310746 274898 310982 275134
rect 311066 274898 311302 275134
rect 310746 257218 310982 257454
rect 311066 257218 311302 257454
rect 310746 256898 310982 257134
rect 311066 256898 311302 257134
rect 310746 239218 310982 239454
rect 311066 239218 311302 239454
rect 310746 238898 310982 239134
rect 311066 238898 311302 239134
rect 310746 221218 310982 221454
rect 311066 221218 311302 221454
rect 310746 220898 310982 221134
rect 311066 220898 311302 221134
rect 310746 203218 310982 203454
rect 311066 203218 311302 203454
rect 310746 202898 310982 203134
rect 311066 202898 311302 203134
rect 310746 185218 310982 185454
rect 311066 185218 311302 185454
rect 310746 184898 310982 185134
rect 311066 184898 311302 185134
rect 310746 167218 310982 167454
rect 311066 167218 311302 167454
rect 310746 166898 310982 167134
rect 311066 166898 311302 167134
rect 310746 149218 310982 149454
rect 311066 149218 311302 149454
rect 310746 148898 310982 149134
rect 311066 148898 311302 149134
rect 310746 131218 310982 131454
rect 311066 131218 311302 131454
rect 310746 130898 310982 131134
rect 311066 130898 311302 131134
rect 310746 113218 310982 113454
rect 311066 113218 311302 113454
rect 310746 112898 310982 113134
rect 311066 112898 311302 113134
rect 310746 95218 310982 95454
rect 311066 95218 311302 95454
rect 310746 94898 310982 95134
rect 311066 94898 311302 95134
rect 310746 77218 310982 77454
rect 311066 77218 311302 77454
rect 310746 76898 310982 77134
rect 311066 76898 311302 77134
rect 310746 59218 310982 59454
rect 311066 59218 311302 59454
rect 310746 58898 310982 59134
rect 311066 58898 311302 59134
rect 310746 41218 310982 41454
rect 311066 41218 311302 41454
rect 310746 40898 310982 41134
rect 311066 40898 311302 41134
rect 310746 23218 310982 23454
rect 311066 23218 311302 23454
rect 310746 22898 310982 23134
rect 311066 22898 311302 23134
rect 310746 5218 310982 5454
rect 311066 5218 311302 5454
rect 310746 4898 310982 5134
rect 311066 4898 311302 5134
rect 310746 -1092 310982 -856
rect 311066 -1092 311302 -856
rect 310746 -1412 310982 -1176
rect 311066 -1412 311302 -1176
rect 314466 461816 314702 462052
rect 314786 461816 315022 462052
rect 314466 461496 314702 461732
rect 314786 461496 315022 461732
rect 314466 440938 314702 441174
rect 314786 440938 315022 441174
rect 314466 440618 314702 440854
rect 314786 440618 315022 440854
rect 314466 422938 314702 423174
rect 314786 422938 315022 423174
rect 314466 422618 314702 422854
rect 314786 422618 315022 422854
rect 314466 404938 314702 405174
rect 314786 404938 315022 405174
rect 314466 404618 314702 404854
rect 314786 404618 315022 404854
rect 314466 386938 314702 387174
rect 314786 386938 315022 387174
rect 314466 386618 314702 386854
rect 314786 386618 315022 386854
rect 314466 368938 314702 369174
rect 314786 368938 315022 369174
rect 314466 368618 314702 368854
rect 314786 368618 315022 368854
rect 314466 350938 314702 351174
rect 314786 350938 315022 351174
rect 314466 350618 314702 350854
rect 314786 350618 315022 350854
rect 314466 332938 314702 333174
rect 314786 332938 315022 333174
rect 314466 332618 314702 332854
rect 314786 332618 315022 332854
rect 314466 314938 314702 315174
rect 314786 314938 315022 315174
rect 314466 314618 314702 314854
rect 314786 314618 315022 314854
rect 314466 296938 314702 297174
rect 314786 296938 315022 297174
rect 314466 296618 314702 296854
rect 314786 296618 315022 296854
rect 314466 278938 314702 279174
rect 314786 278938 315022 279174
rect 314466 278618 314702 278854
rect 314786 278618 315022 278854
rect 314466 260938 314702 261174
rect 314786 260938 315022 261174
rect 314466 260618 314702 260854
rect 314786 260618 315022 260854
rect 314466 242938 314702 243174
rect 314786 242938 315022 243174
rect 314466 242618 314702 242854
rect 314786 242618 315022 242854
rect 314466 224938 314702 225174
rect 314786 224938 315022 225174
rect 314466 224618 314702 224854
rect 314786 224618 315022 224854
rect 314466 206938 314702 207174
rect 314786 206938 315022 207174
rect 314466 206618 314702 206854
rect 314786 206618 315022 206854
rect 314466 188938 314702 189174
rect 314786 188938 315022 189174
rect 314466 188618 314702 188854
rect 314786 188618 315022 188854
rect 314466 170938 314702 171174
rect 314786 170938 315022 171174
rect 314466 170618 314702 170854
rect 314786 170618 315022 170854
rect 314466 152938 314702 153174
rect 314786 152938 315022 153174
rect 314466 152618 314702 152854
rect 314786 152618 315022 152854
rect 314466 134938 314702 135174
rect 314786 134938 315022 135174
rect 314466 134618 314702 134854
rect 314786 134618 315022 134854
rect 314466 116938 314702 117174
rect 314786 116938 315022 117174
rect 314466 116618 314702 116854
rect 314786 116618 315022 116854
rect 314466 98938 314702 99174
rect 314786 98938 315022 99174
rect 314466 98618 314702 98854
rect 314786 98618 315022 98854
rect 314466 80938 314702 81174
rect 314786 80938 315022 81174
rect 314466 80618 314702 80854
rect 314786 80618 315022 80854
rect 314466 62938 314702 63174
rect 314786 62938 315022 63174
rect 314466 62618 314702 62854
rect 314786 62618 315022 62854
rect 314466 44938 314702 45174
rect 314786 44938 315022 45174
rect 314466 44618 314702 44854
rect 314786 44618 315022 44854
rect 314466 26938 314702 27174
rect 314786 26938 315022 27174
rect 314466 26618 314702 26854
rect 314786 26618 315022 26854
rect 314466 8938 314702 9174
rect 314786 8938 315022 9174
rect 314466 8618 314702 8854
rect 314786 8618 315022 8854
rect 314466 -2052 314702 -1816
rect 314786 -2052 315022 -1816
rect 314466 -2372 314702 -2136
rect 314786 -2372 315022 -2136
rect 318186 462776 318422 463012
rect 318506 462776 318742 463012
rect 318186 462456 318422 462692
rect 318506 462456 318742 462692
rect 318186 444658 318422 444894
rect 318506 444658 318742 444894
rect 318186 444338 318422 444574
rect 318506 444338 318742 444574
rect 318186 426658 318422 426894
rect 318506 426658 318742 426894
rect 318186 426338 318422 426574
rect 318506 426338 318742 426574
rect 318186 408658 318422 408894
rect 318506 408658 318742 408894
rect 318186 408338 318422 408574
rect 318506 408338 318742 408574
rect 318186 390658 318422 390894
rect 318506 390658 318742 390894
rect 318186 390338 318422 390574
rect 318506 390338 318742 390574
rect 318186 372658 318422 372894
rect 318506 372658 318742 372894
rect 318186 372338 318422 372574
rect 318506 372338 318742 372574
rect 318186 354658 318422 354894
rect 318506 354658 318742 354894
rect 318186 354338 318422 354574
rect 318506 354338 318742 354574
rect 318186 336658 318422 336894
rect 318506 336658 318742 336894
rect 318186 336338 318422 336574
rect 318506 336338 318742 336574
rect 318186 318658 318422 318894
rect 318506 318658 318742 318894
rect 318186 318338 318422 318574
rect 318506 318338 318742 318574
rect 318186 300658 318422 300894
rect 318506 300658 318742 300894
rect 318186 300338 318422 300574
rect 318506 300338 318742 300574
rect 318186 282658 318422 282894
rect 318506 282658 318742 282894
rect 318186 282338 318422 282574
rect 318506 282338 318742 282574
rect 318186 264658 318422 264894
rect 318506 264658 318742 264894
rect 318186 264338 318422 264574
rect 318506 264338 318742 264574
rect 318186 246658 318422 246894
rect 318506 246658 318742 246894
rect 318186 246338 318422 246574
rect 318506 246338 318742 246574
rect 318186 228658 318422 228894
rect 318506 228658 318742 228894
rect 318186 228338 318422 228574
rect 318506 228338 318742 228574
rect 318186 210658 318422 210894
rect 318506 210658 318742 210894
rect 318186 210338 318422 210574
rect 318506 210338 318742 210574
rect 318186 192658 318422 192894
rect 318506 192658 318742 192894
rect 318186 192338 318422 192574
rect 318506 192338 318742 192574
rect 318186 174658 318422 174894
rect 318506 174658 318742 174894
rect 318186 174338 318422 174574
rect 318506 174338 318742 174574
rect 318186 156658 318422 156894
rect 318506 156658 318742 156894
rect 318186 156338 318422 156574
rect 318506 156338 318742 156574
rect 318186 138658 318422 138894
rect 318506 138658 318742 138894
rect 318186 138338 318422 138574
rect 318506 138338 318742 138574
rect 318186 120658 318422 120894
rect 318506 120658 318742 120894
rect 318186 120338 318422 120574
rect 318506 120338 318742 120574
rect 318186 102658 318422 102894
rect 318506 102658 318742 102894
rect 318186 102338 318422 102574
rect 318506 102338 318742 102574
rect 318186 84658 318422 84894
rect 318506 84658 318742 84894
rect 318186 84338 318422 84574
rect 318506 84338 318742 84574
rect 318186 66658 318422 66894
rect 318506 66658 318742 66894
rect 318186 66338 318422 66574
rect 318506 66338 318742 66574
rect 318186 48658 318422 48894
rect 318506 48658 318742 48894
rect 318186 48338 318422 48574
rect 318506 48338 318742 48574
rect 318186 30658 318422 30894
rect 318506 30658 318742 30894
rect 318186 30338 318422 30574
rect 318506 30338 318742 30574
rect 318186 12658 318422 12894
rect 318506 12658 318742 12894
rect 318186 12338 318422 12574
rect 318506 12338 318742 12574
rect 318186 -3012 318422 -2776
rect 318506 -3012 318742 -2776
rect 318186 -3332 318422 -3096
rect 318506 -3332 318742 -3096
rect 321906 463736 322142 463972
rect 322226 463736 322462 463972
rect 321906 463416 322142 463652
rect 322226 463416 322462 463652
rect 321906 448378 322142 448614
rect 322226 448378 322462 448614
rect 321906 448058 322142 448294
rect 322226 448058 322462 448294
rect 321906 430378 322142 430614
rect 322226 430378 322462 430614
rect 321906 430058 322142 430294
rect 322226 430058 322462 430294
rect 321906 412378 322142 412614
rect 322226 412378 322462 412614
rect 321906 412058 322142 412294
rect 322226 412058 322462 412294
rect 321906 394378 322142 394614
rect 322226 394378 322462 394614
rect 321906 394058 322142 394294
rect 322226 394058 322462 394294
rect 321906 376378 322142 376614
rect 322226 376378 322462 376614
rect 321906 376058 322142 376294
rect 322226 376058 322462 376294
rect 321906 358378 322142 358614
rect 322226 358378 322462 358614
rect 321906 358058 322142 358294
rect 322226 358058 322462 358294
rect 321906 340378 322142 340614
rect 322226 340378 322462 340614
rect 321906 340058 322142 340294
rect 322226 340058 322462 340294
rect 321906 322378 322142 322614
rect 322226 322378 322462 322614
rect 321906 322058 322142 322294
rect 322226 322058 322462 322294
rect 321906 304378 322142 304614
rect 322226 304378 322462 304614
rect 321906 304058 322142 304294
rect 322226 304058 322462 304294
rect 321906 286378 322142 286614
rect 322226 286378 322462 286614
rect 321906 286058 322142 286294
rect 322226 286058 322462 286294
rect 321906 268378 322142 268614
rect 322226 268378 322462 268614
rect 321906 268058 322142 268294
rect 322226 268058 322462 268294
rect 321906 250378 322142 250614
rect 322226 250378 322462 250614
rect 321906 250058 322142 250294
rect 322226 250058 322462 250294
rect 321906 232378 322142 232614
rect 322226 232378 322462 232614
rect 321906 232058 322142 232294
rect 322226 232058 322462 232294
rect 321906 214378 322142 214614
rect 322226 214378 322462 214614
rect 321906 214058 322142 214294
rect 322226 214058 322462 214294
rect 321906 196378 322142 196614
rect 322226 196378 322462 196614
rect 321906 196058 322142 196294
rect 322226 196058 322462 196294
rect 321906 178378 322142 178614
rect 322226 178378 322462 178614
rect 321906 178058 322142 178294
rect 322226 178058 322462 178294
rect 321906 160378 322142 160614
rect 322226 160378 322462 160614
rect 321906 160058 322142 160294
rect 322226 160058 322462 160294
rect 321906 142378 322142 142614
rect 322226 142378 322462 142614
rect 321906 142058 322142 142294
rect 322226 142058 322462 142294
rect 321906 124378 322142 124614
rect 322226 124378 322462 124614
rect 321906 124058 322142 124294
rect 322226 124058 322462 124294
rect 321906 106378 322142 106614
rect 322226 106378 322462 106614
rect 321906 106058 322142 106294
rect 322226 106058 322462 106294
rect 321906 88378 322142 88614
rect 322226 88378 322462 88614
rect 321906 88058 322142 88294
rect 322226 88058 322462 88294
rect 321906 70378 322142 70614
rect 322226 70378 322462 70614
rect 321906 70058 322142 70294
rect 322226 70058 322462 70294
rect 321906 52378 322142 52614
rect 322226 52378 322462 52614
rect 321906 52058 322142 52294
rect 322226 52058 322462 52294
rect 321906 34378 322142 34614
rect 322226 34378 322462 34614
rect 321906 34058 322142 34294
rect 322226 34058 322462 34294
rect 321906 16378 322142 16614
rect 322226 16378 322462 16614
rect 321906 16058 322142 16294
rect 322226 16058 322462 16294
rect 321906 -3972 322142 -3736
rect 322226 -3972 322462 -3736
rect 321906 -4292 322142 -4056
rect 322226 -4292 322462 -4056
rect 328746 460856 328982 461092
rect 329066 460856 329302 461092
rect 328746 460536 328982 460772
rect 329066 460536 329302 460772
rect 354186 462776 354422 463012
rect 354506 462776 354742 463012
rect 354186 462456 354422 462692
rect 354506 462456 354742 462692
rect 328746 455218 328982 455454
rect 329066 455218 329302 455454
rect 328746 454898 328982 455134
rect 329066 454898 329302 455134
rect 328746 437218 328982 437454
rect 329066 437218 329302 437454
rect 328746 436898 328982 437134
rect 329066 436898 329302 437134
rect 328746 419218 328982 419454
rect 329066 419218 329302 419454
rect 328746 418898 328982 419134
rect 329066 418898 329302 419134
rect 328746 401218 328982 401454
rect 329066 401218 329302 401454
rect 328746 400898 328982 401134
rect 329066 400898 329302 401134
rect 328746 383218 328982 383454
rect 329066 383218 329302 383454
rect 328746 382898 328982 383134
rect 329066 382898 329302 383134
rect 328746 365218 328982 365454
rect 329066 365218 329302 365454
rect 328746 364898 328982 365134
rect 329066 364898 329302 365134
rect 328746 347218 328982 347454
rect 329066 347218 329302 347454
rect 328746 346898 328982 347134
rect 329066 346898 329302 347134
rect 328746 329218 328982 329454
rect 329066 329218 329302 329454
rect 328746 328898 328982 329134
rect 329066 328898 329302 329134
rect 328746 311218 328982 311454
rect 329066 311218 329302 311454
rect 328746 310898 328982 311134
rect 329066 310898 329302 311134
rect 328746 293218 328982 293454
rect 329066 293218 329302 293454
rect 328746 292898 328982 293134
rect 329066 292898 329302 293134
rect 328746 275218 328982 275454
rect 329066 275218 329302 275454
rect 328746 274898 328982 275134
rect 329066 274898 329302 275134
rect 328746 257218 328982 257454
rect 329066 257218 329302 257454
rect 328746 256898 328982 257134
rect 329066 256898 329302 257134
rect 328746 239218 328982 239454
rect 329066 239218 329302 239454
rect 328746 238898 328982 239134
rect 329066 238898 329302 239134
rect 328746 221218 328982 221454
rect 329066 221218 329302 221454
rect 328746 220898 328982 221134
rect 329066 220898 329302 221134
rect 328746 203218 328982 203454
rect 329066 203218 329302 203454
rect 328746 202898 328982 203134
rect 329066 202898 329302 203134
rect 328746 185218 328982 185454
rect 329066 185218 329302 185454
rect 328746 184898 328982 185134
rect 329066 184898 329302 185134
rect 328746 167218 328982 167454
rect 329066 167218 329302 167454
rect 328746 166898 328982 167134
rect 329066 166898 329302 167134
rect 328746 149218 328982 149454
rect 329066 149218 329302 149454
rect 328746 148898 328982 149134
rect 329066 148898 329302 149134
rect 328746 131218 328982 131454
rect 329066 131218 329302 131454
rect 328746 130898 328982 131134
rect 329066 130898 329302 131134
rect 328746 113218 328982 113454
rect 329066 113218 329302 113454
rect 328746 112898 328982 113134
rect 329066 112898 329302 113134
rect 328746 95218 328982 95454
rect 329066 95218 329302 95454
rect 328746 94898 328982 95134
rect 329066 94898 329302 95134
rect 328746 77218 328982 77454
rect 329066 77218 329302 77454
rect 328746 76898 328982 77134
rect 329066 76898 329302 77134
rect 328746 59218 328982 59454
rect 329066 59218 329302 59454
rect 328746 58898 328982 59134
rect 329066 58898 329302 59134
rect 328746 41218 328982 41454
rect 329066 41218 329302 41454
rect 328746 40898 328982 41134
rect 329066 40898 329302 41134
rect 328746 23218 328982 23454
rect 329066 23218 329302 23454
rect 328746 22898 328982 23134
rect 329066 22898 329302 23134
rect 328746 5218 328982 5454
rect 329066 5218 329302 5454
rect 328746 4898 328982 5134
rect 329066 4898 329302 5134
rect 328746 -1092 328982 -856
rect 329066 -1092 329302 -856
rect 328746 -1412 328982 -1176
rect 329066 -1412 329302 -1176
rect 332466 440938 332702 441174
rect 332786 440938 333022 441174
rect 332466 440618 332702 440854
rect 332786 440618 333022 440854
rect 332466 422938 332702 423174
rect 332786 422938 333022 423174
rect 332466 422618 332702 422854
rect 332786 422618 333022 422854
rect 332466 404938 332702 405174
rect 332786 404938 333022 405174
rect 332466 404618 332702 404854
rect 332786 404618 333022 404854
rect 332466 386938 332702 387174
rect 332786 386938 333022 387174
rect 332466 386618 332702 386854
rect 332786 386618 333022 386854
rect 332466 368938 332702 369174
rect 332786 368938 333022 369174
rect 332466 368618 332702 368854
rect 332786 368618 333022 368854
rect 332466 350938 332702 351174
rect 332786 350938 333022 351174
rect 332466 350618 332702 350854
rect 332786 350618 333022 350854
rect 332466 332938 332702 333174
rect 332786 332938 333022 333174
rect 332466 332618 332702 332854
rect 332786 332618 333022 332854
rect 332466 314938 332702 315174
rect 332786 314938 333022 315174
rect 332466 314618 332702 314854
rect 332786 314618 333022 314854
rect 332466 296938 332702 297174
rect 332786 296938 333022 297174
rect 332466 296618 332702 296854
rect 332786 296618 333022 296854
rect 332466 278938 332702 279174
rect 332786 278938 333022 279174
rect 332466 278618 332702 278854
rect 332786 278618 333022 278854
rect 332466 260938 332702 261174
rect 332786 260938 333022 261174
rect 332466 260618 332702 260854
rect 332786 260618 333022 260854
rect 332466 242938 332702 243174
rect 332786 242938 333022 243174
rect 332466 242618 332702 242854
rect 332786 242618 333022 242854
rect 332466 224938 332702 225174
rect 332786 224938 333022 225174
rect 332466 224618 332702 224854
rect 332786 224618 333022 224854
rect 332466 206938 332702 207174
rect 332786 206938 333022 207174
rect 332466 206618 332702 206854
rect 332786 206618 333022 206854
rect 332466 188938 332702 189174
rect 332786 188938 333022 189174
rect 332466 188618 332702 188854
rect 332786 188618 333022 188854
rect 332466 170938 332702 171174
rect 332786 170938 333022 171174
rect 332466 170618 332702 170854
rect 332786 170618 333022 170854
rect 332466 152938 332702 153174
rect 332786 152938 333022 153174
rect 332466 152618 332702 152854
rect 332786 152618 333022 152854
rect 332466 134938 332702 135174
rect 332786 134938 333022 135174
rect 332466 134618 332702 134854
rect 332786 134618 333022 134854
rect 332466 116938 332702 117174
rect 332786 116938 333022 117174
rect 332466 116618 332702 116854
rect 332786 116618 333022 116854
rect 332466 98938 332702 99174
rect 332786 98938 333022 99174
rect 332466 98618 332702 98854
rect 332786 98618 333022 98854
rect 332466 80938 332702 81174
rect 332786 80938 333022 81174
rect 332466 80618 332702 80854
rect 332786 80618 333022 80854
rect 332466 62938 332702 63174
rect 332786 62938 333022 63174
rect 332466 62618 332702 62854
rect 332786 62618 333022 62854
rect 332466 44938 332702 45174
rect 332786 44938 333022 45174
rect 332466 44618 332702 44854
rect 332786 44618 333022 44854
rect 332466 26938 332702 27174
rect 332786 26938 333022 27174
rect 332466 26618 332702 26854
rect 332786 26618 333022 26854
rect 332466 8938 332702 9174
rect 332786 8938 333022 9174
rect 332466 8618 332702 8854
rect 332786 8618 333022 8854
rect 332466 -2052 332702 -1816
rect 332786 -2052 333022 -1816
rect 332466 -2372 332702 -2136
rect 332786 -2372 333022 -2136
rect 336186 444658 336422 444894
rect 336506 444658 336742 444894
rect 336186 444338 336422 444574
rect 336506 444338 336742 444574
rect 336186 426658 336422 426894
rect 336506 426658 336742 426894
rect 336186 426338 336422 426574
rect 336506 426338 336742 426574
rect 336186 408658 336422 408894
rect 336506 408658 336742 408894
rect 336186 408338 336422 408574
rect 336506 408338 336742 408574
rect 336186 390658 336422 390894
rect 336506 390658 336742 390894
rect 336186 390338 336422 390574
rect 336506 390338 336742 390574
rect 336186 372658 336422 372894
rect 336506 372658 336742 372894
rect 336186 372338 336422 372574
rect 336506 372338 336742 372574
rect 336186 354658 336422 354894
rect 336506 354658 336742 354894
rect 336186 354338 336422 354574
rect 336506 354338 336742 354574
rect 336186 336658 336422 336894
rect 336506 336658 336742 336894
rect 336186 336338 336422 336574
rect 336506 336338 336742 336574
rect 336186 318658 336422 318894
rect 336506 318658 336742 318894
rect 336186 318338 336422 318574
rect 336506 318338 336742 318574
rect 336186 300658 336422 300894
rect 336506 300658 336742 300894
rect 336186 300338 336422 300574
rect 336506 300338 336742 300574
rect 336186 282658 336422 282894
rect 336506 282658 336742 282894
rect 336186 282338 336422 282574
rect 336506 282338 336742 282574
rect 336186 264658 336422 264894
rect 336506 264658 336742 264894
rect 336186 264338 336422 264574
rect 336506 264338 336742 264574
rect 336186 246658 336422 246894
rect 336506 246658 336742 246894
rect 336186 246338 336422 246574
rect 336506 246338 336742 246574
rect 336186 228658 336422 228894
rect 336506 228658 336742 228894
rect 336186 228338 336422 228574
rect 336506 228338 336742 228574
rect 336186 210658 336422 210894
rect 336506 210658 336742 210894
rect 336186 210338 336422 210574
rect 336506 210338 336742 210574
rect 336186 192658 336422 192894
rect 336506 192658 336742 192894
rect 336186 192338 336422 192574
rect 336506 192338 336742 192574
rect 336186 174658 336422 174894
rect 336506 174658 336742 174894
rect 336186 174338 336422 174574
rect 336506 174338 336742 174574
rect 336186 156658 336422 156894
rect 336506 156658 336742 156894
rect 336186 156338 336422 156574
rect 336506 156338 336742 156574
rect 336186 138658 336422 138894
rect 336506 138658 336742 138894
rect 336186 138338 336422 138574
rect 336506 138338 336742 138574
rect 336186 120658 336422 120894
rect 336506 120658 336742 120894
rect 336186 120338 336422 120574
rect 336506 120338 336742 120574
rect 336186 102658 336422 102894
rect 336506 102658 336742 102894
rect 336186 102338 336422 102574
rect 336506 102338 336742 102574
rect 336186 84658 336422 84894
rect 336506 84658 336742 84894
rect 336186 84338 336422 84574
rect 336506 84338 336742 84574
rect 336186 66658 336422 66894
rect 336506 66658 336742 66894
rect 336186 66338 336422 66574
rect 336506 66338 336742 66574
rect 336186 48658 336422 48894
rect 336506 48658 336742 48894
rect 336186 48338 336422 48574
rect 336506 48338 336742 48574
rect 336186 30658 336422 30894
rect 336506 30658 336742 30894
rect 336186 30338 336422 30574
rect 336506 30338 336742 30574
rect 336186 12658 336422 12894
rect 336506 12658 336742 12894
rect 336186 12338 336422 12574
rect 336506 12338 336742 12574
rect 336186 -3012 336422 -2776
rect 336506 -3012 336742 -2776
rect 336186 -3332 336422 -3096
rect 336506 -3332 336742 -3096
rect 339906 448378 340142 448614
rect 340226 448378 340462 448614
rect 339906 448058 340142 448294
rect 340226 448058 340462 448294
rect 339906 430378 340142 430614
rect 340226 430378 340462 430614
rect 339906 430058 340142 430294
rect 340226 430058 340462 430294
rect 339906 412378 340142 412614
rect 340226 412378 340462 412614
rect 339906 412058 340142 412294
rect 340226 412058 340462 412294
rect 339906 394378 340142 394614
rect 340226 394378 340462 394614
rect 339906 394058 340142 394294
rect 340226 394058 340462 394294
rect 339906 376378 340142 376614
rect 340226 376378 340462 376614
rect 339906 376058 340142 376294
rect 340226 376058 340462 376294
rect 339906 358378 340142 358614
rect 340226 358378 340462 358614
rect 339906 358058 340142 358294
rect 340226 358058 340462 358294
rect 339906 340378 340142 340614
rect 340226 340378 340462 340614
rect 339906 340058 340142 340294
rect 340226 340058 340462 340294
rect 339906 322378 340142 322614
rect 340226 322378 340462 322614
rect 339906 322058 340142 322294
rect 340226 322058 340462 322294
rect 339906 304378 340142 304614
rect 340226 304378 340462 304614
rect 339906 304058 340142 304294
rect 340226 304058 340462 304294
rect 339906 286378 340142 286614
rect 340226 286378 340462 286614
rect 339906 286058 340142 286294
rect 340226 286058 340462 286294
rect 339906 268378 340142 268614
rect 340226 268378 340462 268614
rect 339906 268058 340142 268294
rect 340226 268058 340462 268294
rect 339906 250378 340142 250614
rect 340226 250378 340462 250614
rect 339906 250058 340142 250294
rect 340226 250058 340462 250294
rect 339906 232378 340142 232614
rect 340226 232378 340462 232614
rect 339906 232058 340142 232294
rect 340226 232058 340462 232294
rect 339906 214378 340142 214614
rect 340226 214378 340462 214614
rect 339906 214058 340142 214294
rect 340226 214058 340462 214294
rect 339906 196378 340142 196614
rect 340226 196378 340462 196614
rect 339906 196058 340142 196294
rect 340226 196058 340462 196294
rect 339906 178378 340142 178614
rect 340226 178378 340462 178614
rect 339906 178058 340142 178294
rect 340226 178058 340462 178294
rect 339906 160378 340142 160614
rect 340226 160378 340462 160614
rect 339906 160058 340142 160294
rect 340226 160058 340462 160294
rect 339906 142378 340142 142614
rect 340226 142378 340462 142614
rect 339906 142058 340142 142294
rect 340226 142058 340462 142294
rect 339906 124378 340142 124614
rect 340226 124378 340462 124614
rect 339906 124058 340142 124294
rect 340226 124058 340462 124294
rect 339906 106378 340142 106614
rect 340226 106378 340462 106614
rect 339906 106058 340142 106294
rect 340226 106058 340462 106294
rect 339906 88378 340142 88614
rect 340226 88378 340462 88614
rect 339906 88058 340142 88294
rect 340226 88058 340462 88294
rect 339906 70378 340142 70614
rect 340226 70378 340462 70614
rect 339906 70058 340142 70294
rect 340226 70058 340462 70294
rect 339906 52378 340142 52614
rect 340226 52378 340462 52614
rect 339906 52058 340142 52294
rect 340226 52058 340462 52294
rect 339906 34378 340142 34614
rect 340226 34378 340462 34614
rect 339906 34058 340142 34294
rect 340226 34058 340462 34294
rect 339906 16378 340142 16614
rect 340226 16378 340462 16614
rect 339906 16058 340142 16294
rect 340226 16058 340462 16294
rect 339906 -3972 340142 -3736
rect 340226 -3972 340462 -3736
rect 339906 -4292 340142 -4056
rect 340226 -4292 340462 -4056
rect 346746 455218 346982 455454
rect 347066 455218 347302 455454
rect 346746 454898 346982 455134
rect 347066 454898 347302 455134
rect 346746 437218 346982 437454
rect 347066 437218 347302 437454
rect 346746 436898 346982 437134
rect 347066 436898 347302 437134
rect 346746 419218 346982 419454
rect 347066 419218 347302 419454
rect 346746 418898 346982 419134
rect 347066 418898 347302 419134
rect 346746 401218 346982 401454
rect 347066 401218 347302 401454
rect 346746 400898 346982 401134
rect 347066 400898 347302 401134
rect 346746 383218 346982 383454
rect 347066 383218 347302 383454
rect 346746 382898 346982 383134
rect 347066 382898 347302 383134
rect 346746 365218 346982 365454
rect 347066 365218 347302 365454
rect 346746 364898 346982 365134
rect 347066 364898 347302 365134
rect 346746 347218 346982 347454
rect 347066 347218 347302 347454
rect 346746 346898 346982 347134
rect 347066 346898 347302 347134
rect 346746 329218 346982 329454
rect 347066 329218 347302 329454
rect 346746 328898 346982 329134
rect 347066 328898 347302 329134
rect 346746 311218 346982 311454
rect 347066 311218 347302 311454
rect 346746 310898 346982 311134
rect 347066 310898 347302 311134
rect 346746 293218 346982 293454
rect 347066 293218 347302 293454
rect 346746 292898 346982 293134
rect 347066 292898 347302 293134
rect 346746 275218 346982 275454
rect 347066 275218 347302 275454
rect 346746 274898 346982 275134
rect 347066 274898 347302 275134
rect 346746 257218 346982 257454
rect 347066 257218 347302 257454
rect 346746 256898 346982 257134
rect 347066 256898 347302 257134
rect 346746 239218 346982 239454
rect 347066 239218 347302 239454
rect 346746 238898 346982 239134
rect 347066 238898 347302 239134
rect 346746 221218 346982 221454
rect 347066 221218 347302 221454
rect 346746 220898 346982 221134
rect 347066 220898 347302 221134
rect 346746 203218 346982 203454
rect 347066 203218 347302 203454
rect 346746 202898 346982 203134
rect 347066 202898 347302 203134
rect 346746 185218 346982 185454
rect 347066 185218 347302 185454
rect 346746 184898 346982 185134
rect 347066 184898 347302 185134
rect 346746 167218 346982 167454
rect 347066 167218 347302 167454
rect 346746 166898 346982 167134
rect 347066 166898 347302 167134
rect 346746 149218 346982 149454
rect 347066 149218 347302 149454
rect 346746 148898 346982 149134
rect 347066 148898 347302 149134
rect 346746 131218 346982 131454
rect 347066 131218 347302 131454
rect 346746 130898 346982 131134
rect 347066 130898 347302 131134
rect 346746 113218 346982 113454
rect 347066 113218 347302 113454
rect 346746 112898 346982 113134
rect 347066 112898 347302 113134
rect 346746 95218 346982 95454
rect 347066 95218 347302 95454
rect 346746 94898 346982 95134
rect 347066 94898 347302 95134
rect 346746 77218 346982 77454
rect 347066 77218 347302 77454
rect 346746 76898 346982 77134
rect 347066 76898 347302 77134
rect 346746 59218 346982 59454
rect 347066 59218 347302 59454
rect 346746 58898 346982 59134
rect 347066 58898 347302 59134
rect 346746 41218 346982 41454
rect 347066 41218 347302 41454
rect 346746 40898 346982 41134
rect 347066 40898 347302 41134
rect 346746 23218 346982 23454
rect 347066 23218 347302 23454
rect 346746 22898 346982 23134
rect 347066 22898 347302 23134
rect 346746 5218 346982 5454
rect 347066 5218 347302 5454
rect 346746 4898 346982 5134
rect 347066 4898 347302 5134
rect 346746 -1092 346982 -856
rect 347066 -1092 347302 -856
rect 346746 -1412 346982 -1176
rect 347066 -1412 347302 -1176
rect 350466 440938 350702 441174
rect 350786 440938 351022 441174
rect 350466 440618 350702 440854
rect 350786 440618 351022 440854
rect 350466 422938 350702 423174
rect 350786 422938 351022 423174
rect 350466 422618 350702 422854
rect 350786 422618 351022 422854
rect 350466 404938 350702 405174
rect 350786 404938 351022 405174
rect 350466 404618 350702 404854
rect 350786 404618 351022 404854
rect 350466 386938 350702 387174
rect 350786 386938 351022 387174
rect 350466 386618 350702 386854
rect 350786 386618 351022 386854
rect 350466 368938 350702 369174
rect 350786 368938 351022 369174
rect 350466 368618 350702 368854
rect 350786 368618 351022 368854
rect 350466 350938 350702 351174
rect 350786 350938 351022 351174
rect 350466 350618 350702 350854
rect 350786 350618 351022 350854
rect 350466 332938 350702 333174
rect 350786 332938 351022 333174
rect 350466 332618 350702 332854
rect 350786 332618 351022 332854
rect 350466 314938 350702 315174
rect 350786 314938 351022 315174
rect 350466 314618 350702 314854
rect 350786 314618 351022 314854
rect 350466 296938 350702 297174
rect 350786 296938 351022 297174
rect 350466 296618 350702 296854
rect 350786 296618 351022 296854
rect 350466 278938 350702 279174
rect 350786 278938 351022 279174
rect 350466 278618 350702 278854
rect 350786 278618 351022 278854
rect 350466 260938 350702 261174
rect 350786 260938 351022 261174
rect 350466 260618 350702 260854
rect 350786 260618 351022 260854
rect 350466 242938 350702 243174
rect 350786 242938 351022 243174
rect 350466 242618 350702 242854
rect 350786 242618 351022 242854
rect 350466 224938 350702 225174
rect 350786 224938 351022 225174
rect 350466 224618 350702 224854
rect 350786 224618 351022 224854
rect 350466 206938 350702 207174
rect 350786 206938 351022 207174
rect 350466 206618 350702 206854
rect 350786 206618 351022 206854
rect 350466 188938 350702 189174
rect 350786 188938 351022 189174
rect 350466 188618 350702 188854
rect 350786 188618 351022 188854
rect 350466 170938 350702 171174
rect 350786 170938 351022 171174
rect 350466 170618 350702 170854
rect 350786 170618 351022 170854
rect 350466 152938 350702 153174
rect 350786 152938 351022 153174
rect 350466 152618 350702 152854
rect 350786 152618 351022 152854
rect 350466 134938 350702 135174
rect 350786 134938 351022 135174
rect 350466 134618 350702 134854
rect 350786 134618 351022 134854
rect 350466 116938 350702 117174
rect 350786 116938 351022 117174
rect 350466 116618 350702 116854
rect 350786 116618 351022 116854
rect 350466 98938 350702 99174
rect 350786 98938 351022 99174
rect 350466 98618 350702 98854
rect 350786 98618 351022 98854
rect 350466 80938 350702 81174
rect 350786 80938 351022 81174
rect 350466 80618 350702 80854
rect 350786 80618 351022 80854
rect 350466 62938 350702 63174
rect 350786 62938 351022 63174
rect 350466 62618 350702 62854
rect 350786 62618 351022 62854
rect 350466 44938 350702 45174
rect 350786 44938 351022 45174
rect 350466 44618 350702 44854
rect 350786 44618 351022 44854
rect 350466 26938 350702 27174
rect 350786 26938 351022 27174
rect 350466 26618 350702 26854
rect 350786 26618 351022 26854
rect 350466 8938 350702 9174
rect 350786 8938 351022 9174
rect 350466 8618 350702 8854
rect 350786 8618 351022 8854
rect 350466 -2052 350702 -1816
rect 350786 -2052 351022 -1816
rect 350466 -2372 350702 -2136
rect 350786 -2372 351022 -2136
rect 354186 444658 354422 444894
rect 354506 444658 354742 444894
rect 354186 444338 354422 444574
rect 354506 444338 354742 444574
rect 354186 426658 354422 426894
rect 354506 426658 354742 426894
rect 354186 426338 354422 426574
rect 354506 426338 354742 426574
rect 354186 408658 354422 408894
rect 354506 408658 354742 408894
rect 354186 408338 354422 408574
rect 354506 408338 354742 408574
rect 354186 390658 354422 390894
rect 354506 390658 354742 390894
rect 354186 390338 354422 390574
rect 354506 390338 354742 390574
rect 354186 372658 354422 372894
rect 354506 372658 354742 372894
rect 354186 372338 354422 372574
rect 354506 372338 354742 372574
rect 354186 354658 354422 354894
rect 354506 354658 354742 354894
rect 354186 354338 354422 354574
rect 354506 354338 354742 354574
rect 354186 336658 354422 336894
rect 354506 336658 354742 336894
rect 354186 336338 354422 336574
rect 354506 336338 354742 336574
rect 354186 318658 354422 318894
rect 354506 318658 354742 318894
rect 354186 318338 354422 318574
rect 354506 318338 354742 318574
rect 354186 300658 354422 300894
rect 354506 300658 354742 300894
rect 354186 300338 354422 300574
rect 354506 300338 354742 300574
rect 354186 282658 354422 282894
rect 354506 282658 354742 282894
rect 354186 282338 354422 282574
rect 354506 282338 354742 282574
rect 354186 264658 354422 264894
rect 354506 264658 354742 264894
rect 354186 264338 354422 264574
rect 354506 264338 354742 264574
rect 354186 246658 354422 246894
rect 354506 246658 354742 246894
rect 354186 246338 354422 246574
rect 354506 246338 354742 246574
rect 354186 228658 354422 228894
rect 354506 228658 354742 228894
rect 354186 228338 354422 228574
rect 354506 228338 354742 228574
rect 354186 210658 354422 210894
rect 354506 210658 354742 210894
rect 354186 210338 354422 210574
rect 354506 210338 354742 210574
rect 354186 192658 354422 192894
rect 354506 192658 354742 192894
rect 354186 192338 354422 192574
rect 354506 192338 354742 192574
rect 354186 174658 354422 174894
rect 354506 174658 354742 174894
rect 354186 174338 354422 174574
rect 354506 174338 354742 174574
rect 354186 156658 354422 156894
rect 354506 156658 354742 156894
rect 354186 156338 354422 156574
rect 354506 156338 354742 156574
rect 354186 138658 354422 138894
rect 354506 138658 354742 138894
rect 354186 138338 354422 138574
rect 354506 138338 354742 138574
rect 354186 120658 354422 120894
rect 354506 120658 354742 120894
rect 354186 120338 354422 120574
rect 354506 120338 354742 120574
rect 354186 102658 354422 102894
rect 354506 102658 354742 102894
rect 354186 102338 354422 102574
rect 354506 102338 354742 102574
rect 354186 84658 354422 84894
rect 354506 84658 354742 84894
rect 354186 84338 354422 84574
rect 354506 84338 354742 84574
rect 354186 66658 354422 66894
rect 354506 66658 354742 66894
rect 354186 66338 354422 66574
rect 354506 66338 354742 66574
rect 354186 48658 354422 48894
rect 354506 48658 354742 48894
rect 354186 48338 354422 48574
rect 354506 48338 354742 48574
rect 354186 30658 354422 30894
rect 354506 30658 354742 30894
rect 354186 30338 354422 30574
rect 354506 30338 354742 30574
rect 354186 12658 354422 12894
rect 354506 12658 354742 12894
rect 354186 12338 354422 12574
rect 354506 12338 354742 12574
rect 354186 -3012 354422 -2776
rect 354506 -3012 354742 -2776
rect 354186 -3332 354422 -3096
rect 354506 -3332 354742 -3096
rect 357906 463736 358142 463972
rect 358226 463736 358462 463972
rect 357906 463416 358142 463652
rect 358226 463416 358462 463652
rect 357906 448378 358142 448614
rect 358226 448378 358462 448614
rect 357906 448058 358142 448294
rect 358226 448058 358462 448294
rect 357906 430378 358142 430614
rect 358226 430378 358462 430614
rect 357906 430058 358142 430294
rect 358226 430058 358462 430294
rect 357906 412378 358142 412614
rect 358226 412378 358462 412614
rect 357906 412058 358142 412294
rect 358226 412058 358462 412294
rect 357906 394378 358142 394614
rect 358226 394378 358462 394614
rect 357906 394058 358142 394294
rect 358226 394058 358462 394294
rect 357906 376378 358142 376614
rect 358226 376378 358462 376614
rect 357906 376058 358142 376294
rect 358226 376058 358462 376294
rect 357906 358378 358142 358614
rect 358226 358378 358462 358614
rect 357906 358058 358142 358294
rect 358226 358058 358462 358294
rect 357906 340378 358142 340614
rect 358226 340378 358462 340614
rect 357906 340058 358142 340294
rect 358226 340058 358462 340294
rect 357906 322378 358142 322614
rect 358226 322378 358462 322614
rect 357906 322058 358142 322294
rect 358226 322058 358462 322294
rect 357906 304378 358142 304614
rect 358226 304378 358462 304614
rect 357906 304058 358142 304294
rect 358226 304058 358462 304294
rect 357906 286378 358142 286614
rect 358226 286378 358462 286614
rect 357906 286058 358142 286294
rect 358226 286058 358462 286294
rect 357906 268378 358142 268614
rect 358226 268378 358462 268614
rect 357906 268058 358142 268294
rect 358226 268058 358462 268294
rect 357906 250378 358142 250614
rect 358226 250378 358462 250614
rect 357906 250058 358142 250294
rect 358226 250058 358462 250294
rect 357906 232378 358142 232614
rect 358226 232378 358462 232614
rect 357906 232058 358142 232294
rect 358226 232058 358462 232294
rect 357906 214378 358142 214614
rect 358226 214378 358462 214614
rect 357906 214058 358142 214294
rect 358226 214058 358462 214294
rect 357906 196378 358142 196614
rect 358226 196378 358462 196614
rect 357906 196058 358142 196294
rect 358226 196058 358462 196294
rect 357906 178378 358142 178614
rect 358226 178378 358462 178614
rect 357906 178058 358142 178294
rect 358226 178058 358462 178294
rect 357906 160378 358142 160614
rect 358226 160378 358462 160614
rect 357906 160058 358142 160294
rect 358226 160058 358462 160294
rect 357906 142378 358142 142614
rect 358226 142378 358462 142614
rect 357906 142058 358142 142294
rect 358226 142058 358462 142294
rect 357906 124378 358142 124614
rect 358226 124378 358462 124614
rect 357906 124058 358142 124294
rect 358226 124058 358462 124294
rect 357906 106378 358142 106614
rect 358226 106378 358462 106614
rect 357906 106058 358142 106294
rect 358226 106058 358462 106294
rect 357906 88378 358142 88614
rect 358226 88378 358462 88614
rect 357906 88058 358142 88294
rect 358226 88058 358462 88294
rect 357906 70378 358142 70614
rect 358226 70378 358462 70614
rect 357906 70058 358142 70294
rect 358226 70058 358462 70294
rect 357906 52378 358142 52614
rect 358226 52378 358462 52614
rect 357906 52058 358142 52294
rect 358226 52058 358462 52294
rect 357906 34378 358142 34614
rect 358226 34378 358462 34614
rect 357906 34058 358142 34294
rect 358226 34058 358462 34294
rect 357906 16378 358142 16614
rect 358226 16378 358462 16614
rect 357906 16058 358142 16294
rect 358226 16058 358462 16294
rect 357906 -3972 358142 -3736
rect 358226 -3972 358462 -3736
rect 357906 -4292 358142 -4056
rect 358226 -4292 358462 -4056
rect 364746 460856 364982 461092
rect 365066 460856 365302 461092
rect 364746 460536 364982 460772
rect 365066 460536 365302 460772
rect 364746 455218 364982 455454
rect 365066 455218 365302 455454
rect 364746 454898 364982 455134
rect 365066 454898 365302 455134
rect 364746 437218 364982 437454
rect 365066 437218 365302 437454
rect 364746 436898 364982 437134
rect 365066 436898 365302 437134
rect 364746 419218 364982 419454
rect 365066 419218 365302 419454
rect 364746 418898 364982 419134
rect 365066 418898 365302 419134
rect 364746 401218 364982 401454
rect 365066 401218 365302 401454
rect 364746 400898 364982 401134
rect 365066 400898 365302 401134
rect 364746 383218 364982 383454
rect 365066 383218 365302 383454
rect 364746 382898 364982 383134
rect 365066 382898 365302 383134
rect 364746 365218 364982 365454
rect 365066 365218 365302 365454
rect 364746 364898 364982 365134
rect 365066 364898 365302 365134
rect 364746 347218 364982 347454
rect 365066 347218 365302 347454
rect 364746 346898 364982 347134
rect 365066 346898 365302 347134
rect 364746 329218 364982 329454
rect 365066 329218 365302 329454
rect 364746 328898 364982 329134
rect 365066 328898 365302 329134
rect 364746 311218 364982 311454
rect 365066 311218 365302 311454
rect 364746 310898 364982 311134
rect 365066 310898 365302 311134
rect 364746 293218 364982 293454
rect 365066 293218 365302 293454
rect 364746 292898 364982 293134
rect 365066 292898 365302 293134
rect 364746 275218 364982 275454
rect 365066 275218 365302 275454
rect 364746 274898 364982 275134
rect 365066 274898 365302 275134
rect 364746 257218 364982 257454
rect 365066 257218 365302 257454
rect 364746 256898 364982 257134
rect 365066 256898 365302 257134
rect 364746 239218 364982 239454
rect 365066 239218 365302 239454
rect 364746 238898 364982 239134
rect 365066 238898 365302 239134
rect 364746 221218 364982 221454
rect 365066 221218 365302 221454
rect 364746 220898 364982 221134
rect 365066 220898 365302 221134
rect 364746 203218 364982 203454
rect 365066 203218 365302 203454
rect 364746 202898 364982 203134
rect 365066 202898 365302 203134
rect 364746 185218 364982 185454
rect 365066 185218 365302 185454
rect 364746 184898 364982 185134
rect 365066 184898 365302 185134
rect 364746 167218 364982 167454
rect 365066 167218 365302 167454
rect 364746 166898 364982 167134
rect 365066 166898 365302 167134
rect 364746 149218 364982 149454
rect 365066 149218 365302 149454
rect 364746 148898 364982 149134
rect 365066 148898 365302 149134
rect 364746 131218 364982 131454
rect 365066 131218 365302 131454
rect 364746 130898 364982 131134
rect 365066 130898 365302 131134
rect 364746 113218 364982 113454
rect 365066 113218 365302 113454
rect 364746 112898 364982 113134
rect 365066 112898 365302 113134
rect 364746 95218 364982 95454
rect 365066 95218 365302 95454
rect 364746 94898 364982 95134
rect 365066 94898 365302 95134
rect 364746 77218 364982 77454
rect 365066 77218 365302 77454
rect 364746 76898 364982 77134
rect 365066 76898 365302 77134
rect 364746 59218 364982 59454
rect 365066 59218 365302 59454
rect 364746 58898 364982 59134
rect 365066 58898 365302 59134
rect 364746 41218 364982 41454
rect 365066 41218 365302 41454
rect 364746 40898 364982 41134
rect 365066 40898 365302 41134
rect 364746 23218 364982 23454
rect 365066 23218 365302 23454
rect 364746 22898 364982 23134
rect 365066 22898 365302 23134
rect 364746 5218 364982 5454
rect 365066 5218 365302 5454
rect 364746 4898 364982 5134
rect 365066 4898 365302 5134
rect 364746 -1092 364982 -856
rect 365066 -1092 365302 -856
rect 364746 -1412 364982 -1176
rect 365066 -1412 365302 -1176
rect 368466 461816 368702 462052
rect 368786 461816 369022 462052
rect 368466 461496 368702 461732
rect 368786 461496 369022 461732
rect 368466 440938 368702 441174
rect 368786 440938 369022 441174
rect 368466 440618 368702 440854
rect 368786 440618 369022 440854
rect 368466 422938 368702 423174
rect 368786 422938 369022 423174
rect 368466 422618 368702 422854
rect 368786 422618 369022 422854
rect 368466 404938 368702 405174
rect 368786 404938 369022 405174
rect 368466 404618 368702 404854
rect 368786 404618 369022 404854
rect 368466 386938 368702 387174
rect 368786 386938 369022 387174
rect 368466 386618 368702 386854
rect 368786 386618 369022 386854
rect 368466 368938 368702 369174
rect 368786 368938 369022 369174
rect 368466 368618 368702 368854
rect 368786 368618 369022 368854
rect 368466 350938 368702 351174
rect 368786 350938 369022 351174
rect 368466 350618 368702 350854
rect 368786 350618 369022 350854
rect 368466 332938 368702 333174
rect 368786 332938 369022 333174
rect 368466 332618 368702 332854
rect 368786 332618 369022 332854
rect 368466 314938 368702 315174
rect 368786 314938 369022 315174
rect 368466 314618 368702 314854
rect 368786 314618 369022 314854
rect 368466 296938 368702 297174
rect 368786 296938 369022 297174
rect 368466 296618 368702 296854
rect 368786 296618 369022 296854
rect 368466 278938 368702 279174
rect 368786 278938 369022 279174
rect 368466 278618 368702 278854
rect 368786 278618 369022 278854
rect 368466 260938 368702 261174
rect 368786 260938 369022 261174
rect 368466 260618 368702 260854
rect 368786 260618 369022 260854
rect 368466 242938 368702 243174
rect 368786 242938 369022 243174
rect 368466 242618 368702 242854
rect 368786 242618 369022 242854
rect 368466 224938 368702 225174
rect 368786 224938 369022 225174
rect 368466 224618 368702 224854
rect 368786 224618 369022 224854
rect 368466 206938 368702 207174
rect 368786 206938 369022 207174
rect 368466 206618 368702 206854
rect 368786 206618 369022 206854
rect 368466 188938 368702 189174
rect 368786 188938 369022 189174
rect 368466 188618 368702 188854
rect 368786 188618 369022 188854
rect 368466 170938 368702 171174
rect 368786 170938 369022 171174
rect 368466 170618 368702 170854
rect 368786 170618 369022 170854
rect 368466 152938 368702 153174
rect 368786 152938 369022 153174
rect 368466 152618 368702 152854
rect 368786 152618 369022 152854
rect 368466 134938 368702 135174
rect 368786 134938 369022 135174
rect 368466 134618 368702 134854
rect 368786 134618 369022 134854
rect 368466 116938 368702 117174
rect 368786 116938 369022 117174
rect 368466 116618 368702 116854
rect 368786 116618 369022 116854
rect 368466 98938 368702 99174
rect 368786 98938 369022 99174
rect 368466 98618 368702 98854
rect 368786 98618 369022 98854
rect 368466 80938 368702 81174
rect 368786 80938 369022 81174
rect 368466 80618 368702 80854
rect 368786 80618 369022 80854
rect 368466 62938 368702 63174
rect 368786 62938 369022 63174
rect 368466 62618 368702 62854
rect 368786 62618 369022 62854
rect 368466 44938 368702 45174
rect 368786 44938 369022 45174
rect 368466 44618 368702 44854
rect 368786 44618 369022 44854
rect 368466 26938 368702 27174
rect 368786 26938 369022 27174
rect 368466 26618 368702 26854
rect 368786 26618 369022 26854
rect 368466 8938 368702 9174
rect 368786 8938 369022 9174
rect 368466 8618 368702 8854
rect 368786 8618 369022 8854
rect 368466 -2052 368702 -1816
rect 368786 -2052 369022 -1816
rect 368466 -2372 368702 -2136
rect 368786 -2372 369022 -2136
rect 372186 462776 372422 463012
rect 372506 462776 372742 463012
rect 372186 462456 372422 462692
rect 372506 462456 372742 462692
rect 372186 444658 372422 444894
rect 372506 444658 372742 444894
rect 372186 444338 372422 444574
rect 372506 444338 372742 444574
rect 372186 426658 372422 426894
rect 372506 426658 372742 426894
rect 372186 426338 372422 426574
rect 372506 426338 372742 426574
rect 372186 408658 372422 408894
rect 372506 408658 372742 408894
rect 372186 408338 372422 408574
rect 372506 408338 372742 408574
rect 372186 390658 372422 390894
rect 372506 390658 372742 390894
rect 372186 390338 372422 390574
rect 372506 390338 372742 390574
rect 372186 372658 372422 372894
rect 372506 372658 372742 372894
rect 372186 372338 372422 372574
rect 372506 372338 372742 372574
rect 372186 354658 372422 354894
rect 372506 354658 372742 354894
rect 372186 354338 372422 354574
rect 372506 354338 372742 354574
rect 372186 336658 372422 336894
rect 372506 336658 372742 336894
rect 372186 336338 372422 336574
rect 372506 336338 372742 336574
rect 372186 318658 372422 318894
rect 372506 318658 372742 318894
rect 372186 318338 372422 318574
rect 372506 318338 372742 318574
rect 372186 300658 372422 300894
rect 372506 300658 372742 300894
rect 372186 300338 372422 300574
rect 372506 300338 372742 300574
rect 372186 282658 372422 282894
rect 372506 282658 372742 282894
rect 372186 282338 372422 282574
rect 372506 282338 372742 282574
rect 372186 264658 372422 264894
rect 372506 264658 372742 264894
rect 372186 264338 372422 264574
rect 372506 264338 372742 264574
rect 372186 246658 372422 246894
rect 372506 246658 372742 246894
rect 372186 246338 372422 246574
rect 372506 246338 372742 246574
rect 372186 228658 372422 228894
rect 372506 228658 372742 228894
rect 372186 228338 372422 228574
rect 372506 228338 372742 228574
rect 372186 210658 372422 210894
rect 372506 210658 372742 210894
rect 372186 210338 372422 210574
rect 372506 210338 372742 210574
rect 372186 192658 372422 192894
rect 372506 192658 372742 192894
rect 372186 192338 372422 192574
rect 372506 192338 372742 192574
rect 372186 174658 372422 174894
rect 372506 174658 372742 174894
rect 372186 174338 372422 174574
rect 372506 174338 372742 174574
rect 372186 156658 372422 156894
rect 372506 156658 372742 156894
rect 372186 156338 372422 156574
rect 372506 156338 372742 156574
rect 372186 138658 372422 138894
rect 372506 138658 372742 138894
rect 372186 138338 372422 138574
rect 372506 138338 372742 138574
rect 372186 120658 372422 120894
rect 372506 120658 372742 120894
rect 372186 120338 372422 120574
rect 372506 120338 372742 120574
rect 372186 102658 372422 102894
rect 372506 102658 372742 102894
rect 372186 102338 372422 102574
rect 372506 102338 372742 102574
rect 372186 84658 372422 84894
rect 372506 84658 372742 84894
rect 372186 84338 372422 84574
rect 372506 84338 372742 84574
rect 372186 66658 372422 66894
rect 372506 66658 372742 66894
rect 372186 66338 372422 66574
rect 372506 66338 372742 66574
rect 372186 48658 372422 48894
rect 372506 48658 372742 48894
rect 372186 48338 372422 48574
rect 372506 48338 372742 48574
rect 372186 30658 372422 30894
rect 372506 30658 372742 30894
rect 372186 30338 372422 30574
rect 372506 30338 372742 30574
rect 372186 12658 372422 12894
rect 372506 12658 372742 12894
rect 372186 12338 372422 12574
rect 372506 12338 372742 12574
rect 372186 -3012 372422 -2776
rect 372506 -3012 372742 -2776
rect 372186 -3332 372422 -3096
rect 372506 -3332 372742 -3096
rect 375906 463736 376142 463972
rect 376226 463736 376462 463972
rect 375906 463416 376142 463652
rect 376226 463416 376462 463652
rect 375906 448378 376142 448614
rect 376226 448378 376462 448614
rect 375906 448058 376142 448294
rect 376226 448058 376462 448294
rect 375906 430378 376142 430614
rect 376226 430378 376462 430614
rect 375906 430058 376142 430294
rect 376226 430058 376462 430294
rect 375906 412378 376142 412614
rect 376226 412378 376462 412614
rect 375906 412058 376142 412294
rect 376226 412058 376462 412294
rect 375906 394378 376142 394614
rect 376226 394378 376462 394614
rect 375906 394058 376142 394294
rect 376226 394058 376462 394294
rect 375906 376378 376142 376614
rect 376226 376378 376462 376614
rect 375906 376058 376142 376294
rect 376226 376058 376462 376294
rect 375906 358378 376142 358614
rect 376226 358378 376462 358614
rect 375906 358058 376142 358294
rect 376226 358058 376462 358294
rect 375906 340378 376142 340614
rect 376226 340378 376462 340614
rect 375906 340058 376142 340294
rect 376226 340058 376462 340294
rect 375906 322378 376142 322614
rect 376226 322378 376462 322614
rect 375906 322058 376142 322294
rect 376226 322058 376462 322294
rect 375906 304378 376142 304614
rect 376226 304378 376462 304614
rect 375906 304058 376142 304294
rect 376226 304058 376462 304294
rect 375906 286378 376142 286614
rect 376226 286378 376462 286614
rect 375906 286058 376142 286294
rect 376226 286058 376462 286294
rect 375906 268378 376142 268614
rect 376226 268378 376462 268614
rect 375906 268058 376142 268294
rect 376226 268058 376462 268294
rect 375906 250378 376142 250614
rect 376226 250378 376462 250614
rect 375906 250058 376142 250294
rect 376226 250058 376462 250294
rect 375906 232378 376142 232614
rect 376226 232378 376462 232614
rect 375906 232058 376142 232294
rect 376226 232058 376462 232294
rect 375906 214378 376142 214614
rect 376226 214378 376462 214614
rect 375906 214058 376142 214294
rect 376226 214058 376462 214294
rect 375906 196378 376142 196614
rect 376226 196378 376462 196614
rect 375906 196058 376142 196294
rect 376226 196058 376462 196294
rect 375906 178378 376142 178614
rect 376226 178378 376462 178614
rect 375906 178058 376142 178294
rect 376226 178058 376462 178294
rect 375906 160378 376142 160614
rect 376226 160378 376462 160614
rect 375906 160058 376142 160294
rect 376226 160058 376462 160294
rect 375906 142378 376142 142614
rect 376226 142378 376462 142614
rect 375906 142058 376142 142294
rect 376226 142058 376462 142294
rect 375906 124378 376142 124614
rect 376226 124378 376462 124614
rect 375906 124058 376142 124294
rect 376226 124058 376462 124294
rect 375906 106378 376142 106614
rect 376226 106378 376462 106614
rect 375906 106058 376142 106294
rect 376226 106058 376462 106294
rect 375906 88378 376142 88614
rect 376226 88378 376462 88614
rect 375906 88058 376142 88294
rect 376226 88058 376462 88294
rect 375906 70378 376142 70614
rect 376226 70378 376462 70614
rect 375906 70058 376142 70294
rect 376226 70058 376462 70294
rect 375906 52378 376142 52614
rect 376226 52378 376462 52614
rect 375906 52058 376142 52294
rect 376226 52058 376462 52294
rect 375906 34378 376142 34614
rect 376226 34378 376462 34614
rect 375906 34058 376142 34294
rect 376226 34058 376462 34294
rect 375906 16378 376142 16614
rect 376226 16378 376462 16614
rect 375906 16058 376142 16294
rect 376226 16058 376462 16294
rect 375906 -3972 376142 -3736
rect 376226 -3972 376462 -3736
rect 375906 -4292 376142 -4056
rect 376226 -4292 376462 -4056
rect 382746 460856 382982 461092
rect 383066 460856 383302 461092
rect 382746 460536 382982 460772
rect 383066 460536 383302 460772
rect 382746 455218 382982 455454
rect 383066 455218 383302 455454
rect 382746 454898 382982 455134
rect 383066 454898 383302 455134
rect 382746 437218 382982 437454
rect 383066 437218 383302 437454
rect 382746 436898 382982 437134
rect 383066 436898 383302 437134
rect 382746 419218 382982 419454
rect 383066 419218 383302 419454
rect 382746 418898 382982 419134
rect 383066 418898 383302 419134
rect 382746 401218 382982 401454
rect 383066 401218 383302 401454
rect 382746 400898 382982 401134
rect 383066 400898 383302 401134
rect 382746 383218 382982 383454
rect 383066 383218 383302 383454
rect 382746 382898 382982 383134
rect 383066 382898 383302 383134
rect 382746 365218 382982 365454
rect 383066 365218 383302 365454
rect 382746 364898 382982 365134
rect 383066 364898 383302 365134
rect 382746 347218 382982 347454
rect 383066 347218 383302 347454
rect 382746 346898 382982 347134
rect 383066 346898 383302 347134
rect 382746 329218 382982 329454
rect 383066 329218 383302 329454
rect 382746 328898 382982 329134
rect 383066 328898 383302 329134
rect 382746 311218 382982 311454
rect 383066 311218 383302 311454
rect 382746 310898 382982 311134
rect 383066 310898 383302 311134
rect 382746 293218 382982 293454
rect 383066 293218 383302 293454
rect 382746 292898 382982 293134
rect 383066 292898 383302 293134
rect 382746 275218 382982 275454
rect 383066 275218 383302 275454
rect 382746 274898 382982 275134
rect 383066 274898 383302 275134
rect 382746 257218 382982 257454
rect 383066 257218 383302 257454
rect 382746 256898 382982 257134
rect 383066 256898 383302 257134
rect 382746 239218 382982 239454
rect 383066 239218 383302 239454
rect 382746 238898 382982 239134
rect 383066 238898 383302 239134
rect 382746 221218 382982 221454
rect 383066 221218 383302 221454
rect 382746 220898 382982 221134
rect 383066 220898 383302 221134
rect 382746 203218 382982 203454
rect 383066 203218 383302 203454
rect 382746 202898 382982 203134
rect 383066 202898 383302 203134
rect 382746 185218 382982 185454
rect 383066 185218 383302 185454
rect 382746 184898 382982 185134
rect 383066 184898 383302 185134
rect 382746 167218 382982 167454
rect 383066 167218 383302 167454
rect 382746 166898 382982 167134
rect 383066 166898 383302 167134
rect 382746 149218 382982 149454
rect 383066 149218 383302 149454
rect 382746 148898 382982 149134
rect 383066 148898 383302 149134
rect 382746 131218 382982 131454
rect 383066 131218 383302 131454
rect 382746 130898 382982 131134
rect 383066 130898 383302 131134
rect 382746 113218 382982 113454
rect 383066 113218 383302 113454
rect 382746 112898 382982 113134
rect 383066 112898 383302 113134
rect 382746 95218 382982 95454
rect 383066 95218 383302 95454
rect 382746 94898 382982 95134
rect 383066 94898 383302 95134
rect 382746 77218 382982 77454
rect 383066 77218 383302 77454
rect 382746 76898 382982 77134
rect 383066 76898 383302 77134
rect 382746 59218 382982 59454
rect 383066 59218 383302 59454
rect 382746 58898 382982 59134
rect 383066 58898 383302 59134
rect 382746 41218 382982 41454
rect 383066 41218 383302 41454
rect 382746 40898 382982 41134
rect 383066 40898 383302 41134
rect 382746 23218 382982 23454
rect 383066 23218 383302 23454
rect 382746 22898 382982 23134
rect 383066 22898 383302 23134
rect 382746 5218 382982 5454
rect 383066 5218 383302 5454
rect 382746 4898 382982 5134
rect 383066 4898 383302 5134
rect 382746 -1092 382982 -856
rect 383066 -1092 383302 -856
rect 382746 -1412 382982 -1176
rect 383066 -1412 383302 -1176
rect 386466 461816 386702 462052
rect 386786 461816 387022 462052
rect 386466 461496 386702 461732
rect 386786 461496 387022 461732
rect 386466 440938 386702 441174
rect 386786 440938 387022 441174
rect 386466 440618 386702 440854
rect 386786 440618 387022 440854
rect 386466 422938 386702 423174
rect 386786 422938 387022 423174
rect 386466 422618 386702 422854
rect 386786 422618 387022 422854
rect 386466 404938 386702 405174
rect 386786 404938 387022 405174
rect 386466 404618 386702 404854
rect 386786 404618 387022 404854
rect 386466 386938 386702 387174
rect 386786 386938 387022 387174
rect 386466 386618 386702 386854
rect 386786 386618 387022 386854
rect 386466 368938 386702 369174
rect 386786 368938 387022 369174
rect 386466 368618 386702 368854
rect 386786 368618 387022 368854
rect 386466 350938 386702 351174
rect 386786 350938 387022 351174
rect 386466 350618 386702 350854
rect 386786 350618 387022 350854
rect 386466 332938 386702 333174
rect 386786 332938 387022 333174
rect 386466 332618 386702 332854
rect 386786 332618 387022 332854
rect 386466 314938 386702 315174
rect 386786 314938 387022 315174
rect 386466 314618 386702 314854
rect 386786 314618 387022 314854
rect 386466 296938 386702 297174
rect 386786 296938 387022 297174
rect 386466 296618 386702 296854
rect 386786 296618 387022 296854
rect 386466 278938 386702 279174
rect 386786 278938 387022 279174
rect 386466 278618 386702 278854
rect 386786 278618 387022 278854
rect 386466 260938 386702 261174
rect 386786 260938 387022 261174
rect 386466 260618 386702 260854
rect 386786 260618 387022 260854
rect 386466 242938 386702 243174
rect 386786 242938 387022 243174
rect 386466 242618 386702 242854
rect 386786 242618 387022 242854
rect 386466 224938 386702 225174
rect 386786 224938 387022 225174
rect 386466 224618 386702 224854
rect 386786 224618 387022 224854
rect 386466 206938 386702 207174
rect 386786 206938 387022 207174
rect 386466 206618 386702 206854
rect 386786 206618 387022 206854
rect 386466 188938 386702 189174
rect 386786 188938 387022 189174
rect 386466 188618 386702 188854
rect 386786 188618 387022 188854
rect 386466 170938 386702 171174
rect 386786 170938 387022 171174
rect 386466 170618 386702 170854
rect 386786 170618 387022 170854
rect 386466 152938 386702 153174
rect 386786 152938 387022 153174
rect 386466 152618 386702 152854
rect 386786 152618 387022 152854
rect 386466 134938 386702 135174
rect 386786 134938 387022 135174
rect 386466 134618 386702 134854
rect 386786 134618 387022 134854
rect 386466 116938 386702 117174
rect 386786 116938 387022 117174
rect 386466 116618 386702 116854
rect 386786 116618 387022 116854
rect 386466 98938 386702 99174
rect 386786 98938 387022 99174
rect 386466 98618 386702 98854
rect 386786 98618 387022 98854
rect 386466 80938 386702 81174
rect 386786 80938 387022 81174
rect 386466 80618 386702 80854
rect 386786 80618 387022 80854
rect 386466 62938 386702 63174
rect 386786 62938 387022 63174
rect 386466 62618 386702 62854
rect 386786 62618 387022 62854
rect 386466 44938 386702 45174
rect 386786 44938 387022 45174
rect 386466 44618 386702 44854
rect 386786 44618 387022 44854
rect 386466 26938 386702 27174
rect 386786 26938 387022 27174
rect 386466 26618 386702 26854
rect 386786 26618 387022 26854
rect 386466 8938 386702 9174
rect 386786 8938 387022 9174
rect 386466 8618 386702 8854
rect 386786 8618 387022 8854
rect 386466 -2052 386702 -1816
rect 386786 -2052 387022 -1816
rect 386466 -2372 386702 -2136
rect 386786 -2372 387022 -2136
rect 390186 462776 390422 463012
rect 390506 462776 390742 463012
rect 390186 462456 390422 462692
rect 390506 462456 390742 462692
rect 390186 444658 390422 444894
rect 390506 444658 390742 444894
rect 390186 444338 390422 444574
rect 390506 444338 390742 444574
rect 390186 426658 390422 426894
rect 390506 426658 390742 426894
rect 390186 426338 390422 426574
rect 390506 426338 390742 426574
rect 390186 408658 390422 408894
rect 390506 408658 390742 408894
rect 390186 408338 390422 408574
rect 390506 408338 390742 408574
rect 390186 390658 390422 390894
rect 390506 390658 390742 390894
rect 390186 390338 390422 390574
rect 390506 390338 390742 390574
rect 390186 372658 390422 372894
rect 390506 372658 390742 372894
rect 390186 372338 390422 372574
rect 390506 372338 390742 372574
rect 390186 354658 390422 354894
rect 390506 354658 390742 354894
rect 390186 354338 390422 354574
rect 390506 354338 390742 354574
rect 390186 336658 390422 336894
rect 390506 336658 390742 336894
rect 390186 336338 390422 336574
rect 390506 336338 390742 336574
rect 390186 318658 390422 318894
rect 390506 318658 390742 318894
rect 390186 318338 390422 318574
rect 390506 318338 390742 318574
rect 390186 300658 390422 300894
rect 390506 300658 390742 300894
rect 390186 300338 390422 300574
rect 390506 300338 390742 300574
rect 390186 282658 390422 282894
rect 390506 282658 390742 282894
rect 390186 282338 390422 282574
rect 390506 282338 390742 282574
rect 390186 264658 390422 264894
rect 390506 264658 390742 264894
rect 390186 264338 390422 264574
rect 390506 264338 390742 264574
rect 390186 246658 390422 246894
rect 390506 246658 390742 246894
rect 390186 246338 390422 246574
rect 390506 246338 390742 246574
rect 390186 228658 390422 228894
rect 390506 228658 390742 228894
rect 390186 228338 390422 228574
rect 390506 228338 390742 228574
rect 390186 210658 390422 210894
rect 390506 210658 390742 210894
rect 390186 210338 390422 210574
rect 390506 210338 390742 210574
rect 390186 192658 390422 192894
rect 390506 192658 390742 192894
rect 390186 192338 390422 192574
rect 390506 192338 390742 192574
rect 390186 174658 390422 174894
rect 390506 174658 390742 174894
rect 390186 174338 390422 174574
rect 390506 174338 390742 174574
rect 390186 156658 390422 156894
rect 390506 156658 390742 156894
rect 390186 156338 390422 156574
rect 390506 156338 390742 156574
rect 390186 138658 390422 138894
rect 390506 138658 390742 138894
rect 390186 138338 390422 138574
rect 390506 138338 390742 138574
rect 390186 120658 390422 120894
rect 390506 120658 390742 120894
rect 390186 120338 390422 120574
rect 390506 120338 390742 120574
rect 390186 102658 390422 102894
rect 390506 102658 390742 102894
rect 390186 102338 390422 102574
rect 390506 102338 390742 102574
rect 390186 84658 390422 84894
rect 390506 84658 390742 84894
rect 390186 84338 390422 84574
rect 390506 84338 390742 84574
rect 390186 66658 390422 66894
rect 390506 66658 390742 66894
rect 390186 66338 390422 66574
rect 390506 66338 390742 66574
rect 390186 48658 390422 48894
rect 390506 48658 390742 48894
rect 390186 48338 390422 48574
rect 390506 48338 390742 48574
rect 390186 30658 390422 30894
rect 390506 30658 390742 30894
rect 390186 30338 390422 30574
rect 390506 30338 390742 30574
rect 390186 12658 390422 12894
rect 390506 12658 390742 12894
rect 390186 12338 390422 12574
rect 390506 12338 390742 12574
rect 390186 -3012 390422 -2776
rect 390506 -3012 390742 -2776
rect 390186 -3332 390422 -3096
rect 390506 -3332 390742 -3096
rect 393906 463736 394142 463972
rect 394226 463736 394462 463972
rect 393906 463416 394142 463652
rect 394226 463416 394462 463652
rect 393906 448378 394142 448614
rect 394226 448378 394462 448614
rect 393906 448058 394142 448294
rect 394226 448058 394462 448294
rect 393906 430378 394142 430614
rect 394226 430378 394462 430614
rect 393906 430058 394142 430294
rect 394226 430058 394462 430294
rect 393906 412378 394142 412614
rect 394226 412378 394462 412614
rect 393906 412058 394142 412294
rect 394226 412058 394462 412294
rect 393906 394378 394142 394614
rect 394226 394378 394462 394614
rect 393906 394058 394142 394294
rect 394226 394058 394462 394294
rect 393906 376378 394142 376614
rect 394226 376378 394462 376614
rect 393906 376058 394142 376294
rect 394226 376058 394462 376294
rect 393906 358378 394142 358614
rect 394226 358378 394462 358614
rect 393906 358058 394142 358294
rect 394226 358058 394462 358294
rect 393906 340378 394142 340614
rect 394226 340378 394462 340614
rect 393906 340058 394142 340294
rect 394226 340058 394462 340294
rect 393906 322378 394142 322614
rect 394226 322378 394462 322614
rect 393906 322058 394142 322294
rect 394226 322058 394462 322294
rect 393906 304378 394142 304614
rect 394226 304378 394462 304614
rect 393906 304058 394142 304294
rect 394226 304058 394462 304294
rect 393906 286378 394142 286614
rect 394226 286378 394462 286614
rect 393906 286058 394142 286294
rect 394226 286058 394462 286294
rect 393906 268378 394142 268614
rect 394226 268378 394462 268614
rect 393906 268058 394142 268294
rect 394226 268058 394462 268294
rect 393906 250378 394142 250614
rect 394226 250378 394462 250614
rect 393906 250058 394142 250294
rect 394226 250058 394462 250294
rect 393906 232378 394142 232614
rect 394226 232378 394462 232614
rect 393906 232058 394142 232294
rect 394226 232058 394462 232294
rect 393906 214378 394142 214614
rect 394226 214378 394462 214614
rect 393906 214058 394142 214294
rect 394226 214058 394462 214294
rect 393906 196378 394142 196614
rect 394226 196378 394462 196614
rect 393906 196058 394142 196294
rect 394226 196058 394462 196294
rect 393906 178378 394142 178614
rect 394226 178378 394462 178614
rect 393906 178058 394142 178294
rect 394226 178058 394462 178294
rect 393906 160378 394142 160614
rect 394226 160378 394462 160614
rect 393906 160058 394142 160294
rect 394226 160058 394462 160294
rect 393906 142378 394142 142614
rect 394226 142378 394462 142614
rect 393906 142058 394142 142294
rect 394226 142058 394462 142294
rect 393906 124378 394142 124614
rect 394226 124378 394462 124614
rect 393906 124058 394142 124294
rect 394226 124058 394462 124294
rect 393906 106378 394142 106614
rect 394226 106378 394462 106614
rect 393906 106058 394142 106294
rect 394226 106058 394462 106294
rect 393906 88378 394142 88614
rect 394226 88378 394462 88614
rect 393906 88058 394142 88294
rect 394226 88058 394462 88294
rect 393906 70378 394142 70614
rect 394226 70378 394462 70614
rect 393906 70058 394142 70294
rect 394226 70058 394462 70294
rect 393906 52378 394142 52614
rect 394226 52378 394462 52614
rect 393906 52058 394142 52294
rect 394226 52058 394462 52294
rect 393906 34378 394142 34614
rect 394226 34378 394462 34614
rect 393906 34058 394142 34294
rect 394226 34058 394462 34294
rect 393906 16378 394142 16614
rect 394226 16378 394462 16614
rect 393906 16058 394142 16294
rect 394226 16058 394462 16294
rect 393906 -3972 394142 -3736
rect 394226 -3972 394462 -3736
rect 393906 -4292 394142 -4056
rect 394226 -4292 394462 -4056
rect 400746 460856 400982 461092
rect 401066 460856 401302 461092
rect 400746 460536 400982 460772
rect 401066 460536 401302 460772
rect 400746 455218 400982 455454
rect 401066 455218 401302 455454
rect 400746 454898 400982 455134
rect 401066 454898 401302 455134
rect 400746 437218 400982 437454
rect 401066 437218 401302 437454
rect 400746 436898 400982 437134
rect 401066 436898 401302 437134
rect 400746 419218 400982 419454
rect 401066 419218 401302 419454
rect 400746 418898 400982 419134
rect 401066 418898 401302 419134
rect 400746 401218 400982 401454
rect 401066 401218 401302 401454
rect 400746 400898 400982 401134
rect 401066 400898 401302 401134
rect 400746 383218 400982 383454
rect 401066 383218 401302 383454
rect 400746 382898 400982 383134
rect 401066 382898 401302 383134
rect 400746 365218 400982 365454
rect 401066 365218 401302 365454
rect 400746 364898 400982 365134
rect 401066 364898 401302 365134
rect 400746 347218 400982 347454
rect 401066 347218 401302 347454
rect 400746 346898 400982 347134
rect 401066 346898 401302 347134
rect 400746 329218 400982 329454
rect 401066 329218 401302 329454
rect 400746 328898 400982 329134
rect 401066 328898 401302 329134
rect 400746 311218 400982 311454
rect 401066 311218 401302 311454
rect 400746 310898 400982 311134
rect 401066 310898 401302 311134
rect 400746 293218 400982 293454
rect 401066 293218 401302 293454
rect 400746 292898 400982 293134
rect 401066 292898 401302 293134
rect 400746 275218 400982 275454
rect 401066 275218 401302 275454
rect 400746 274898 400982 275134
rect 401066 274898 401302 275134
rect 400746 257218 400982 257454
rect 401066 257218 401302 257454
rect 400746 256898 400982 257134
rect 401066 256898 401302 257134
rect 400746 239218 400982 239454
rect 401066 239218 401302 239454
rect 400746 238898 400982 239134
rect 401066 238898 401302 239134
rect 400746 221218 400982 221454
rect 401066 221218 401302 221454
rect 400746 220898 400982 221134
rect 401066 220898 401302 221134
rect 400746 203218 400982 203454
rect 401066 203218 401302 203454
rect 400746 202898 400982 203134
rect 401066 202898 401302 203134
rect 400746 185218 400982 185454
rect 401066 185218 401302 185454
rect 400746 184898 400982 185134
rect 401066 184898 401302 185134
rect 400746 167218 400982 167454
rect 401066 167218 401302 167454
rect 400746 166898 400982 167134
rect 401066 166898 401302 167134
rect 400746 149218 400982 149454
rect 401066 149218 401302 149454
rect 400746 148898 400982 149134
rect 401066 148898 401302 149134
rect 400746 131218 400982 131454
rect 401066 131218 401302 131454
rect 400746 130898 400982 131134
rect 401066 130898 401302 131134
rect 400746 113218 400982 113454
rect 401066 113218 401302 113454
rect 400746 112898 400982 113134
rect 401066 112898 401302 113134
rect 400746 95218 400982 95454
rect 401066 95218 401302 95454
rect 400746 94898 400982 95134
rect 401066 94898 401302 95134
rect 400746 77218 400982 77454
rect 401066 77218 401302 77454
rect 400746 76898 400982 77134
rect 401066 76898 401302 77134
rect 400746 59218 400982 59454
rect 401066 59218 401302 59454
rect 400746 58898 400982 59134
rect 401066 58898 401302 59134
rect 400746 41218 400982 41454
rect 401066 41218 401302 41454
rect 400746 40898 400982 41134
rect 401066 40898 401302 41134
rect 400746 23218 400982 23454
rect 401066 23218 401302 23454
rect 400746 22898 400982 23134
rect 401066 22898 401302 23134
rect 400746 5218 400982 5454
rect 401066 5218 401302 5454
rect 400746 4898 400982 5134
rect 401066 4898 401302 5134
rect 400746 -1092 400982 -856
rect 401066 -1092 401302 -856
rect 400746 -1412 400982 -1176
rect 401066 -1412 401302 -1176
rect 404466 461816 404702 462052
rect 404786 461816 405022 462052
rect 404466 461496 404702 461732
rect 404786 461496 405022 461732
rect 404466 440938 404702 441174
rect 404786 440938 405022 441174
rect 404466 440618 404702 440854
rect 404786 440618 405022 440854
rect 404466 422938 404702 423174
rect 404786 422938 405022 423174
rect 404466 422618 404702 422854
rect 404786 422618 405022 422854
rect 404466 404938 404702 405174
rect 404786 404938 405022 405174
rect 404466 404618 404702 404854
rect 404786 404618 405022 404854
rect 404466 386938 404702 387174
rect 404786 386938 405022 387174
rect 404466 386618 404702 386854
rect 404786 386618 405022 386854
rect 404466 368938 404702 369174
rect 404786 368938 405022 369174
rect 404466 368618 404702 368854
rect 404786 368618 405022 368854
rect 404466 350938 404702 351174
rect 404786 350938 405022 351174
rect 404466 350618 404702 350854
rect 404786 350618 405022 350854
rect 404466 332938 404702 333174
rect 404786 332938 405022 333174
rect 404466 332618 404702 332854
rect 404786 332618 405022 332854
rect 404466 314938 404702 315174
rect 404786 314938 405022 315174
rect 404466 314618 404702 314854
rect 404786 314618 405022 314854
rect 404466 296938 404702 297174
rect 404786 296938 405022 297174
rect 404466 296618 404702 296854
rect 404786 296618 405022 296854
rect 404466 278938 404702 279174
rect 404786 278938 405022 279174
rect 404466 278618 404702 278854
rect 404786 278618 405022 278854
rect 404466 260938 404702 261174
rect 404786 260938 405022 261174
rect 404466 260618 404702 260854
rect 404786 260618 405022 260854
rect 404466 242938 404702 243174
rect 404786 242938 405022 243174
rect 404466 242618 404702 242854
rect 404786 242618 405022 242854
rect 404466 224938 404702 225174
rect 404786 224938 405022 225174
rect 404466 224618 404702 224854
rect 404786 224618 405022 224854
rect 404466 206938 404702 207174
rect 404786 206938 405022 207174
rect 404466 206618 404702 206854
rect 404786 206618 405022 206854
rect 404466 188938 404702 189174
rect 404786 188938 405022 189174
rect 404466 188618 404702 188854
rect 404786 188618 405022 188854
rect 404466 170938 404702 171174
rect 404786 170938 405022 171174
rect 404466 170618 404702 170854
rect 404786 170618 405022 170854
rect 404466 152938 404702 153174
rect 404786 152938 405022 153174
rect 404466 152618 404702 152854
rect 404786 152618 405022 152854
rect 404466 134938 404702 135174
rect 404786 134938 405022 135174
rect 404466 134618 404702 134854
rect 404786 134618 405022 134854
rect 404466 116938 404702 117174
rect 404786 116938 405022 117174
rect 404466 116618 404702 116854
rect 404786 116618 405022 116854
rect 404466 98938 404702 99174
rect 404786 98938 405022 99174
rect 404466 98618 404702 98854
rect 404786 98618 405022 98854
rect 404466 80938 404702 81174
rect 404786 80938 405022 81174
rect 404466 80618 404702 80854
rect 404786 80618 405022 80854
rect 404466 62938 404702 63174
rect 404786 62938 405022 63174
rect 404466 62618 404702 62854
rect 404786 62618 405022 62854
rect 404466 44938 404702 45174
rect 404786 44938 405022 45174
rect 404466 44618 404702 44854
rect 404786 44618 405022 44854
rect 404466 26938 404702 27174
rect 404786 26938 405022 27174
rect 404466 26618 404702 26854
rect 404786 26618 405022 26854
rect 404466 8938 404702 9174
rect 404786 8938 405022 9174
rect 404466 8618 404702 8854
rect 404786 8618 405022 8854
rect 404466 -2052 404702 -1816
rect 404786 -2052 405022 -1816
rect 404466 -2372 404702 -2136
rect 404786 -2372 405022 -2136
rect 408186 462776 408422 463012
rect 408506 462776 408742 463012
rect 408186 462456 408422 462692
rect 408506 462456 408742 462692
rect 408186 444658 408422 444894
rect 408506 444658 408742 444894
rect 408186 444338 408422 444574
rect 408506 444338 408742 444574
rect 408186 426658 408422 426894
rect 408506 426658 408742 426894
rect 408186 426338 408422 426574
rect 408506 426338 408742 426574
rect 408186 408658 408422 408894
rect 408506 408658 408742 408894
rect 408186 408338 408422 408574
rect 408506 408338 408742 408574
rect 408186 390658 408422 390894
rect 408506 390658 408742 390894
rect 408186 390338 408422 390574
rect 408506 390338 408742 390574
rect 408186 372658 408422 372894
rect 408506 372658 408742 372894
rect 408186 372338 408422 372574
rect 408506 372338 408742 372574
rect 408186 354658 408422 354894
rect 408506 354658 408742 354894
rect 408186 354338 408422 354574
rect 408506 354338 408742 354574
rect 408186 336658 408422 336894
rect 408506 336658 408742 336894
rect 408186 336338 408422 336574
rect 408506 336338 408742 336574
rect 408186 318658 408422 318894
rect 408506 318658 408742 318894
rect 408186 318338 408422 318574
rect 408506 318338 408742 318574
rect 408186 300658 408422 300894
rect 408506 300658 408742 300894
rect 408186 300338 408422 300574
rect 408506 300338 408742 300574
rect 408186 282658 408422 282894
rect 408506 282658 408742 282894
rect 408186 282338 408422 282574
rect 408506 282338 408742 282574
rect 408186 264658 408422 264894
rect 408506 264658 408742 264894
rect 408186 264338 408422 264574
rect 408506 264338 408742 264574
rect 408186 246658 408422 246894
rect 408506 246658 408742 246894
rect 408186 246338 408422 246574
rect 408506 246338 408742 246574
rect 408186 228658 408422 228894
rect 408506 228658 408742 228894
rect 408186 228338 408422 228574
rect 408506 228338 408742 228574
rect 408186 210658 408422 210894
rect 408506 210658 408742 210894
rect 408186 210338 408422 210574
rect 408506 210338 408742 210574
rect 408186 192658 408422 192894
rect 408506 192658 408742 192894
rect 408186 192338 408422 192574
rect 408506 192338 408742 192574
rect 408186 174658 408422 174894
rect 408506 174658 408742 174894
rect 408186 174338 408422 174574
rect 408506 174338 408742 174574
rect 408186 156658 408422 156894
rect 408506 156658 408742 156894
rect 408186 156338 408422 156574
rect 408506 156338 408742 156574
rect 408186 138658 408422 138894
rect 408506 138658 408742 138894
rect 408186 138338 408422 138574
rect 408506 138338 408742 138574
rect 408186 120658 408422 120894
rect 408506 120658 408742 120894
rect 408186 120338 408422 120574
rect 408506 120338 408742 120574
rect 408186 102658 408422 102894
rect 408506 102658 408742 102894
rect 408186 102338 408422 102574
rect 408506 102338 408742 102574
rect 408186 84658 408422 84894
rect 408506 84658 408742 84894
rect 408186 84338 408422 84574
rect 408506 84338 408742 84574
rect 408186 66658 408422 66894
rect 408506 66658 408742 66894
rect 408186 66338 408422 66574
rect 408506 66338 408742 66574
rect 408186 48658 408422 48894
rect 408506 48658 408742 48894
rect 408186 48338 408422 48574
rect 408506 48338 408742 48574
rect 408186 30658 408422 30894
rect 408506 30658 408742 30894
rect 408186 30338 408422 30574
rect 408506 30338 408742 30574
rect 408186 12658 408422 12894
rect 408506 12658 408742 12894
rect 408186 12338 408422 12574
rect 408506 12338 408742 12574
rect 408186 -3012 408422 -2776
rect 408506 -3012 408742 -2776
rect 408186 -3332 408422 -3096
rect 408506 -3332 408742 -3096
rect 411906 463736 412142 463972
rect 412226 463736 412462 463972
rect 411906 463416 412142 463652
rect 412226 463416 412462 463652
rect 411906 448378 412142 448614
rect 412226 448378 412462 448614
rect 411906 448058 412142 448294
rect 412226 448058 412462 448294
rect 411906 430378 412142 430614
rect 412226 430378 412462 430614
rect 411906 430058 412142 430294
rect 412226 430058 412462 430294
rect 411906 412378 412142 412614
rect 412226 412378 412462 412614
rect 411906 412058 412142 412294
rect 412226 412058 412462 412294
rect 411906 394378 412142 394614
rect 412226 394378 412462 394614
rect 411906 394058 412142 394294
rect 412226 394058 412462 394294
rect 411906 376378 412142 376614
rect 412226 376378 412462 376614
rect 411906 376058 412142 376294
rect 412226 376058 412462 376294
rect 411906 358378 412142 358614
rect 412226 358378 412462 358614
rect 411906 358058 412142 358294
rect 412226 358058 412462 358294
rect 411906 340378 412142 340614
rect 412226 340378 412462 340614
rect 411906 340058 412142 340294
rect 412226 340058 412462 340294
rect 411906 322378 412142 322614
rect 412226 322378 412462 322614
rect 411906 322058 412142 322294
rect 412226 322058 412462 322294
rect 411906 304378 412142 304614
rect 412226 304378 412462 304614
rect 411906 304058 412142 304294
rect 412226 304058 412462 304294
rect 411906 286378 412142 286614
rect 412226 286378 412462 286614
rect 411906 286058 412142 286294
rect 412226 286058 412462 286294
rect 411906 268378 412142 268614
rect 412226 268378 412462 268614
rect 411906 268058 412142 268294
rect 412226 268058 412462 268294
rect 411906 250378 412142 250614
rect 412226 250378 412462 250614
rect 411906 250058 412142 250294
rect 412226 250058 412462 250294
rect 411906 232378 412142 232614
rect 412226 232378 412462 232614
rect 411906 232058 412142 232294
rect 412226 232058 412462 232294
rect 411906 214378 412142 214614
rect 412226 214378 412462 214614
rect 411906 214058 412142 214294
rect 412226 214058 412462 214294
rect 411906 196378 412142 196614
rect 412226 196378 412462 196614
rect 411906 196058 412142 196294
rect 412226 196058 412462 196294
rect 411906 178378 412142 178614
rect 412226 178378 412462 178614
rect 411906 178058 412142 178294
rect 412226 178058 412462 178294
rect 411906 160378 412142 160614
rect 412226 160378 412462 160614
rect 411906 160058 412142 160294
rect 412226 160058 412462 160294
rect 411906 142378 412142 142614
rect 412226 142378 412462 142614
rect 411906 142058 412142 142294
rect 412226 142058 412462 142294
rect 411906 124378 412142 124614
rect 412226 124378 412462 124614
rect 411906 124058 412142 124294
rect 412226 124058 412462 124294
rect 411906 106378 412142 106614
rect 412226 106378 412462 106614
rect 411906 106058 412142 106294
rect 412226 106058 412462 106294
rect 411906 88378 412142 88614
rect 412226 88378 412462 88614
rect 411906 88058 412142 88294
rect 412226 88058 412462 88294
rect 411906 70378 412142 70614
rect 412226 70378 412462 70614
rect 411906 70058 412142 70294
rect 412226 70058 412462 70294
rect 411906 52378 412142 52614
rect 412226 52378 412462 52614
rect 411906 52058 412142 52294
rect 412226 52058 412462 52294
rect 411906 34378 412142 34614
rect 412226 34378 412462 34614
rect 411906 34058 412142 34294
rect 412226 34058 412462 34294
rect 411906 16378 412142 16614
rect 412226 16378 412462 16614
rect 411906 16058 412142 16294
rect 412226 16058 412462 16294
rect 411906 -3972 412142 -3736
rect 412226 -3972 412462 -3736
rect 411906 -4292 412142 -4056
rect 412226 -4292 412462 -4056
rect 418746 460856 418982 461092
rect 419066 460856 419302 461092
rect 418746 460536 418982 460772
rect 419066 460536 419302 460772
rect 418746 455218 418982 455454
rect 419066 455218 419302 455454
rect 418746 454898 418982 455134
rect 419066 454898 419302 455134
rect 418746 437218 418982 437454
rect 419066 437218 419302 437454
rect 418746 436898 418982 437134
rect 419066 436898 419302 437134
rect 418746 419218 418982 419454
rect 419066 419218 419302 419454
rect 418746 418898 418982 419134
rect 419066 418898 419302 419134
rect 418746 401218 418982 401454
rect 419066 401218 419302 401454
rect 418746 400898 418982 401134
rect 419066 400898 419302 401134
rect 418746 383218 418982 383454
rect 419066 383218 419302 383454
rect 418746 382898 418982 383134
rect 419066 382898 419302 383134
rect 418746 365218 418982 365454
rect 419066 365218 419302 365454
rect 418746 364898 418982 365134
rect 419066 364898 419302 365134
rect 418746 347218 418982 347454
rect 419066 347218 419302 347454
rect 418746 346898 418982 347134
rect 419066 346898 419302 347134
rect 418746 329218 418982 329454
rect 419066 329218 419302 329454
rect 418746 328898 418982 329134
rect 419066 328898 419302 329134
rect 418746 311218 418982 311454
rect 419066 311218 419302 311454
rect 418746 310898 418982 311134
rect 419066 310898 419302 311134
rect 418746 293218 418982 293454
rect 419066 293218 419302 293454
rect 418746 292898 418982 293134
rect 419066 292898 419302 293134
rect 418746 275218 418982 275454
rect 419066 275218 419302 275454
rect 418746 274898 418982 275134
rect 419066 274898 419302 275134
rect 418746 257218 418982 257454
rect 419066 257218 419302 257454
rect 418746 256898 418982 257134
rect 419066 256898 419302 257134
rect 418746 239218 418982 239454
rect 419066 239218 419302 239454
rect 418746 238898 418982 239134
rect 419066 238898 419302 239134
rect 418746 221218 418982 221454
rect 419066 221218 419302 221454
rect 418746 220898 418982 221134
rect 419066 220898 419302 221134
rect 418746 203218 418982 203454
rect 419066 203218 419302 203454
rect 418746 202898 418982 203134
rect 419066 202898 419302 203134
rect 418746 185218 418982 185454
rect 419066 185218 419302 185454
rect 418746 184898 418982 185134
rect 419066 184898 419302 185134
rect 418746 167218 418982 167454
rect 419066 167218 419302 167454
rect 418746 166898 418982 167134
rect 419066 166898 419302 167134
rect 418746 149218 418982 149454
rect 419066 149218 419302 149454
rect 418746 148898 418982 149134
rect 419066 148898 419302 149134
rect 418746 131218 418982 131454
rect 419066 131218 419302 131454
rect 418746 130898 418982 131134
rect 419066 130898 419302 131134
rect 418746 113218 418982 113454
rect 419066 113218 419302 113454
rect 418746 112898 418982 113134
rect 419066 112898 419302 113134
rect 418746 95218 418982 95454
rect 419066 95218 419302 95454
rect 418746 94898 418982 95134
rect 419066 94898 419302 95134
rect 418746 77218 418982 77454
rect 419066 77218 419302 77454
rect 418746 76898 418982 77134
rect 419066 76898 419302 77134
rect 418746 59218 418982 59454
rect 419066 59218 419302 59454
rect 418746 58898 418982 59134
rect 419066 58898 419302 59134
rect 418746 41218 418982 41454
rect 419066 41218 419302 41454
rect 418746 40898 418982 41134
rect 419066 40898 419302 41134
rect 418746 23218 418982 23454
rect 419066 23218 419302 23454
rect 418746 22898 418982 23134
rect 419066 22898 419302 23134
rect 418746 5218 418982 5454
rect 419066 5218 419302 5454
rect 418746 4898 418982 5134
rect 419066 4898 419302 5134
rect 418746 -1092 418982 -856
rect 419066 -1092 419302 -856
rect 418746 -1412 418982 -1176
rect 419066 -1412 419302 -1176
rect 422466 461816 422702 462052
rect 422786 461816 423022 462052
rect 422466 461496 422702 461732
rect 422786 461496 423022 461732
rect 422466 440938 422702 441174
rect 422786 440938 423022 441174
rect 422466 440618 422702 440854
rect 422786 440618 423022 440854
rect 422466 422938 422702 423174
rect 422786 422938 423022 423174
rect 422466 422618 422702 422854
rect 422786 422618 423022 422854
rect 422466 404938 422702 405174
rect 422786 404938 423022 405174
rect 422466 404618 422702 404854
rect 422786 404618 423022 404854
rect 422466 386938 422702 387174
rect 422786 386938 423022 387174
rect 422466 386618 422702 386854
rect 422786 386618 423022 386854
rect 422466 368938 422702 369174
rect 422786 368938 423022 369174
rect 422466 368618 422702 368854
rect 422786 368618 423022 368854
rect 422466 350938 422702 351174
rect 422786 350938 423022 351174
rect 422466 350618 422702 350854
rect 422786 350618 423022 350854
rect 422466 332938 422702 333174
rect 422786 332938 423022 333174
rect 422466 332618 422702 332854
rect 422786 332618 423022 332854
rect 422466 314938 422702 315174
rect 422786 314938 423022 315174
rect 422466 314618 422702 314854
rect 422786 314618 423022 314854
rect 422466 296938 422702 297174
rect 422786 296938 423022 297174
rect 422466 296618 422702 296854
rect 422786 296618 423022 296854
rect 422466 278938 422702 279174
rect 422786 278938 423022 279174
rect 422466 278618 422702 278854
rect 422786 278618 423022 278854
rect 422466 260938 422702 261174
rect 422786 260938 423022 261174
rect 422466 260618 422702 260854
rect 422786 260618 423022 260854
rect 422466 242938 422702 243174
rect 422786 242938 423022 243174
rect 422466 242618 422702 242854
rect 422786 242618 423022 242854
rect 422466 224938 422702 225174
rect 422786 224938 423022 225174
rect 422466 224618 422702 224854
rect 422786 224618 423022 224854
rect 422466 206938 422702 207174
rect 422786 206938 423022 207174
rect 422466 206618 422702 206854
rect 422786 206618 423022 206854
rect 422466 188938 422702 189174
rect 422786 188938 423022 189174
rect 422466 188618 422702 188854
rect 422786 188618 423022 188854
rect 422466 170938 422702 171174
rect 422786 170938 423022 171174
rect 422466 170618 422702 170854
rect 422786 170618 423022 170854
rect 422466 152938 422702 153174
rect 422786 152938 423022 153174
rect 422466 152618 422702 152854
rect 422786 152618 423022 152854
rect 422466 134938 422702 135174
rect 422786 134938 423022 135174
rect 422466 134618 422702 134854
rect 422786 134618 423022 134854
rect 422466 116938 422702 117174
rect 422786 116938 423022 117174
rect 422466 116618 422702 116854
rect 422786 116618 423022 116854
rect 422466 98938 422702 99174
rect 422786 98938 423022 99174
rect 422466 98618 422702 98854
rect 422786 98618 423022 98854
rect 422466 80938 422702 81174
rect 422786 80938 423022 81174
rect 422466 80618 422702 80854
rect 422786 80618 423022 80854
rect 422466 62938 422702 63174
rect 422786 62938 423022 63174
rect 422466 62618 422702 62854
rect 422786 62618 423022 62854
rect 422466 44938 422702 45174
rect 422786 44938 423022 45174
rect 422466 44618 422702 44854
rect 422786 44618 423022 44854
rect 422466 26938 422702 27174
rect 422786 26938 423022 27174
rect 422466 26618 422702 26854
rect 422786 26618 423022 26854
rect 422466 8938 422702 9174
rect 422786 8938 423022 9174
rect 422466 8618 422702 8854
rect 422786 8618 423022 8854
rect 422466 -2052 422702 -1816
rect 422786 -2052 423022 -1816
rect 422466 -2372 422702 -2136
rect 422786 -2372 423022 -2136
rect 426186 462776 426422 463012
rect 426506 462776 426742 463012
rect 426186 462456 426422 462692
rect 426506 462456 426742 462692
rect 426186 444658 426422 444894
rect 426506 444658 426742 444894
rect 426186 444338 426422 444574
rect 426506 444338 426742 444574
rect 426186 426658 426422 426894
rect 426506 426658 426742 426894
rect 426186 426338 426422 426574
rect 426506 426338 426742 426574
rect 426186 408658 426422 408894
rect 426506 408658 426742 408894
rect 426186 408338 426422 408574
rect 426506 408338 426742 408574
rect 426186 390658 426422 390894
rect 426506 390658 426742 390894
rect 426186 390338 426422 390574
rect 426506 390338 426742 390574
rect 426186 372658 426422 372894
rect 426506 372658 426742 372894
rect 426186 372338 426422 372574
rect 426506 372338 426742 372574
rect 426186 354658 426422 354894
rect 426506 354658 426742 354894
rect 426186 354338 426422 354574
rect 426506 354338 426742 354574
rect 426186 336658 426422 336894
rect 426506 336658 426742 336894
rect 426186 336338 426422 336574
rect 426506 336338 426742 336574
rect 426186 318658 426422 318894
rect 426506 318658 426742 318894
rect 426186 318338 426422 318574
rect 426506 318338 426742 318574
rect 426186 300658 426422 300894
rect 426506 300658 426742 300894
rect 426186 300338 426422 300574
rect 426506 300338 426742 300574
rect 426186 282658 426422 282894
rect 426506 282658 426742 282894
rect 426186 282338 426422 282574
rect 426506 282338 426742 282574
rect 426186 264658 426422 264894
rect 426506 264658 426742 264894
rect 426186 264338 426422 264574
rect 426506 264338 426742 264574
rect 426186 246658 426422 246894
rect 426506 246658 426742 246894
rect 426186 246338 426422 246574
rect 426506 246338 426742 246574
rect 426186 228658 426422 228894
rect 426506 228658 426742 228894
rect 426186 228338 426422 228574
rect 426506 228338 426742 228574
rect 426186 210658 426422 210894
rect 426506 210658 426742 210894
rect 426186 210338 426422 210574
rect 426506 210338 426742 210574
rect 426186 192658 426422 192894
rect 426506 192658 426742 192894
rect 426186 192338 426422 192574
rect 426506 192338 426742 192574
rect 426186 174658 426422 174894
rect 426506 174658 426742 174894
rect 426186 174338 426422 174574
rect 426506 174338 426742 174574
rect 426186 156658 426422 156894
rect 426506 156658 426742 156894
rect 426186 156338 426422 156574
rect 426506 156338 426742 156574
rect 426186 138658 426422 138894
rect 426506 138658 426742 138894
rect 426186 138338 426422 138574
rect 426506 138338 426742 138574
rect 426186 120658 426422 120894
rect 426506 120658 426742 120894
rect 426186 120338 426422 120574
rect 426506 120338 426742 120574
rect 426186 102658 426422 102894
rect 426506 102658 426742 102894
rect 426186 102338 426422 102574
rect 426506 102338 426742 102574
rect 426186 84658 426422 84894
rect 426506 84658 426742 84894
rect 426186 84338 426422 84574
rect 426506 84338 426742 84574
rect 426186 66658 426422 66894
rect 426506 66658 426742 66894
rect 426186 66338 426422 66574
rect 426506 66338 426742 66574
rect 426186 48658 426422 48894
rect 426506 48658 426742 48894
rect 426186 48338 426422 48574
rect 426506 48338 426742 48574
rect 426186 30658 426422 30894
rect 426506 30658 426742 30894
rect 426186 30338 426422 30574
rect 426506 30338 426742 30574
rect 426186 12658 426422 12894
rect 426506 12658 426742 12894
rect 426186 12338 426422 12574
rect 426506 12338 426742 12574
rect 426186 -3012 426422 -2776
rect 426506 -3012 426742 -2776
rect 426186 -3332 426422 -3096
rect 426506 -3332 426742 -3096
rect 429906 463736 430142 463972
rect 430226 463736 430462 463972
rect 429906 463416 430142 463652
rect 430226 463416 430462 463652
rect 429906 448378 430142 448614
rect 430226 448378 430462 448614
rect 429906 448058 430142 448294
rect 430226 448058 430462 448294
rect 429906 430378 430142 430614
rect 430226 430378 430462 430614
rect 429906 430058 430142 430294
rect 430226 430058 430462 430294
rect 429906 412378 430142 412614
rect 430226 412378 430462 412614
rect 429906 412058 430142 412294
rect 430226 412058 430462 412294
rect 429906 394378 430142 394614
rect 430226 394378 430462 394614
rect 429906 394058 430142 394294
rect 430226 394058 430462 394294
rect 429906 376378 430142 376614
rect 430226 376378 430462 376614
rect 429906 376058 430142 376294
rect 430226 376058 430462 376294
rect 429906 358378 430142 358614
rect 430226 358378 430462 358614
rect 429906 358058 430142 358294
rect 430226 358058 430462 358294
rect 429906 340378 430142 340614
rect 430226 340378 430462 340614
rect 429906 340058 430142 340294
rect 430226 340058 430462 340294
rect 429906 322378 430142 322614
rect 430226 322378 430462 322614
rect 429906 322058 430142 322294
rect 430226 322058 430462 322294
rect 429906 304378 430142 304614
rect 430226 304378 430462 304614
rect 429906 304058 430142 304294
rect 430226 304058 430462 304294
rect 429906 286378 430142 286614
rect 430226 286378 430462 286614
rect 429906 286058 430142 286294
rect 430226 286058 430462 286294
rect 429906 268378 430142 268614
rect 430226 268378 430462 268614
rect 429906 268058 430142 268294
rect 430226 268058 430462 268294
rect 429906 250378 430142 250614
rect 430226 250378 430462 250614
rect 429906 250058 430142 250294
rect 430226 250058 430462 250294
rect 429906 232378 430142 232614
rect 430226 232378 430462 232614
rect 429906 232058 430142 232294
rect 430226 232058 430462 232294
rect 429906 214378 430142 214614
rect 430226 214378 430462 214614
rect 429906 214058 430142 214294
rect 430226 214058 430462 214294
rect 429906 196378 430142 196614
rect 430226 196378 430462 196614
rect 429906 196058 430142 196294
rect 430226 196058 430462 196294
rect 429906 178378 430142 178614
rect 430226 178378 430462 178614
rect 429906 178058 430142 178294
rect 430226 178058 430462 178294
rect 429906 160378 430142 160614
rect 430226 160378 430462 160614
rect 429906 160058 430142 160294
rect 430226 160058 430462 160294
rect 429906 142378 430142 142614
rect 430226 142378 430462 142614
rect 429906 142058 430142 142294
rect 430226 142058 430462 142294
rect 429906 124378 430142 124614
rect 430226 124378 430462 124614
rect 429906 124058 430142 124294
rect 430226 124058 430462 124294
rect 429906 106378 430142 106614
rect 430226 106378 430462 106614
rect 429906 106058 430142 106294
rect 430226 106058 430462 106294
rect 429906 88378 430142 88614
rect 430226 88378 430462 88614
rect 429906 88058 430142 88294
rect 430226 88058 430462 88294
rect 429906 70378 430142 70614
rect 430226 70378 430462 70614
rect 429906 70058 430142 70294
rect 430226 70058 430462 70294
rect 429906 52378 430142 52614
rect 430226 52378 430462 52614
rect 429906 52058 430142 52294
rect 430226 52058 430462 52294
rect 429906 34378 430142 34614
rect 430226 34378 430462 34614
rect 429906 34058 430142 34294
rect 430226 34058 430462 34294
rect 429906 16378 430142 16614
rect 430226 16378 430462 16614
rect 429906 16058 430142 16294
rect 430226 16058 430462 16294
rect 429906 -3972 430142 -3736
rect 430226 -3972 430462 -3736
rect 429906 -4292 430142 -4056
rect 430226 -4292 430462 -4056
rect 436746 460856 436982 461092
rect 437066 460856 437302 461092
rect 436746 460536 436982 460772
rect 437066 460536 437302 460772
rect 436746 455218 436982 455454
rect 437066 455218 437302 455454
rect 436746 454898 436982 455134
rect 437066 454898 437302 455134
rect 436746 437218 436982 437454
rect 437066 437218 437302 437454
rect 436746 436898 436982 437134
rect 437066 436898 437302 437134
rect 436746 419218 436982 419454
rect 437066 419218 437302 419454
rect 436746 418898 436982 419134
rect 437066 418898 437302 419134
rect 436746 401218 436982 401454
rect 437066 401218 437302 401454
rect 436746 400898 436982 401134
rect 437066 400898 437302 401134
rect 436746 383218 436982 383454
rect 437066 383218 437302 383454
rect 436746 382898 436982 383134
rect 437066 382898 437302 383134
rect 436746 365218 436982 365454
rect 437066 365218 437302 365454
rect 436746 364898 436982 365134
rect 437066 364898 437302 365134
rect 436746 347218 436982 347454
rect 437066 347218 437302 347454
rect 436746 346898 436982 347134
rect 437066 346898 437302 347134
rect 436746 329218 436982 329454
rect 437066 329218 437302 329454
rect 436746 328898 436982 329134
rect 437066 328898 437302 329134
rect 436746 311218 436982 311454
rect 437066 311218 437302 311454
rect 436746 310898 436982 311134
rect 437066 310898 437302 311134
rect 436746 293218 436982 293454
rect 437066 293218 437302 293454
rect 436746 292898 436982 293134
rect 437066 292898 437302 293134
rect 436746 275218 436982 275454
rect 437066 275218 437302 275454
rect 436746 274898 436982 275134
rect 437066 274898 437302 275134
rect 436746 257218 436982 257454
rect 437066 257218 437302 257454
rect 436746 256898 436982 257134
rect 437066 256898 437302 257134
rect 436746 239218 436982 239454
rect 437066 239218 437302 239454
rect 436746 238898 436982 239134
rect 437066 238898 437302 239134
rect 436746 221218 436982 221454
rect 437066 221218 437302 221454
rect 436746 220898 436982 221134
rect 437066 220898 437302 221134
rect 436746 203218 436982 203454
rect 437066 203218 437302 203454
rect 436746 202898 436982 203134
rect 437066 202898 437302 203134
rect 436746 185218 436982 185454
rect 437066 185218 437302 185454
rect 436746 184898 436982 185134
rect 437066 184898 437302 185134
rect 436746 167218 436982 167454
rect 437066 167218 437302 167454
rect 436746 166898 436982 167134
rect 437066 166898 437302 167134
rect 436746 149218 436982 149454
rect 437066 149218 437302 149454
rect 436746 148898 436982 149134
rect 437066 148898 437302 149134
rect 436746 131218 436982 131454
rect 437066 131218 437302 131454
rect 436746 130898 436982 131134
rect 437066 130898 437302 131134
rect 436746 113218 436982 113454
rect 437066 113218 437302 113454
rect 436746 112898 436982 113134
rect 437066 112898 437302 113134
rect 436746 95218 436982 95454
rect 437066 95218 437302 95454
rect 436746 94898 436982 95134
rect 437066 94898 437302 95134
rect 436746 77218 436982 77454
rect 437066 77218 437302 77454
rect 436746 76898 436982 77134
rect 437066 76898 437302 77134
rect 436746 59218 436982 59454
rect 437066 59218 437302 59454
rect 436746 58898 436982 59134
rect 437066 58898 437302 59134
rect 436746 41218 436982 41454
rect 437066 41218 437302 41454
rect 436746 40898 436982 41134
rect 437066 40898 437302 41134
rect 436746 23218 436982 23454
rect 437066 23218 437302 23454
rect 436746 22898 436982 23134
rect 437066 22898 437302 23134
rect 436746 5218 436982 5454
rect 437066 5218 437302 5454
rect 436746 4898 436982 5134
rect 437066 4898 437302 5134
rect 436746 -1092 436982 -856
rect 437066 -1092 437302 -856
rect 436746 -1412 436982 -1176
rect 437066 -1412 437302 -1176
rect 440466 461816 440702 462052
rect 440786 461816 441022 462052
rect 440466 461496 440702 461732
rect 440786 461496 441022 461732
rect 440466 440938 440702 441174
rect 440786 440938 441022 441174
rect 440466 440618 440702 440854
rect 440786 440618 441022 440854
rect 440466 422938 440702 423174
rect 440786 422938 441022 423174
rect 440466 422618 440702 422854
rect 440786 422618 441022 422854
rect 440466 404938 440702 405174
rect 440786 404938 441022 405174
rect 440466 404618 440702 404854
rect 440786 404618 441022 404854
rect 440466 386938 440702 387174
rect 440786 386938 441022 387174
rect 440466 386618 440702 386854
rect 440786 386618 441022 386854
rect 440466 368938 440702 369174
rect 440786 368938 441022 369174
rect 440466 368618 440702 368854
rect 440786 368618 441022 368854
rect 440466 350938 440702 351174
rect 440786 350938 441022 351174
rect 440466 350618 440702 350854
rect 440786 350618 441022 350854
rect 440466 332938 440702 333174
rect 440786 332938 441022 333174
rect 440466 332618 440702 332854
rect 440786 332618 441022 332854
rect 440466 314938 440702 315174
rect 440786 314938 441022 315174
rect 440466 314618 440702 314854
rect 440786 314618 441022 314854
rect 440466 296938 440702 297174
rect 440786 296938 441022 297174
rect 440466 296618 440702 296854
rect 440786 296618 441022 296854
rect 440466 278938 440702 279174
rect 440786 278938 441022 279174
rect 440466 278618 440702 278854
rect 440786 278618 441022 278854
rect 440466 260938 440702 261174
rect 440786 260938 441022 261174
rect 440466 260618 440702 260854
rect 440786 260618 441022 260854
rect 440466 242938 440702 243174
rect 440786 242938 441022 243174
rect 440466 242618 440702 242854
rect 440786 242618 441022 242854
rect 440466 224938 440702 225174
rect 440786 224938 441022 225174
rect 440466 224618 440702 224854
rect 440786 224618 441022 224854
rect 440466 206938 440702 207174
rect 440786 206938 441022 207174
rect 440466 206618 440702 206854
rect 440786 206618 441022 206854
rect 440466 188938 440702 189174
rect 440786 188938 441022 189174
rect 440466 188618 440702 188854
rect 440786 188618 441022 188854
rect 440466 170938 440702 171174
rect 440786 170938 441022 171174
rect 440466 170618 440702 170854
rect 440786 170618 441022 170854
rect 440466 152938 440702 153174
rect 440786 152938 441022 153174
rect 440466 152618 440702 152854
rect 440786 152618 441022 152854
rect 440466 134938 440702 135174
rect 440786 134938 441022 135174
rect 440466 134618 440702 134854
rect 440786 134618 441022 134854
rect 440466 116938 440702 117174
rect 440786 116938 441022 117174
rect 440466 116618 440702 116854
rect 440786 116618 441022 116854
rect 440466 98938 440702 99174
rect 440786 98938 441022 99174
rect 440466 98618 440702 98854
rect 440786 98618 441022 98854
rect 440466 80938 440702 81174
rect 440786 80938 441022 81174
rect 440466 80618 440702 80854
rect 440786 80618 441022 80854
rect 440466 62938 440702 63174
rect 440786 62938 441022 63174
rect 440466 62618 440702 62854
rect 440786 62618 441022 62854
rect 440466 44938 440702 45174
rect 440786 44938 441022 45174
rect 440466 44618 440702 44854
rect 440786 44618 441022 44854
rect 440466 26938 440702 27174
rect 440786 26938 441022 27174
rect 440466 26618 440702 26854
rect 440786 26618 441022 26854
rect 440466 8938 440702 9174
rect 440786 8938 441022 9174
rect 440466 8618 440702 8854
rect 440786 8618 441022 8854
rect 440466 -2052 440702 -1816
rect 440786 -2052 441022 -1816
rect 440466 -2372 440702 -2136
rect 440786 -2372 441022 -2136
rect 444186 462776 444422 463012
rect 444506 462776 444742 463012
rect 444186 462456 444422 462692
rect 444506 462456 444742 462692
rect 444186 444658 444422 444894
rect 444506 444658 444742 444894
rect 444186 444338 444422 444574
rect 444506 444338 444742 444574
rect 444186 426658 444422 426894
rect 444506 426658 444742 426894
rect 444186 426338 444422 426574
rect 444506 426338 444742 426574
rect 444186 408658 444422 408894
rect 444506 408658 444742 408894
rect 444186 408338 444422 408574
rect 444506 408338 444742 408574
rect 444186 390658 444422 390894
rect 444506 390658 444742 390894
rect 444186 390338 444422 390574
rect 444506 390338 444742 390574
rect 444186 372658 444422 372894
rect 444506 372658 444742 372894
rect 444186 372338 444422 372574
rect 444506 372338 444742 372574
rect 444186 354658 444422 354894
rect 444506 354658 444742 354894
rect 444186 354338 444422 354574
rect 444506 354338 444742 354574
rect 444186 336658 444422 336894
rect 444506 336658 444742 336894
rect 444186 336338 444422 336574
rect 444506 336338 444742 336574
rect 444186 318658 444422 318894
rect 444506 318658 444742 318894
rect 444186 318338 444422 318574
rect 444506 318338 444742 318574
rect 444186 300658 444422 300894
rect 444506 300658 444742 300894
rect 444186 300338 444422 300574
rect 444506 300338 444742 300574
rect 444186 282658 444422 282894
rect 444506 282658 444742 282894
rect 444186 282338 444422 282574
rect 444506 282338 444742 282574
rect 444186 264658 444422 264894
rect 444506 264658 444742 264894
rect 444186 264338 444422 264574
rect 444506 264338 444742 264574
rect 444186 246658 444422 246894
rect 444506 246658 444742 246894
rect 444186 246338 444422 246574
rect 444506 246338 444742 246574
rect 444186 228658 444422 228894
rect 444506 228658 444742 228894
rect 444186 228338 444422 228574
rect 444506 228338 444742 228574
rect 444186 210658 444422 210894
rect 444506 210658 444742 210894
rect 444186 210338 444422 210574
rect 444506 210338 444742 210574
rect 444186 192658 444422 192894
rect 444506 192658 444742 192894
rect 444186 192338 444422 192574
rect 444506 192338 444742 192574
rect 444186 174658 444422 174894
rect 444506 174658 444742 174894
rect 444186 174338 444422 174574
rect 444506 174338 444742 174574
rect 444186 156658 444422 156894
rect 444506 156658 444742 156894
rect 444186 156338 444422 156574
rect 444506 156338 444742 156574
rect 444186 138658 444422 138894
rect 444506 138658 444742 138894
rect 444186 138338 444422 138574
rect 444506 138338 444742 138574
rect 444186 120658 444422 120894
rect 444506 120658 444742 120894
rect 444186 120338 444422 120574
rect 444506 120338 444742 120574
rect 444186 102658 444422 102894
rect 444506 102658 444742 102894
rect 444186 102338 444422 102574
rect 444506 102338 444742 102574
rect 444186 84658 444422 84894
rect 444506 84658 444742 84894
rect 444186 84338 444422 84574
rect 444506 84338 444742 84574
rect 444186 66658 444422 66894
rect 444506 66658 444742 66894
rect 444186 66338 444422 66574
rect 444506 66338 444742 66574
rect 444186 48658 444422 48894
rect 444506 48658 444742 48894
rect 444186 48338 444422 48574
rect 444506 48338 444742 48574
rect 444186 30658 444422 30894
rect 444506 30658 444742 30894
rect 444186 30338 444422 30574
rect 444506 30338 444742 30574
rect 444186 12658 444422 12894
rect 444506 12658 444742 12894
rect 444186 12338 444422 12574
rect 444506 12338 444742 12574
rect 444186 -3012 444422 -2776
rect 444506 -3012 444742 -2776
rect 444186 -3332 444422 -3096
rect 444506 -3332 444742 -3096
rect 447906 463736 448142 463972
rect 448226 463736 448462 463972
rect 447906 463416 448142 463652
rect 448226 463416 448462 463652
rect 447906 448378 448142 448614
rect 448226 448378 448462 448614
rect 447906 448058 448142 448294
rect 448226 448058 448462 448294
rect 447906 430378 448142 430614
rect 448226 430378 448462 430614
rect 447906 430058 448142 430294
rect 448226 430058 448462 430294
rect 447906 412378 448142 412614
rect 448226 412378 448462 412614
rect 447906 412058 448142 412294
rect 448226 412058 448462 412294
rect 447906 394378 448142 394614
rect 448226 394378 448462 394614
rect 447906 394058 448142 394294
rect 448226 394058 448462 394294
rect 447906 376378 448142 376614
rect 448226 376378 448462 376614
rect 447906 376058 448142 376294
rect 448226 376058 448462 376294
rect 447906 358378 448142 358614
rect 448226 358378 448462 358614
rect 447906 358058 448142 358294
rect 448226 358058 448462 358294
rect 447906 340378 448142 340614
rect 448226 340378 448462 340614
rect 447906 340058 448142 340294
rect 448226 340058 448462 340294
rect 447906 322378 448142 322614
rect 448226 322378 448462 322614
rect 447906 322058 448142 322294
rect 448226 322058 448462 322294
rect 447906 304378 448142 304614
rect 448226 304378 448462 304614
rect 447906 304058 448142 304294
rect 448226 304058 448462 304294
rect 447906 286378 448142 286614
rect 448226 286378 448462 286614
rect 447906 286058 448142 286294
rect 448226 286058 448462 286294
rect 447906 268378 448142 268614
rect 448226 268378 448462 268614
rect 447906 268058 448142 268294
rect 448226 268058 448462 268294
rect 447906 250378 448142 250614
rect 448226 250378 448462 250614
rect 447906 250058 448142 250294
rect 448226 250058 448462 250294
rect 447906 232378 448142 232614
rect 448226 232378 448462 232614
rect 447906 232058 448142 232294
rect 448226 232058 448462 232294
rect 447906 214378 448142 214614
rect 448226 214378 448462 214614
rect 447906 214058 448142 214294
rect 448226 214058 448462 214294
rect 447906 196378 448142 196614
rect 448226 196378 448462 196614
rect 447906 196058 448142 196294
rect 448226 196058 448462 196294
rect 447906 178378 448142 178614
rect 448226 178378 448462 178614
rect 447906 178058 448142 178294
rect 448226 178058 448462 178294
rect 447906 160378 448142 160614
rect 448226 160378 448462 160614
rect 447906 160058 448142 160294
rect 448226 160058 448462 160294
rect 447906 142378 448142 142614
rect 448226 142378 448462 142614
rect 447906 142058 448142 142294
rect 448226 142058 448462 142294
rect 447906 124378 448142 124614
rect 448226 124378 448462 124614
rect 447906 124058 448142 124294
rect 448226 124058 448462 124294
rect 447906 106378 448142 106614
rect 448226 106378 448462 106614
rect 447906 106058 448142 106294
rect 448226 106058 448462 106294
rect 447906 88378 448142 88614
rect 448226 88378 448462 88614
rect 447906 88058 448142 88294
rect 448226 88058 448462 88294
rect 447906 70378 448142 70614
rect 448226 70378 448462 70614
rect 447906 70058 448142 70294
rect 448226 70058 448462 70294
rect 447906 52378 448142 52614
rect 448226 52378 448462 52614
rect 447906 52058 448142 52294
rect 448226 52058 448462 52294
rect 447906 34378 448142 34614
rect 448226 34378 448462 34614
rect 447906 34058 448142 34294
rect 448226 34058 448462 34294
rect 447906 16378 448142 16614
rect 448226 16378 448462 16614
rect 447906 16058 448142 16294
rect 448226 16058 448462 16294
rect 447906 -3972 448142 -3736
rect 448226 -3972 448462 -3736
rect 447906 -4292 448142 -4056
rect 448226 -4292 448462 -4056
rect 454746 460856 454982 461092
rect 455066 460856 455302 461092
rect 454746 460536 454982 460772
rect 455066 460536 455302 460772
rect 454746 455218 454982 455454
rect 455066 455218 455302 455454
rect 454746 454898 454982 455134
rect 455066 454898 455302 455134
rect 454746 437218 454982 437454
rect 455066 437218 455302 437454
rect 454746 436898 454982 437134
rect 455066 436898 455302 437134
rect 454746 419218 454982 419454
rect 455066 419218 455302 419454
rect 454746 418898 454982 419134
rect 455066 418898 455302 419134
rect 454746 401218 454982 401454
rect 455066 401218 455302 401454
rect 454746 400898 454982 401134
rect 455066 400898 455302 401134
rect 454746 383218 454982 383454
rect 455066 383218 455302 383454
rect 454746 382898 454982 383134
rect 455066 382898 455302 383134
rect 454746 365218 454982 365454
rect 455066 365218 455302 365454
rect 454746 364898 454982 365134
rect 455066 364898 455302 365134
rect 454746 347218 454982 347454
rect 455066 347218 455302 347454
rect 454746 346898 454982 347134
rect 455066 346898 455302 347134
rect 454746 329218 454982 329454
rect 455066 329218 455302 329454
rect 454746 328898 454982 329134
rect 455066 328898 455302 329134
rect 454746 311218 454982 311454
rect 455066 311218 455302 311454
rect 454746 310898 454982 311134
rect 455066 310898 455302 311134
rect 454746 293218 454982 293454
rect 455066 293218 455302 293454
rect 454746 292898 454982 293134
rect 455066 292898 455302 293134
rect 454746 275218 454982 275454
rect 455066 275218 455302 275454
rect 454746 274898 454982 275134
rect 455066 274898 455302 275134
rect 454746 257218 454982 257454
rect 455066 257218 455302 257454
rect 454746 256898 454982 257134
rect 455066 256898 455302 257134
rect 454746 239218 454982 239454
rect 455066 239218 455302 239454
rect 454746 238898 454982 239134
rect 455066 238898 455302 239134
rect 454746 221218 454982 221454
rect 455066 221218 455302 221454
rect 454746 220898 454982 221134
rect 455066 220898 455302 221134
rect 454746 203218 454982 203454
rect 455066 203218 455302 203454
rect 454746 202898 454982 203134
rect 455066 202898 455302 203134
rect 454746 185218 454982 185454
rect 455066 185218 455302 185454
rect 454746 184898 454982 185134
rect 455066 184898 455302 185134
rect 454746 167218 454982 167454
rect 455066 167218 455302 167454
rect 454746 166898 454982 167134
rect 455066 166898 455302 167134
rect 454746 149218 454982 149454
rect 455066 149218 455302 149454
rect 454746 148898 454982 149134
rect 455066 148898 455302 149134
rect 454746 131218 454982 131454
rect 455066 131218 455302 131454
rect 454746 130898 454982 131134
rect 455066 130898 455302 131134
rect 454746 113218 454982 113454
rect 455066 113218 455302 113454
rect 454746 112898 454982 113134
rect 455066 112898 455302 113134
rect 454746 95218 454982 95454
rect 455066 95218 455302 95454
rect 454746 94898 454982 95134
rect 455066 94898 455302 95134
rect 454746 77218 454982 77454
rect 455066 77218 455302 77454
rect 454746 76898 454982 77134
rect 455066 76898 455302 77134
rect 454746 59218 454982 59454
rect 455066 59218 455302 59454
rect 454746 58898 454982 59134
rect 455066 58898 455302 59134
rect 454746 41218 454982 41454
rect 455066 41218 455302 41454
rect 454746 40898 454982 41134
rect 455066 40898 455302 41134
rect 454746 23218 454982 23454
rect 455066 23218 455302 23454
rect 454746 22898 454982 23134
rect 455066 22898 455302 23134
rect 454746 5218 454982 5454
rect 455066 5218 455302 5454
rect 454746 4898 454982 5134
rect 455066 4898 455302 5134
rect 454746 -1092 454982 -856
rect 455066 -1092 455302 -856
rect 454746 -1412 454982 -1176
rect 455066 -1412 455302 -1176
rect 458466 461816 458702 462052
rect 458786 461816 459022 462052
rect 458466 461496 458702 461732
rect 458786 461496 459022 461732
rect 458466 440938 458702 441174
rect 458786 440938 459022 441174
rect 458466 440618 458702 440854
rect 458786 440618 459022 440854
rect 458466 422938 458702 423174
rect 458786 422938 459022 423174
rect 458466 422618 458702 422854
rect 458786 422618 459022 422854
rect 458466 404938 458702 405174
rect 458786 404938 459022 405174
rect 458466 404618 458702 404854
rect 458786 404618 459022 404854
rect 458466 386938 458702 387174
rect 458786 386938 459022 387174
rect 458466 386618 458702 386854
rect 458786 386618 459022 386854
rect 458466 368938 458702 369174
rect 458786 368938 459022 369174
rect 458466 368618 458702 368854
rect 458786 368618 459022 368854
rect 458466 350938 458702 351174
rect 458786 350938 459022 351174
rect 458466 350618 458702 350854
rect 458786 350618 459022 350854
rect 458466 332938 458702 333174
rect 458786 332938 459022 333174
rect 458466 332618 458702 332854
rect 458786 332618 459022 332854
rect 458466 314938 458702 315174
rect 458786 314938 459022 315174
rect 458466 314618 458702 314854
rect 458786 314618 459022 314854
rect 458466 296938 458702 297174
rect 458786 296938 459022 297174
rect 458466 296618 458702 296854
rect 458786 296618 459022 296854
rect 458466 278938 458702 279174
rect 458786 278938 459022 279174
rect 458466 278618 458702 278854
rect 458786 278618 459022 278854
rect 458466 260938 458702 261174
rect 458786 260938 459022 261174
rect 458466 260618 458702 260854
rect 458786 260618 459022 260854
rect 458466 242938 458702 243174
rect 458786 242938 459022 243174
rect 458466 242618 458702 242854
rect 458786 242618 459022 242854
rect 458466 224938 458702 225174
rect 458786 224938 459022 225174
rect 458466 224618 458702 224854
rect 458786 224618 459022 224854
rect 458466 206938 458702 207174
rect 458786 206938 459022 207174
rect 458466 206618 458702 206854
rect 458786 206618 459022 206854
rect 458466 188938 458702 189174
rect 458786 188938 459022 189174
rect 458466 188618 458702 188854
rect 458786 188618 459022 188854
rect 458466 170938 458702 171174
rect 458786 170938 459022 171174
rect 458466 170618 458702 170854
rect 458786 170618 459022 170854
rect 458466 152938 458702 153174
rect 458786 152938 459022 153174
rect 458466 152618 458702 152854
rect 458786 152618 459022 152854
rect 458466 134938 458702 135174
rect 458786 134938 459022 135174
rect 458466 134618 458702 134854
rect 458786 134618 459022 134854
rect 458466 116938 458702 117174
rect 458786 116938 459022 117174
rect 458466 116618 458702 116854
rect 458786 116618 459022 116854
rect 458466 98938 458702 99174
rect 458786 98938 459022 99174
rect 458466 98618 458702 98854
rect 458786 98618 459022 98854
rect 458466 80938 458702 81174
rect 458786 80938 459022 81174
rect 458466 80618 458702 80854
rect 458786 80618 459022 80854
rect 458466 62938 458702 63174
rect 458786 62938 459022 63174
rect 458466 62618 458702 62854
rect 458786 62618 459022 62854
rect 458466 44938 458702 45174
rect 458786 44938 459022 45174
rect 458466 44618 458702 44854
rect 458786 44618 459022 44854
rect 458466 26938 458702 27174
rect 458786 26938 459022 27174
rect 458466 26618 458702 26854
rect 458786 26618 459022 26854
rect 458466 8938 458702 9174
rect 458786 8938 459022 9174
rect 458466 8618 458702 8854
rect 458786 8618 459022 8854
rect 458466 -2052 458702 -1816
rect 458786 -2052 459022 -1816
rect 458466 -2372 458702 -2136
rect 458786 -2372 459022 -2136
rect 462186 462776 462422 463012
rect 462506 462776 462742 463012
rect 462186 462456 462422 462692
rect 462506 462456 462742 462692
rect 462186 444658 462422 444894
rect 462506 444658 462742 444894
rect 462186 444338 462422 444574
rect 462506 444338 462742 444574
rect 462186 426658 462422 426894
rect 462506 426658 462742 426894
rect 462186 426338 462422 426574
rect 462506 426338 462742 426574
rect 462186 408658 462422 408894
rect 462506 408658 462742 408894
rect 462186 408338 462422 408574
rect 462506 408338 462742 408574
rect 462186 390658 462422 390894
rect 462506 390658 462742 390894
rect 462186 390338 462422 390574
rect 462506 390338 462742 390574
rect 462186 372658 462422 372894
rect 462506 372658 462742 372894
rect 462186 372338 462422 372574
rect 462506 372338 462742 372574
rect 462186 354658 462422 354894
rect 462506 354658 462742 354894
rect 462186 354338 462422 354574
rect 462506 354338 462742 354574
rect 462186 336658 462422 336894
rect 462506 336658 462742 336894
rect 462186 336338 462422 336574
rect 462506 336338 462742 336574
rect 462186 318658 462422 318894
rect 462506 318658 462742 318894
rect 462186 318338 462422 318574
rect 462506 318338 462742 318574
rect 462186 300658 462422 300894
rect 462506 300658 462742 300894
rect 462186 300338 462422 300574
rect 462506 300338 462742 300574
rect 462186 282658 462422 282894
rect 462506 282658 462742 282894
rect 462186 282338 462422 282574
rect 462506 282338 462742 282574
rect 462186 264658 462422 264894
rect 462506 264658 462742 264894
rect 462186 264338 462422 264574
rect 462506 264338 462742 264574
rect 462186 246658 462422 246894
rect 462506 246658 462742 246894
rect 462186 246338 462422 246574
rect 462506 246338 462742 246574
rect 462186 228658 462422 228894
rect 462506 228658 462742 228894
rect 462186 228338 462422 228574
rect 462506 228338 462742 228574
rect 462186 210658 462422 210894
rect 462506 210658 462742 210894
rect 462186 210338 462422 210574
rect 462506 210338 462742 210574
rect 462186 192658 462422 192894
rect 462506 192658 462742 192894
rect 462186 192338 462422 192574
rect 462506 192338 462742 192574
rect 462186 174658 462422 174894
rect 462506 174658 462742 174894
rect 462186 174338 462422 174574
rect 462506 174338 462742 174574
rect 462186 156658 462422 156894
rect 462506 156658 462742 156894
rect 462186 156338 462422 156574
rect 462506 156338 462742 156574
rect 462186 138658 462422 138894
rect 462506 138658 462742 138894
rect 462186 138338 462422 138574
rect 462506 138338 462742 138574
rect 462186 120658 462422 120894
rect 462506 120658 462742 120894
rect 462186 120338 462422 120574
rect 462506 120338 462742 120574
rect 462186 102658 462422 102894
rect 462506 102658 462742 102894
rect 462186 102338 462422 102574
rect 462506 102338 462742 102574
rect 462186 84658 462422 84894
rect 462506 84658 462742 84894
rect 462186 84338 462422 84574
rect 462506 84338 462742 84574
rect 462186 66658 462422 66894
rect 462506 66658 462742 66894
rect 462186 66338 462422 66574
rect 462506 66338 462742 66574
rect 462186 48658 462422 48894
rect 462506 48658 462742 48894
rect 462186 48338 462422 48574
rect 462506 48338 462742 48574
rect 462186 30658 462422 30894
rect 462506 30658 462742 30894
rect 462186 30338 462422 30574
rect 462506 30338 462742 30574
rect 462186 12658 462422 12894
rect 462506 12658 462742 12894
rect 462186 12338 462422 12574
rect 462506 12338 462742 12574
rect 462186 -3012 462422 -2776
rect 462506 -3012 462742 -2776
rect 462186 -3332 462422 -3096
rect 462506 -3332 462742 -3096
rect 465906 463736 466142 463972
rect 466226 463736 466462 463972
rect 465906 463416 466142 463652
rect 466226 463416 466462 463652
rect 465906 448378 466142 448614
rect 466226 448378 466462 448614
rect 465906 448058 466142 448294
rect 466226 448058 466462 448294
rect 465906 430378 466142 430614
rect 466226 430378 466462 430614
rect 465906 430058 466142 430294
rect 466226 430058 466462 430294
rect 465906 412378 466142 412614
rect 466226 412378 466462 412614
rect 465906 412058 466142 412294
rect 466226 412058 466462 412294
rect 465906 394378 466142 394614
rect 466226 394378 466462 394614
rect 465906 394058 466142 394294
rect 466226 394058 466462 394294
rect 465906 376378 466142 376614
rect 466226 376378 466462 376614
rect 465906 376058 466142 376294
rect 466226 376058 466462 376294
rect 465906 358378 466142 358614
rect 466226 358378 466462 358614
rect 465906 358058 466142 358294
rect 466226 358058 466462 358294
rect 465906 340378 466142 340614
rect 466226 340378 466462 340614
rect 465906 340058 466142 340294
rect 466226 340058 466462 340294
rect 465906 322378 466142 322614
rect 466226 322378 466462 322614
rect 465906 322058 466142 322294
rect 466226 322058 466462 322294
rect 465906 304378 466142 304614
rect 466226 304378 466462 304614
rect 465906 304058 466142 304294
rect 466226 304058 466462 304294
rect 465906 286378 466142 286614
rect 466226 286378 466462 286614
rect 465906 286058 466142 286294
rect 466226 286058 466462 286294
rect 465906 268378 466142 268614
rect 466226 268378 466462 268614
rect 465906 268058 466142 268294
rect 466226 268058 466462 268294
rect 465906 250378 466142 250614
rect 466226 250378 466462 250614
rect 465906 250058 466142 250294
rect 466226 250058 466462 250294
rect 465906 232378 466142 232614
rect 466226 232378 466462 232614
rect 465906 232058 466142 232294
rect 466226 232058 466462 232294
rect 465906 214378 466142 214614
rect 466226 214378 466462 214614
rect 465906 214058 466142 214294
rect 466226 214058 466462 214294
rect 465906 196378 466142 196614
rect 466226 196378 466462 196614
rect 465906 196058 466142 196294
rect 466226 196058 466462 196294
rect 465906 178378 466142 178614
rect 466226 178378 466462 178614
rect 465906 178058 466142 178294
rect 466226 178058 466462 178294
rect 465906 160378 466142 160614
rect 466226 160378 466462 160614
rect 465906 160058 466142 160294
rect 466226 160058 466462 160294
rect 465906 142378 466142 142614
rect 466226 142378 466462 142614
rect 465906 142058 466142 142294
rect 466226 142058 466462 142294
rect 465906 124378 466142 124614
rect 466226 124378 466462 124614
rect 465906 124058 466142 124294
rect 466226 124058 466462 124294
rect 465906 106378 466142 106614
rect 466226 106378 466462 106614
rect 465906 106058 466142 106294
rect 466226 106058 466462 106294
rect 465906 88378 466142 88614
rect 466226 88378 466462 88614
rect 465906 88058 466142 88294
rect 466226 88058 466462 88294
rect 465906 70378 466142 70614
rect 466226 70378 466462 70614
rect 465906 70058 466142 70294
rect 466226 70058 466462 70294
rect 465906 52378 466142 52614
rect 466226 52378 466462 52614
rect 465906 52058 466142 52294
rect 466226 52058 466462 52294
rect 465906 34378 466142 34614
rect 466226 34378 466462 34614
rect 465906 34058 466142 34294
rect 466226 34058 466462 34294
rect 465906 16378 466142 16614
rect 466226 16378 466462 16614
rect 465906 16058 466142 16294
rect 466226 16058 466462 16294
rect 465906 -3972 466142 -3736
rect 466226 -3972 466462 -3736
rect 465906 -4292 466142 -4056
rect 466226 -4292 466462 -4056
rect 472746 460856 472982 461092
rect 473066 460856 473302 461092
rect 472746 460536 472982 460772
rect 473066 460536 473302 460772
rect 472746 455218 472982 455454
rect 473066 455218 473302 455454
rect 472746 454898 472982 455134
rect 473066 454898 473302 455134
rect 472746 437218 472982 437454
rect 473066 437218 473302 437454
rect 472746 436898 472982 437134
rect 473066 436898 473302 437134
rect 472746 419218 472982 419454
rect 473066 419218 473302 419454
rect 472746 418898 472982 419134
rect 473066 418898 473302 419134
rect 472746 401218 472982 401454
rect 473066 401218 473302 401454
rect 472746 400898 472982 401134
rect 473066 400898 473302 401134
rect 472746 383218 472982 383454
rect 473066 383218 473302 383454
rect 472746 382898 472982 383134
rect 473066 382898 473302 383134
rect 472746 365218 472982 365454
rect 473066 365218 473302 365454
rect 472746 364898 472982 365134
rect 473066 364898 473302 365134
rect 472746 347218 472982 347454
rect 473066 347218 473302 347454
rect 472746 346898 472982 347134
rect 473066 346898 473302 347134
rect 472746 329218 472982 329454
rect 473066 329218 473302 329454
rect 472746 328898 472982 329134
rect 473066 328898 473302 329134
rect 472746 311218 472982 311454
rect 473066 311218 473302 311454
rect 472746 310898 472982 311134
rect 473066 310898 473302 311134
rect 472746 293218 472982 293454
rect 473066 293218 473302 293454
rect 472746 292898 472982 293134
rect 473066 292898 473302 293134
rect 472746 275218 472982 275454
rect 473066 275218 473302 275454
rect 472746 274898 472982 275134
rect 473066 274898 473302 275134
rect 472746 257218 472982 257454
rect 473066 257218 473302 257454
rect 472746 256898 472982 257134
rect 473066 256898 473302 257134
rect 472746 239218 472982 239454
rect 473066 239218 473302 239454
rect 472746 238898 472982 239134
rect 473066 238898 473302 239134
rect 472746 221218 472982 221454
rect 473066 221218 473302 221454
rect 472746 220898 472982 221134
rect 473066 220898 473302 221134
rect 472746 203218 472982 203454
rect 473066 203218 473302 203454
rect 472746 202898 472982 203134
rect 473066 202898 473302 203134
rect 472746 185218 472982 185454
rect 473066 185218 473302 185454
rect 472746 184898 472982 185134
rect 473066 184898 473302 185134
rect 472746 167218 472982 167454
rect 473066 167218 473302 167454
rect 472746 166898 472982 167134
rect 473066 166898 473302 167134
rect 472746 149218 472982 149454
rect 473066 149218 473302 149454
rect 472746 148898 472982 149134
rect 473066 148898 473302 149134
rect 472746 131218 472982 131454
rect 473066 131218 473302 131454
rect 472746 130898 472982 131134
rect 473066 130898 473302 131134
rect 472746 113218 472982 113454
rect 473066 113218 473302 113454
rect 472746 112898 472982 113134
rect 473066 112898 473302 113134
rect 472746 95218 472982 95454
rect 473066 95218 473302 95454
rect 472746 94898 472982 95134
rect 473066 94898 473302 95134
rect 472746 77218 472982 77454
rect 473066 77218 473302 77454
rect 472746 76898 472982 77134
rect 473066 76898 473302 77134
rect 472746 59218 472982 59454
rect 473066 59218 473302 59454
rect 472746 58898 472982 59134
rect 473066 58898 473302 59134
rect 472746 41218 472982 41454
rect 473066 41218 473302 41454
rect 472746 40898 472982 41134
rect 473066 40898 473302 41134
rect 472746 23218 472982 23454
rect 473066 23218 473302 23454
rect 472746 22898 472982 23134
rect 473066 22898 473302 23134
rect 472746 5218 472982 5454
rect 473066 5218 473302 5454
rect 472746 4898 472982 5134
rect 473066 4898 473302 5134
rect 472746 -1092 472982 -856
rect 473066 -1092 473302 -856
rect 472746 -1412 472982 -1176
rect 473066 -1412 473302 -1176
rect 476466 461816 476702 462052
rect 476786 461816 477022 462052
rect 476466 461496 476702 461732
rect 476786 461496 477022 461732
rect 476466 440938 476702 441174
rect 476786 440938 477022 441174
rect 476466 440618 476702 440854
rect 476786 440618 477022 440854
rect 476466 422938 476702 423174
rect 476786 422938 477022 423174
rect 476466 422618 476702 422854
rect 476786 422618 477022 422854
rect 476466 404938 476702 405174
rect 476786 404938 477022 405174
rect 476466 404618 476702 404854
rect 476786 404618 477022 404854
rect 476466 386938 476702 387174
rect 476786 386938 477022 387174
rect 476466 386618 476702 386854
rect 476786 386618 477022 386854
rect 476466 368938 476702 369174
rect 476786 368938 477022 369174
rect 476466 368618 476702 368854
rect 476786 368618 477022 368854
rect 476466 350938 476702 351174
rect 476786 350938 477022 351174
rect 476466 350618 476702 350854
rect 476786 350618 477022 350854
rect 476466 332938 476702 333174
rect 476786 332938 477022 333174
rect 476466 332618 476702 332854
rect 476786 332618 477022 332854
rect 476466 314938 476702 315174
rect 476786 314938 477022 315174
rect 476466 314618 476702 314854
rect 476786 314618 477022 314854
rect 476466 296938 476702 297174
rect 476786 296938 477022 297174
rect 476466 296618 476702 296854
rect 476786 296618 477022 296854
rect 476466 278938 476702 279174
rect 476786 278938 477022 279174
rect 476466 278618 476702 278854
rect 476786 278618 477022 278854
rect 476466 260938 476702 261174
rect 476786 260938 477022 261174
rect 476466 260618 476702 260854
rect 476786 260618 477022 260854
rect 476466 242938 476702 243174
rect 476786 242938 477022 243174
rect 476466 242618 476702 242854
rect 476786 242618 477022 242854
rect 476466 224938 476702 225174
rect 476786 224938 477022 225174
rect 476466 224618 476702 224854
rect 476786 224618 477022 224854
rect 476466 206938 476702 207174
rect 476786 206938 477022 207174
rect 476466 206618 476702 206854
rect 476786 206618 477022 206854
rect 476466 188938 476702 189174
rect 476786 188938 477022 189174
rect 476466 188618 476702 188854
rect 476786 188618 477022 188854
rect 476466 170938 476702 171174
rect 476786 170938 477022 171174
rect 476466 170618 476702 170854
rect 476786 170618 477022 170854
rect 476466 152938 476702 153174
rect 476786 152938 477022 153174
rect 476466 152618 476702 152854
rect 476786 152618 477022 152854
rect 476466 134938 476702 135174
rect 476786 134938 477022 135174
rect 476466 134618 476702 134854
rect 476786 134618 477022 134854
rect 476466 116938 476702 117174
rect 476786 116938 477022 117174
rect 476466 116618 476702 116854
rect 476786 116618 477022 116854
rect 476466 98938 476702 99174
rect 476786 98938 477022 99174
rect 476466 98618 476702 98854
rect 476786 98618 477022 98854
rect 476466 80938 476702 81174
rect 476786 80938 477022 81174
rect 476466 80618 476702 80854
rect 476786 80618 477022 80854
rect 476466 62938 476702 63174
rect 476786 62938 477022 63174
rect 476466 62618 476702 62854
rect 476786 62618 477022 62854
rect 476466 44938 476702 45174
rect 476786 44938 477022 45174
rect 476466 44618 476702 44854
rect 476786 44618 477022 44854
rect 476466 26938 476702 27174
rect 476786 26938 477022 27174
rect 476466 26618 476702 26854
rect 476786 26618 477022 26854
rect 476466 8938 476702 9174
rect 476786 8938 477022 9174
rect 476466 8618 476702 8854
rect 476786 8618 477022 8854
rect 476466 -2052 476702 -1816
rect 476786 -2052 477022 -1816
rect 476466 -2372 476702 -2136
rect 476786 -2372 477022 -2136
rect 480186 462776 480422 463012
rect 480506 462776 480742 463012
rect 480186 462456 480422 462692
rect 480506 462456 480742 462692
rect 480186 444658 480422 444894
rect 480506 444658 480742 444894
rect 480186 444338 480422 444574
rect 480506 444338 480742 444574
rect 480186 426658 480422 426894
rect 480506 426658 480742 426894
rect 480186 426338 480422 426574
rect 480506 426338 480742 426574
rect 480186 408658 480422 408894
rect 480506 408658 480742 408894
rect 480186 408338 480422 408574
rect 480506 408338 480742 408574
rect 480186 390658 480422 390894
rect 480506 390658 480742 390894
rect 480186 390338 480422 390574
rect 480506 390338 480742 390574
rect 480186 372658 480422 372894
rect 480506 372658 480742 372894
rect 480186 372338 480422 372574
rect 480506 372338 480742 372574
rect 480186 354658 480422 354894
rect 480506 354658 480742 354894
rect 480186 354338 480422 354574
rect 480506 354338 480742 354574
rect 480186 336658 480422 336894
rect 480506 336658 480742 336894
rect 480186 336338 480422 336574
rect 480506 336338 480742 336574
rect 480186 318658 480422 318894
rect 480506 318658 480742 318894
rect 480186 318338 480422 318574
rect 480506 318338 480742 318574
rect 480186 300658 480422 300894
rect 480506 300658 480742 300894
rect 480186 300338 480422 300574
rect 480506 300338 480742 300574
rect 480186 282658 480422 282894
rect 480506 282658 480742 282894
rect 480186 282338 480422 282574
rect 480506 282338 480742 282574
rect 480186 264658 480422 264894
rect 480506 264658 480742 264894
rect 480186 264338 480422 264574
rect 480506 264338 480742 264574
rect 480186 246658 480422 246894
rect 480506 246658 480742 246894
rect 480186 246338 480422 246574
rect 480506 246338 480742 246574
rect 480186 228658 480422 228894
rect 480506 228658 480742 228894
rect 480186 228338 480422 228574
rect 480506 228338 480742 228574
rect 480186 210658 480422 210894
rect 480506 210658 480742 210894
rect 480186 210338 480422 210574
rect 480506 210338 480742 210574
rect 480186 192658 480422 192894
rect 480506 192658 480742 192894
rect 480186 192338 480422 192574
rect 480506 192338 480742 192574
rect 480186 174658 480422 174894
rect 480506 174658 480742 174894
rect 480186 174338 480422 174574
rect 480506 174338 480742 174574
rect 480186 156658 480422 156894
rect 480506 156658 480742 156894
rect 480186 156338 480422 156574
rect 480506 156338 480742 156574
rect 480186 138658 480422 138894
rect 480506 138658 480742 138894
rect 480186 138338 480422 138574
rect 480506 138338 480742 138574
rect 480186 120658 480422 120894
rect 480506 120658 480742 120894
rect 480186 120338 480422 120574
rect 480506 120338 480742 120574
rect 480186 102658 480422 102894
rect 480506 102658 480742 102894
rect 480186 102338 480422 102574
rect 480506 102338 480742 102574
rect 480186 84658 480422 84894
rect 480506 84658 480742 84894
rect 480186 84338 480422 84574
rect 480506 84338 480742 84574
rect 480186 66658 480422 66894
rect 480506 66658 480742 66894
rect 480186 66338 480422 66574
rect 480506 66338 480742 66574
rect 480186 48658 480422 48894
rect 480506 48658 480742 48894
rect 480186 48338 480422 48574
rect 480506 48338 480742 48574
rect 480186 30658 480422 30894
rect 480506 30658 480742 30894
rect 480186 30338 480422 30574
rect 480506 30338 480742 30574
rect 480186 12658 480422 12894
rect 480506 12658 480742 12894
rect 480186 12338 480422 12574
rect 480506 12338 480742 12574
rect 480186 -3012 480422 -2776
rect 480506 -3012 480742 -2776
rect 480186 -3332 480422 -3096
rect 480506 -3332 480742 -3096
rect 483906 463736 484142 463972
rect 484226 463736 484462 463972
rect 483906 463416 484142 463652
rect 484226 463416 484462 463652
rect 483906 448378 484142 448614
rect 484226 448378 484462 448614
rect 483906 448058 484142 448294
rect 484226 448058 484462 448294
rect 483906 430378 484142 430614
rect 484226 430378 484462 430614
rect 483906 430058 484142 430294
rect 484226 430058 484462 430294
rect 483906 412378 484142 412614
rect 484226 412378 484462 412614
rect 483906 412058 484142 412294
rect 484226 412058 484462 412294
rect 483906 394378 484142 394614
rect 484226 394378 484462 394614
rect 483906 394058 484142 394294
rect 484226 394058 484462 394294
rect 483906 376378 484142 376614
rect 484226 376378 484462 376614
rect 483906 376058 484142 376294
rect 484226 376058 484462 376294
rect 483906 358378 484142 358614
rect 484226 358378 484462 358614
rect 483906 358058 484142 358294
rect 484226 358058 484462 358294
rect 483906 340378 484142 340614
rect 484226 340378 484462 340614
rect 483906 340058 484142 340294
rect 484226 340058 484462 340294
rect 483906 322378 484142 322614
rect 484226 322378 484462 322614
rect 483906 322058 484142 322294
rect 484226 322058 484462 322294
rect 483906 304378 484142 304614
rect 484226 304378 484462 304614
rect 483906 304058 484142 304294
rect 484226 304058 484462 304294
rect 483906 286378 484142 286614
rect 484226 286378 484462 286614
rect 483906 286058 484142 286294
rect 484226 286058 484462 286294
rect 483906 268378 484142 268614
rect 484226 268378 484462 268614
rect 483906 268058 484142 268294
rect 484226 268058 484462 268294
rect 483906 250378 484142 250614
rect 484226 250378 484462 250614
rect 483906 250058 484142 250294
rect 484226 250058 484462 250294
rect 483906 232378 484142 232614
rect 484226 232378 484462 232614
rect 483906 232058 484142 232294
rect 484226 232058 484462 232294
rect 483906 214378 484142 214614
rect 484226 214378 484462 214614
rect 483906 214058 484142 214294
rect 484226 214058 484462 214294
rect 483906 196378 484142 196614
rect 484226 196378 484462 196614
rect 483906 196058 484142 196294
rect 484226 196058 484462 196294
rect 483906 178378 484142 178614
rect 484226 178378 484462 178614
rect 483906 178058 484142 178294
rect 484226 178058 484462 178294
rect 483906 160378 484142 160614
rect 484226 160378 484462 160614
rect 483906 160058 484142 160294
rect 484226 160058 484462 160294
rect 483906 142378 484142 142614
rect 484226 142378 484462 142614
rect 483906 142058 484142 142294
rect 484226 142058 484462 142294
rect 483906 124378 484142 124614
rect 484226 124378 484462 124614
rect 483906 124058 484142 124294
rect 484226 124058 484462 124294
rect 483906 106378 484142 106614
rect 484226 106378 484462 106614
rect 483906 106058 484142 106294
rect 484226 106058 484462 106294
rect 483906 88378 484142 88614
rect 484226 88378 484462 88614
rect 483906 88058 484142 88294
rect 484226 88058 484462 88294
rect 483906 70378 484142 70614
rect 484226 70378 484462 70614
rect 483906 70058 484142 70294
rect 484226 70058 484462 70294
rect 483906 52378 484142 52614
rect 484226 52378 484462 52614
rect 483906 52058 484142 52294
rect 484226 52058 484462 52294
rect 483906 34378 484142 34614
rect 484226 34378 484462 34614
rect 483906 34058 484142 34294
rect 484226 34058 484462 34294
rect 483906 16378 484142 16614
rect 484226 16378 484462 16614
rect 483906 16058 484142 16294
rect 484226 16058 484462 16294
rect 483906 -3972 484142 -3736
rect 484226 -3972 484462 -3736
rect 483906 -4292 484142 -4056
rect 484226 -4292 484462 -4056
rect 490746 460856 490982 461092
rect 491066 460856 491302 461092
rect 490746 460536 490982 460772
rect 491066 460536 491302 460772
rect 490746 455218 490982 455454
rect 491066 455218 491302 455454
rect 490746 454898 490982 455134
rect 491066 454898 491302 455134
rect 490746 437218 490982 437454
rect 491066 437218 491302 437454
rect 490746 436898 490982 437134
rect 491066 436898 491302 437134
rect 490746 419218 490982 419454
rect 491066 419218 491302 419454
rect 490746 418898 490982 419134
rect 491066 418898 491302 419134
rect 490746 401218 490982 401454
rect 491066 401218 491302 401454
rect 490746 400898 490982 401134
rect 491066 400898 491302 401134
rect 490746 383218 490982 383454
rect 491066 383218 491302 383454
rect 490746 382898 490982 383134
rect 491066 382898 491302 383134
rect 490746 365218 490982 365454
rect 491066 365218 491302 365454
rect 490746 364898 490982 365134
rect 491066 364898 491302 365134
rect 490746 347218 490982 347454
rect 491066 347218 491302 347454
rect 490746 346898 490982 347134
rect 491066 346898 491302 347134
rect 490746 329218 490982 329454
rect 491066 329218 491302 329454
rect 490746 328898 490982 329134
rect 491066 328898 491302 329134
rect 490746 311218 490982 311454
rect 491066 311218 491302 311454
rect 490746 310898 490982 311134
rect 491066 310898 491302 311134
rect 490746 293218 490982 293454
rect 491066 293218 491302 293454
rect 490746 292898 490982 293134
rect 491066 292898 491302 293134
rect 490746 275218 490982 275454
rect 491066 275218 491302 275454
rect 490746 274898 490982 275134
rect 491066 274898 491302 275134
rect 490746 257218 490982 257454
rect 491066 257218 491302 257454
rect 490746 256898 490982 257134
rect 491066 256898 491302 257134
rect 490746 239218 490982 239454
rect 491066 239218 491302 239454
rect 490746 238898 490982 239134
rect 491066 238898 491302 239134
rect 490746 221218 490982 221454
rect 491066 221218 491302 221454
rect 490746 220898 490982 221134
rect 491066 220898 491302 221134
rect 490746 203218 490982 203454
rect 491066 203218 491302 203454
rect 490746 202898 490982 203134
rect 491066 202898 491302 203134
rect 490746 185218 490982 185454
rect 491066 185218 491302 185454
rect 490746 184898 490982 185134
rect 491066 184898 491302 185134
rect 490746 167218 490982 167454
rect 491066 167218 491302 167454
rect 490746 166898 490982 167134
rect 491066 166898 491302 167134
rect 490746 149218 490982 149454
rect 491066 149218 491302 149454
rect 490746 148898 490982 149134
rect 491066 148898 491302 149134
rect 490746 131218 490982 131454
rect 491066 131218 491302 131454
rect 490746 130898 490982 131134
rect 491066 130898 491302 131134
rect 490746 113218 490982 113454
rect 491066 113218 491302 113454
rect 490746 112898 490982 113134
rect 491066 112898 491302 113134
rect 490746 95218 490982 95454
rect 491066 95218 491302 95454
rect 490746 94898 490982 95134
rect 491066 94898 491302 95134
rect 490746 77218 490982 77454
rect 491066 77218 491302 77454
rect 490746 76898 490982 77134
rect 491066 76898 491302 77134
rect 490746 59218 490982 59454
rect 491066 59218 491302 59454
rect 490746 58898 490982 59134
rect 491066 58898 491302 59134
rect 490746 41218 490982 41454
rect 491066 41218 491302 41454
rect 490746 40898 490982 41134
rect 491066 40898 491302 41134
rect 490746 23218 490982 23454
rect 491066 23218 491302 23454
rect 490746 22898 490982 23134
rect 491066 22898 491302 23134
rect 490746 5218 490982 5454
rect 491066 5218 491302 5454
rect 490746 4898 490982 5134
rect 491066 4898 491302 5134
rect 490746 -1092 490982 -856
rect 491066 -1092 491302 -856
rect 490746 -1412 490982 -1176
rect 491066 -1412 491302 -1176
rect 494466 461816 494702 462052
rect 494786 461816 495022 462052
rect 494466 461496 494702 461732
rect 494786 461496 495022 461732
rect 494466 440938 494702 441174
rect 494786 440938 495022 441174
rect 494466 440618 494702 440854
rect 494786 440618 495022 440854
rect 494466 422938 494702 423174
rect 494786 422938 495022 423174
rect 494466 422618 494702 422854
rect 494786 422618 495022 422854
rect 494466 404938 494702 405174
rect 494786 404938 495022 405174
rect 494466 404618 494702 404854
rect 494786 404618 495022 404854
rect 494466 386938 494702 387174
rect 494786 386938 495022 387174
rect 494466 386618 494702 386854
rect 494786 386618 495022 386854
rect 494466 368938 494702 369174
rect 494786 368938 495022 369174
rect 494466 368618 494702 368854
rect 494786 368618 495022 368854
rect 494466 350938 494702 351174
rect 494786 350938 495022 351174
rect 494466 350618 494702 350854
rect 494786 350618 495022 350854
rect 494466 332938 494702 333174
rect 494786 332938 495022 333174
rect 494466 332618 494702 332854
rect 494786 332618 495022 332854
rect 494466 314938 494702 315174
rect 494786 314938 495022 315174
rect 494466 314618 494702 314854
rect 494786 314618 495022 314854
rect 494466 296938 494702 297174
rect 494786 296938 495022 297174
rect 494466 296618 494702 296854
rect 494786 296618 495022 296854
rect 494466 278938 494702 279174
rect 494786 278938 495022 279174
rect 494466 278618 494702 278854
rect 494786 278618 495022 278854
rect 494466 260938 494702 261174
rect 494786 260938 495022 261174
rect 494466 260618 494702 260854
rect 494786 260618 495022 260854
rect 494466 242938 494702 243174
rect 494786 242938 495022 243174
rect 494466 242618 494702 242854
rect 494786 242618 495022 242854
rect 494466 224938 494702 225174
rect 494786 224938 495022 225174
rect 494466 224618 494702 224854
rect 494786 224618 495022 224854
rect 494466 206938 494702 207174
rect 494786 206938 495022 207174
rect 494466 206618 494702 206854
rect 494786 206618 495022 206854
rect 494466 188938 494702 189174
rect 494786 188938 495022 189174
rect 494466 188618 494702 188854
rect 494786 188618 495022 188854
rect 494466 170938 494702 171174
rect 494786 170938 495022 171174
rect 494466 170618 494702 170854
rect 494786 170618 495022 170854
rect 494466 152938 494702 153174
rect 494786 152938 495022 153174
rect 494466 152618 494702 152854
rect 494786 152618 495022 152854
rect 494466 134938 494702 135174
rect 494786 134938 495022 135174
rect 494466 134618 494702 134854
rect 494786 134618 495022 134854
rect 494466 116938 494702 117174
rect 494786 116938 495022 117174
rect 494466 116618 494702 116854
rect 494786 116618 495022 116854
rect 494466 98938 494702 99174
rect 494786 98938 495022 99174
rect 494466 98618 494702 98854
rect 494786 98618 495022 98854
rect 494466 80938 494702 81174
rect 494786 80938 495022 81174
rect 494466 80618 494702 80854
rect 494786 80618 495022 80854
rect 494466 62938 494702 63174
rect 494786 62938 495022 63174
rect 494466 62618 494702 62854
rect 494786 62618 495022 62854
rect 494466 44938 494702 45174
rect 494786 44938 495022 45174
rect 494466 44618 494702 44854
rect 494786 44618 495022 44854
rect 494466 26938 494702 27174
rect 494786 26938 495022 27174
rect 494466 26618 494702 26854
rect 494786 26618 495022 26854
rect 494466 8938 494702 9174
rect 494786 8938 495022 9174
rect 494466 8618 494702 8854
rect 494786 8618 495022 8854
rect 494466 -2052 494702 -1816
rect 494786 -2052 495022 -1816
rect 494466 -2372 494702 -2136
rect 494786 -2372 495022 -2136
rect 498186 462776 498422 463012
rect 498506 462776 498742 463012
rect 498186 462456 498422 462692
rect 498506 462456 498742 462692
rect 498186 444658 498422 444894
rect 498506 444658 498742 444894
rect 498186 444338 498422 444574
rect 498506 444338 498742 444574
rect 498186 426658 498422 426894
rect 498506 426658 498742 426894
rect 498186 426338 498422 426574
rect 498506 426338 498742 426574
rect 498186 408658 498422 408894
rect 498506 408658 498742 408894
rect 498186 408338 498422 408574
rect 498506 408338 498742 408574
rect 498186 390658 498422 390894
rect 498506 390658 498742 390894
rect 498186 390338 498422 390574
rect 498506 390338 498742 390574
rect 498186 372658 498422 372894
rect 498506 372658 498742 372894
rect 498186 372338 498422 372574
rect 498506 372338 498742 372574
rect 498186 354658 498422 354894
rect 498506 354658 498742 354894
rect 498186 354338 498422 354574
rect 498506 354338 498742 354574
rect 498186 336658 498422 336894
rect 498506 336658 498742 336894
rect 498186 336338 498422 336574
rect 498506 336338 498742 336574
rect 498186 318658 498422 318894
rect 498506 318658 498742 318894
rect 498186 318338 498422 318574
rect 498506 318338 498742 318574
rect 498186 300658 498422 300894
rect 498506 300658 498742 300894
rect 498186 300338 498422 300574
rect 498506 300338 498742 300574
rect 498186 282658 498422 282894
rect 498506 282658 498742 282894
rect 498186 282338 498422 282574
rect 498506 282338 498742 282574
rect 498186 264658 498422 264894
rect 498506 264658 498742 264894
rect 498186 264338 498422 264574
rect 498506 264338 498742 264574
rect 498186 246658 498422 246894
rect 498506 246658 498742 246894
rect 498186 246338 498422 246574
rect 498506 246338 498742 246574
rect 498186 228658 498422 228894
rect 498506 228658 498742 228894
rect 498186 228338 498422 228574
rect 498506 228338 498742 228574
rect 498186 210658 498422 210894
rect 498506 210658 498742 210894
rect 498186 210338 498422 210574
rect 498506 210338 498742 210574
rect 498186 192658 498422 192894
rect 498506 192658 498742 192894
rect 498186 192338 498422 192574
rect 498506 192338 498742 192574
rect 498186 174658 498422 174894
rect 498506 174658 498742 174894
rect 498186 174338 498422 174574
rect 498506 174338 498742 174574
rect 498186 156658 498422 156894
rect 498506 156658 498742 156894
rect 498186 156338 498422 156574
rect 498506 156338 498742 156574
rect 498186 138658 498422 138894
rect 498506 138658 498742 138894
rect 498186 138338 498422 138574
rect 498506 138338 498742 138574
rect 498186 120658 498422 120894
rect 498506 120658 498742 120894
rect 498186 120338 498422 120574
rect 498506 120338 498742 120574
rect 498186 102658 498422 102894
rect 498506 102658 498742 102894
rect 498186 102338 498422 102574
rect 498506 102338 498742 102574
rect 498186 84658 498422 84894
rect 498506 84658 498742 84894
rect 498186 84338 498422 84574
rect 498506 84338 498742 84574
rect 498186 66658 498422 66894
rect 498506 66658 498742 66894
rect 498186 66338 498422 66574
rect 498506 66338 498742 66574
rect 498186 48658 498422 48894
rect 498506 48658 498742 48894
rect 498186 48338 498422 48574
rect 498506 48338 498742 48574
rect 498186 30658 498422 30894
rect 498506 30658 498742 30894
rect 498186 30338 498422 30574
rect 498506 30338 498742 30574
rect 498186 12658 498422 12894
rect 498506 12658 498742 12894
rect 498186 12338 498422 12574
rect 498506 12338 498742 12574
rect 501906 463736 502142 463972
rect 502226 463736 502462 463972
rect 501906 463416 502142 463652
rect 502226 463416 502462 463652
rect 501906 448378 502142 448614
rect 502226 448378 502462 448614
rect 501906 448058 502142 448294
rect 502226 448058 502462 448294
rect 501906 430378 502142 430614
rect 502226 430378 502462 430614
rect 501906 430058 502142 430294
rect 502226 430058 502462 430294
rect 501906 412378 502142 412614
rect 502226 412378 502462 412614
rect 501906 412058 502142 412294
rect 502226 412058 502462 412294
rect 501906 394378 502142 394614
rect 502226 394378 502462 394614
rect 501906 394058 502142 394294
rect 502226 394058 502462 394294
rect 501906 376378 502142 376614
rect 502226 376378 502462 376614
rect 501906 376058 502142 376294
rect 502226 376058 502462 376294
rect 501906 358378 502142 358614
rect 502226 358378 502462 358614
rect 501906 358058 502142 358294
rect 502226 358058 502462 358294
rect 501906 340378 502142 340614
rect 502226 340378 502462 340614
rect 501906 340058 502142 340294
rect 502226 340058 502462 340294
rect 501906 322378 502142 322614
rect 502226 322378 502462 322614
rect 501906 322058 502142 322294
rect 502226 322058 502462 322294
rect 501906 304378 502142 304614
rect 502226 304378 502462 304614
rect 501906 304058 502142 304294
rect 502226 304058 502462 304294
rect 501906 286378 502142 286614
rect 502226 286378 502462 286614
rect 501906 286058 502142 286294
rect 502226 286058 502462 286294
rect 501906 268378 502142 268614
rect 502226 268378 502462 268614
rect 501906 268058 502142 268294
rect 502226 268058 502462 268294
rect 501906 250378 502142 250614
rect 502226 250378 502462 250614
rect 501906 250058 502142 250294
rect 502226 250058 502462 250294
rect 501906 232378 502142 232614
rect 502226 232378 502462 232614
rect 501906 232058 502142 232294
rect 502226 232058 502462 232294
rect 501906 214378 502142 214614
rect 502226 214378 502462 214614
rect 501906 214058 502142 214294
rect 502226 214058 502462 214294
rect 501906 196378 502142 196614
rect 502226 196378 502462 196614
rect 501906 196058 502142 196294
rect 502226 196058 502462 196294
rect 501906 178378 502142 178614
rect 502226 178378 502462 178614
rect 501906 178058 502142 178294
rect 502226 178058 502462 178294
rect 501906 160378 502142 160614
rect 502226 160378 502462 160614
rect 501906 160058 502142 160294
rect 502226 160058 502462 160294
rect 501906 142378 502142 142614
rect 502226 142378 502462 142614
rect 501906 142058 502142 142294
rect 502226 142058 502462 142294
rect 501906 124378 502142 124614
rect 502226 124378 502462 124614
rect 501906 124058 502142 124294
rect 502226 124058 502462 124294
rect 501906 106378 502142 106614
rect 502226 106378 502462 106614
rect 501906 106058 502142 106294
rect 502226 106058 502462 106294
rect 501906 88378 502142 88614
rect 502226 88378 502462 88614
rect 501906 88058 502142 88294
rect 502226 88058 502462 88294
rect 501906 70378 502142 70614
rect 502226 70378 502462 70614
rect 501906 70058 502142 70294
rect 502226 70058 502462 70294
rect 501906 52378 502142 52614
rect 502226 52378 502462 52614
rect 501906 52058 502142 52294
rect 502226 52058 502462 52294
rect 501906 34378 502142 34614
rect 502226 34378 502462 34614
rect 501906 34058 502142 34294
rect 502226 34058 502462 34294
rect 501906 16378 502142 16614
rect 502226 16378 502462 16614
rect 501906 16058 502142 16294
rect 502226 16058 502462 16294
rect 508746 460856 508982 461092
rect 509066 460856 509302 461092
rect 508746 460536 508982 460772
rect 509066 460536 509302 460772
rect 508746 455218 508982 455454
rect 509066 455218 509302 455454
rect 508746 454898 508982 455134
rect 509066 454898 509302 455134
rect 508746 437218 508982 437454
rect 509066 437218 509302 437454
rect 508746 436898 508982 437134
rect 509066 436898 509302 437134
rect 508746 419218 508982 419454
rect 509066 419218 509302 419454
rect 508746 418898 508982 419134
rect 509066 418898 509302 419134
rect 508746 401218 508982 401454
rect 509066 401218 509302 401454
rect 508746 400898 508982 401134
rect 509066 400898 509302 401134
rect 508746 383218 508982 383454
rect 509066 383218 509302 383454
rect 508746 382898 508982 383134
rect 509066 382898 509302 383134
rect 508746 365218 508982 365454
rect 509066 365218 509302 365454
rect 508746 364898 508982 365134
rect 509066 364898 509302 365134
rect 508746 347218 508982 347454
rect 509066 347218 509302 347454
rect 508746 346898 508982 347134
rect 509066 346898 509302 347134
rect 508746 329218 508982 329454
rect 509066 329218 509302 329454
rect 508746 328898 508982 329134
rect 509066 328898 509302 329134
rect 508746 311218 508982 311454
rect 509066 311218 509302 311454
rect 508746 310898 508982 311134
rect 509066 310898 509302 311134
rect 508746 293218 508982 293454
rect 509066 293218 509302 293454
rect 508746 292898 508982 293134
rect 509066 292898 509302 293134
rect 508746 275218 508982 275454
rect 509066 275218 509302 275454
rect 508746 274898 508982 275134
rect 509066 274898 509302 275134
rect 508746 257218 508982 257454
rect 509066 257218 509302 257454
rect 508746 256898 508982 257134
rect 509066 256898 509302 257134
rect 508746 239218 508982 239454
rect 509066 239218 509302 239454
rect 508746 238898 508982 239134
rect 509066 238898 509302 239134
rect 508746 221218 508982 221454
rect 509066 221218 509302 221454
rect 508746 220898 508982 221134
rect 509066 220898 509302 221134
rect 508746 203218 508982 203454
rect 509066 203218 509302 203454
rect 508746 202898 508982 203134
rect 509066 202898 509302 203134
rect 508746 185218 508982 185454
rect 509066 185218 509302 185454
rect 508746 184898 508982 185134
rect 509066 184898 509302 185134
rect 508746 167218 508982 167454
rect 509066 167218 509302 167454
rect 508746 166898 508982 167134
rect 509066 166898 509302 167134
rect 508746 149218 508982 149454
rect 509066 149218 509302 149454
rect 508746 148898 508982 149134
rect 509066 148898 509302 149134
rect 508746 131218 508982 131454
rect 509066 131218 509302 131454
rect 508746 130898 508982 131134
rect 509066 130898 509302 131134
rect 508746 113218 508982 113454
rect 509066 113218 509302 113454
rect 508746 112898 508982 113134
rect 509066 112898 509302 113134
rect 508746 95218 508982 95454
rect 509066 95218 509302 95454
rect 508746 94898 508982 95134
rect 509066 94898 509302 95134
rect 508746 77218 508982 77454
rect 509066 77218 509302 77454
rect 508746 76898 508982 77134
rect 509066 76898 509302 77134
rect 508746 59218 508982 59454
rect 509066 59218 509302 59454
rect 508746 58898 508982 59134
rect 509066 58898 509302 59134
rect 508746 41218 508982 41454
rect 509066 41218 509302 41454
rect 508746 40898 508982 41134
rect 509066 40898 509302 41134
rect 508746 23218 508982 23454
rect 509066 23218 509302 23454
rect 508746 22898 508982 23134
rect 509066 22898 509302 23134
rect 508746 5218 508982 5454
rect 509066 5218 509302 5454
rect 508746 4898 508982 5134
rect 509066 4898 509302 5134
rect 512466 461816 512702 462052
rect 512786 461816 513022 462052
rect 512466 461496 512702 461732
rect 512786 461496 513022 461732
rect 512466 440938 512702 441174
rect 512786 440938 513022 441174
rect 512466 440618 512702 440854
rect 512786 440618 513022 440854
rect 512466 422938 512702 423174
rect 512786 422938 513022 423174
rect 512466 422618 512702 422854
rect 512786 422618 513022 422854
rect 512466 404938 512702 405174
rect 512786 404938 513022 405174
rect 512466 404618 512702 404854
rect 512786 404618 513022 404854
rect 512466 386938 512702 387174
rect 512786 386938 513022 387174
rect 512466 386618 512702 386854
rect 512786 386618 513022 386854
rect 512466 368938 512702 369174
rect 512786 368938 513022 369174
rect 512466 368618 512702 368854
rect 512786 368618 513022 368854
rect 512466 350938 512702 351174
rect 512786 350938 513022 351174
rect 512466 350618 512702 350854
rect 512786 350618 513022 350854
rect 512466 332938 512702 333174
rect 512786 332938 513022 333174
rect 512466 332618 512702 332854
rect 512786 332618 513022 332854
rect 512466 314938 512702 315174
rect 512786 314938 513022 315174
rect 512466 314618 512702 314854
rect 512786 314618 513022 314854
rect 512466 296938 512702 297174
rect 512786 296938 513022 297174
rect 512466 296618 512702 296854
rect 512786 296618 513022 296854
rect 512466 278938 512702 279174
rect 512786 278938 513022 279174
rect 512466 278618 512702 278854
rect 512786 278618 513022 278854
rect 512466 260938 512702 261174
rect 512786 260938 513022 261174
rect 512466 260618 512702 260854
rect 512786 260618 513022 260854
rect 512466 242938 512702 243174
rect 512786 242938 513022 243174
rect 512466 242618 512702 242854
rect 512786 242618 513022 242854
rect 512466 224938 512702 225174
rect 512786 224938 513022 225174
rect 512466 224618 512702 224854
rect 512786 224618 513022 224854
rect 512466 206938 512702 207174
rect 512786 206938 513022 207174
rect 512466 206618 512702 206854
rect 512786 206618 513022 206854
rect 512466 188938 512702 189174
rect 512786 188938 513022 189174
rect 512466 188618 512702 188854
rect 512786 188618 513022 188854
rect 512466 170938 512702 171174
rect 512786 170938 513022 171174
rect 512466 170618 512702 170854
rect 512786 170618 513022 170854
rect 512466 152938 512702 153174
rect 512786 152938 513022 153174
rect 512466 152618 512702 152854
rect 512786 152618 513022 152854
rect 512466 134938 512702 135174
rect 512786 134938 513022 135174
rect 512466 134618 512702 134854
rect 512786 134618 513022 134854
rect 512466 116938 512702 117174
rect 512786 116938 513022 117174
rect 512466 116618 512702 116854
rect 512786 116618 513022 116854
rect 512466 98938 512702 99174
rect 512786 98938 513022 99174
rect 512466 98618 512702 98854
rect 512786 98618 513022 98854
rect 512466 80938 512702 81174
rect 512786 80938 513022 81174
rect 512466 80618 512702 80854
rect 512786 80618 513022 80854
rect 512466 62938 512702 63174
rect 512786 62938 513022 63174
rect 512466 62618 512702 62854
rect 512786 62618 513022 62854
rect 512466 44938 512702 45174
rect 512786 44938 513022 45174
rect 512466 44618 512702 44854
rect 512786 44618 513022 44854
rect 512466 26938 512702 27174
rect 512786 26938 513022 27174
rect 512466 26618 512702 26854
rect 512786 26618 513022 26854
rect 512466 8938 512702 9174
rect 512786 8938 513022 9174
rect 512466 8618 512702 8854
rect 512786 8618 513022 8854
rect 516186 462776 516422 463012
rect 516506 462776 516742 463012
rect 516186 462456 516422 462692
rect 516506 462456 516742 462692
rect 516186 444658 516422 444894
rect 516506 444658 516742 444894
rect 516186 444338 516422 444574
rect 516506 444338 516742 444574
rect 516186 426658 516422 426894
rect 516506 426658 516742 426894
rect 516186 426338 516422 426574
rect 516506 426338 516742 426574
rect 516186 408658 516422 408894
rect 516506 408658 516742 408894
rect 516186 408338 516422 408574
rect 516506 408338 516742 408574
rect 516186 390658 516422 390894
rect 516506 390658 516742 390894
rect 516186 390338 516422 390574
rect 516506 390338 516742 390574
rect 516186 372658 516422 372894
rect 516506 372658 516742 372894
rect 516186 372338 516422 372574
rect 516506 372338 516742 372574
rect 516186 354658 516422 354894
rect 516506 354658 516742 354894
rect 516186 354338 516422 354574
rect 516506 354338 516742 354574
rect 516186 336658 516422 336894
rect 516506 336658 516742 336894
rect 516186 336338 516422 336574
rect 516506 336338 516742 336574
rect 516186 318658 516422 318894
rect 516506 318658 516742 318894
rect 516186 318338 516422 318574
rect 516506 318338 516742 318574
rect 516186 300658 516422 300894
rect 516506 300658 516742 300894
rect 516186 300338 516422 300574
rect 516506 300338 516742 300574
rect 516186 282658 516422 282894
rect 516506 282658 516742 282894
rect 516186 282338 516422 282574
rect 516506 282338 516742 282574
rect 516186 264658 516422 264894
rect 516506 264658 516742 264894
rect 516186 264338 516422 264574
rect 516506 264338 516742 264574
rect 516186 246658 516422 246894
rect 516506 246658 516742 246894
rect 516186 246338 516422 246574
rect 516506 246338 516742 246574
rect 516186 228658 516422 228894
rect 516506 228658 516742 228894
rect 516186 228338 516422 228574
rect 516506 228338 516742 228574
rect 516186 210658 516422 210894
rect 516506 210658 516742 210894
rect 516186 210338 516422 210574
rect 516506 210338 516742 210574
rect 516186 192658 516422 192894
rect 516506 192658 516742 192894
rect 516186 192338 516422 192574
rect 516506 192338 516742 192574
rect 516186 174658 516422 174894
rect 516506 174658 516742 174894
rect 516186 174338 516422 174574
rect 516506 174338 516742 174574
rect 516186 156658 516422 156894
rect 516506 156658 516742 156894
rect 516186 156338 516422 156574
rect 516506 156338 516742 156574
rect 516186 138658 516422 138894
rect 516506 138658 516742 138894
rect 516186 138338 516422 138574
rect 516506 138338 516742 138574
rect 516186 120658 516422 120894
rect 516506 120658 516742 120894
rect 516186 120338 516422 120574
rect 516506 120338 516742 120574
rect 516186 102658 516422 102894
rect 516506 102658 516742 102894
rect 516186 102338 516422 102574
rect 516506 102338 516742 102574
rect 516186 84658 516422 84894
rect 516506 84658 516742 84894
rect 516186 84338 516422 84574
rect 516506 84338 516742 84574
rect 516186 66658 516422 66894
rect 516506 66658 516742 66894
rect 516186 66338 516422 66574
rect 516506 66338 516742 66574
rect 516186 48658 516422 48894
rect 516506 48658 516742 48894
rect 516186 48338 516422 48574
rect 516506 48338 516742 48574
rect 516186 30658 516422 30894
rect 516506 30658 516742 30894
rect 516186 30338 516422 30574
rect 516506 30338 516742 30574
rect 516186 12658 516422 12894
rect 516506 12658 516742 12894
rect 516186 12338 516422 12574
rect 516506 12338 516742 12574
rect 519906 463736 520142 463972
rect 520226 463736 520462 463972
rect 519906 463416 520142 463652
rect 520226 463416 520462 463652
rect 519906 448378 520142 448614
rect 520226 448378 520462 448614
rect 519906 448058 520142 448294
rect 520226 448058 520462 448294
rect 519906 430378 520142 430614
rect 520226 430378 520462 430614
rect 519906 430058 520142 430294
rect 520226 430058 520462 430294
rect 519906 412378 520142 412614
rect 520226 412378 520462 412614
rect 519906 412058 520142 412294
rect 520226 412058 520462 412294
rect 519906 394378 520142 394614
rect 520226 394378 520462 394614
rect 519906 394058 520142 394294
rect 520226 394058 520462 394294
rect 519906 376378 520142 376614
rect 520226 376378 520462 376614
rect 519906 376058 520142 376294
rect 520226 376058 520462 376294
rect 519906 358378 520142 358614
rect 520226 358378 520462 358614
rect 519906 358058 520142 358294
rect 520226 358058 520462 358294
rect 519906 340378 520142 340614
rect 520226 340378 520462 340614
rect 519906 340058 520142 340294
rect 520226 340058 520462 340294
rect 519906 322378 520142 322614
rect 520226 322378 520462 322614
rect 519906 322058 520142 322294
rect 520226 322058 520462 322294
rect 519906 304378 520142 304614
rect 520226 304378 520462 304614
rect 519906 304058 520142 304294
rect 520226 304058 520462 304294
rect 519906 286378 520142 286614
rect 520226 286378 520462 286614
rect 519906 286058 520142 286294
rect 520226 286058 520462 286294
rect 519906 268378 520142 268614
rect 520226 268378 520462 268614
rect 519906 268058 520142 268294
rect 520226 268058 520462 268294
rect 519906 250378 520142 250614
rect 520226 250378 520462 250614
rect 519906 250058 520142 250294
rect 520226 250058 520462 250294
rect 519906 232378 520142 232614
rect 520226 232378 520462 232614
rect 519906 232058 520142 232294
rect 520226 232058 520462 232294
rect 519906 214378 520142 214614
rect 520226 214378 520462 214614
rect 519906 214058 520142 214294
rect 520226 214058 520462 214294
rect 519906 196378 520142 196614
rect 520226 196378 520462 196614
rect 519906 196058 520142 196294
rect 520226 196058 520462 196294
rect 519906 178378 520142 178614
rect 520226 178378 520462 178614
rect 519906 178058 520142 178294
rect 520226 178058 520462 178294
rect 519906 160378 520142 160614
rect 520226 160378 520462 160614
rect 519906 160058 520142 160294
rect 520226 160058 520462 160294
rect 519906 142378 520142 142614
rect 520226 142378 520462 142614
rect 519906 142058 520142 142294
rect 520226 142058 520462 142294
rect 519906 124378 520142 124614
rect 520226 124378 520462 124614
rect 519906 124058 520142 124294
rect 520226 124058 520462 124294
rect 519906 106378 520142 106614
rect 520226 106378 520462 106614
rect 519906 106058 520142 106294
rect 520226 106058 520462 106294
rect 519906 88378 520142 88614
rect 520226 88378 520462 88614
rect 519906 88058 520142 88294
rect 520226 88058 520462 88294
rect 519906 70378 520142 70614
rect 520226 70378 520462 70614
rect 519906 70058 520142 70294
rect 520226 70058 520462 70294
rect 519906 52378 520142 52614
rect 520226 52378 520462 52614
rect 519906 52058 520142 52294
rect 520226 52058 520462 52294
rect 519906 34378 520142 34614
rect 520226 34378 520462 34614
rect 519906 34058 520142 34294
rect 520226 34058 520462 34294
rect 519906 16378 520142 16614
rect 520226 16378 520462 16614
rect 519906 16058 520142 16294
rect 520226 16058 520462 16294
rect 526746 460856 526982 461092
rect 527066 460856 527302 461092
rect 526746 460536 526982 460772
rect 527066 460536 527302 460772
rect 526746 455218 526982 455454
rect 527066 455218 527302 455454
rect 526746 454898 526982 455134
rect 527066 454898 527302 455134
rect 526746 437218 526982 437454
rect 527066 437218 527302 437454
rect 526746 436898 526982 437134
rect 527066 436898 527302 437134
rect 526746 419218 526982 419454
rect 527066 419218 527302 419454
rect 526746 418898 526982 419134
rect 527066 418898 527302 419134
rect 526746 401218 526982 401454
rect 527066 401218 527302 401454
rect 526746 400898 526982 401134
rect 527066 400898 527302 401134
rect 526746 383218 526982 383454
rect 527066 383218 527302 383454
rect 526746 382898 526982 383134
rect 527066 382898 527302 383134
rect 526746 365218 526982 365454
rect 527066 365218 527302 365454
rect 526746 364898 526982 365134
rect 527066 364898 527302 365134
rect 526746 347218 526982 347454
rect 527066 347218 527302 347454
rect 526746 346898 526982 347134
rect 527066 346898 527302 347134
rect 526746 329218 526982 329454
rect 527066 329218 527302 329454
rect 526746 328898 526982 329134
rect 527066 328898 527302 329134
rect 526746 311218 526982 311454
rect 527066 311218 527302 311454
rect 526746 310898 526982 311134
rect 527066 310898 527302 311134
rect 526746 293218 526982 293454
rect 527066 293218 527302 293454
rect 526746 292898 526982 293134
rect 527066 292898 527302 293134
rect 526746 275218 526982 275454
rect 527066 275218 527302 275454
rect 526746 274898 526982 275134
rect 527066 274898 527302 275134
rect 526746 257218 526982 257454
rect 527066 257218 527302 257454
rect 526746 256898 526982 257134
rect 527066 256898 527302 257134
rect 526746 239218 526982 239454
rect 527066 239218 527302 239454
rect 526746 238898 526982 239134
rect 527066 238898 527302 239134
rect 526746 221218 526982 221454
rect 527066 221218 527302 221454
rect 526746 220898 526982 221134
rect 527066 220898 527302 221134
rect 526746 203218 526982 203454
rect 527066 203218 527302 203454
rect 526746 202898 526982 203134
rect 527066 202898 527302 203134
rect 526746 185218 526982 185454
rect 527066 185218 527302 185454
rect 526746 184898 526982 185134
rect 527066 184898 527302 185134
rect 526746 167218 526982 167454
rect 527066 167218 527302 167454
rect 526746 166898 526982 167134
rect 527066 166898 527302 167134
rect 526746 149218 526982 149454
rect 527066 149218 527302 149454
rect 526746 148898 526982 149134
rect 527066 148898 527302 149134
rect 526746 131218 526982 131454
rect 527066 131218 527302 131454
rect 526746 130898 526982 131134
rect 527066 130898 527302 131134
rect 526746 113218 526982 113454
rect 527066 113218 527302 113454
rect 526746 112898 526982 113134
rect 527066 112898 527302 113134
rect 526746 95218 526982 95454
rect 527066 95218 527302 95454
rect 526746 94898 526982 95134
rect 527066 94898 527302 95134
rect 526746 77218 526982 77454
rect 527066 77218 527302 77454
rect 526746 76898 526982 77134
rect 527066 76898 527302 77134
rect 526746 59218 526982 59454
rect 527066 59218 527302 59454
rect 526746 58898 526982 59134
rect 527066 58898 527302 59134
rect 526746 41218 526982 41454
rect 527066 41218 527302 41454
rect 526746 40898 526982 41134
rect 527066 40898 527302 41134
rect 526746 23218 526982 23454
rect 527066 23218 527302 23454
rect 526746 22898 526982 23134
rect 527066 22898 527302 23134
rect 526746 5218 526982 5454
rect 527066 5218 527302 5454
rect 526746 4898 526982 5134
rect 527066 4898 527302 5134
rect 530466 461816 530702 462052
rect 530786 461816 531022 462052
rect 530466 461496 530702 461732
rect 530786 461496 531022 461732
rect 530466 440938 530702 441174
rect 530786 440938 531022 441174
rect 530466 440618 530702 440854
rect 530786 440618 531022 440854
rect 530466 422938 530702 423174
rect 530786 422938 531022 423174
rect 530466 422618 530702 422854
rect 530786 422618 531022 422854
rect 530466 404938 530702 405174
rect 530786 404938 531022 405174
rect 530466 404618 530702 404854
rect 530786 404618 531022 404854
rect 530466 386938 530702 387174
rect 530786 386938 531022 387174
rect 530466 386618 530702 386854
rect 530786 386618 531022 386854
rect 530466 368938 530702 369174
rect 530786 368938 531022 369174
rect 530466 368618 530702 368854
rect 530786 368618 531022 368854
rect 530466 350938 530702 351174
rect 530786 350938 531022 351174
rect 530466 350618 530702 350854
rect 530786 350618 531022 350854
rect 530466 332938 530702 333174
rect 530786 332938 531022 333174
rect 530466 332618 530702 332854
rect 530786 332618 531022 332854
rect 530466 314938 530702 315174
rect 530786 314938 531022 315174
rect 530466 314618 530702 314854
rect 530786 314618 531022 314854
rect 530466 296938 530702 297174
rect 530786 296938 531022 297174
rect 530466 296618 530702 296854
rect 530786 296618 531022 296854
rect 530466 278938 530702 279174
rect 530786 278938 531022 279174
rect 530466 278618 530702 278854
rect 530786 278618 531022 278854
rect 530466 260938 530702 261174
rect 530786 260938 531022 261174
rect 530466 260618 530702 260854
rect 530786 260618 531022 260854
rect 530466 242938 530702 243174
rect 530786 242938 531022 243174
rect 530466 242618 530702 242854
rect 530786 242618 531022 242854
rect 530466 224938 530702 225174
rect 530786 224938 531022 225174
rect 530466 224618 530702 224854
rect 530786 224618 531022 224854
rect 530466 206938 530702 207174
rect 530786 206938 531022 207174
rect 530466 206618 530702 206854
rect 530786 206618 531022 206854
rect 530466 188938 530702 189174
rect 530786 188938 531022 189174
rect 530466 188618 530702 188854
rect 530786 188618 531022 188854
rect 530466 170938 530702 171174
rect 530786 170938 531022 171174
rect 530466 170618 530702 170854
rect 530786 170618 531022 170854
rect 530466 152938 530702 153174
rect 530786 152938 531022 153174
rect 530466 152618 530702 152854
rect 530786 152618 531022 152854
rect 530466 134938 530702 135174
rect 530786 134938 531022 135174
rect 530466 134618 530702 134854
rect 530786 134618 531022 134854
rect 530466 116938 530702 117174
rect 530786 116938 531022 117174
rect 530466 116618 530702 116854
rect 530786 116618 531022 116854
rect 530466 98938 530702 99174
rect 530786 98938 531022 99174
rect 530466 98618 530702 98854
rect 530786 98618 531022 98854
rect 530466 80938 530702 81174
rect 530786 80938 531022 81174
rect 530466 80618 530702 80854
rect 530786 80618 531022 80854
rect 530466 62938 530702 63174
rect 530786 62938 531022 63174
rect 530466 62618 530702 62854
rect 530786 62618 531022 62854
rect 530466 44938 530702 45174
rect 530786 44938 531022 45174
rect 530466 44618 530702 44854
rect 530786 44618 531022 44854
rect 530466 26938 530702 27174
rect 530786 26938 531022 27174
rect 530466 26618 530702 26854
rect 530786 26618 531022 26854
rect 530466 8938 530702 9174
rect 530786 8938 531022 9174
rect 530466 8618 530702 8854
rect 530786 8618 531022 8854
rect 534186 462776 534422 463012
rect 534506 462776 534742 463012
rect 534186 462456 534422 462692
rect 534506 462456 534742 462692
rect 534186 444658 534422 444894
rect 534506 444658 534742 444894
rect 534186 444338 534422 444574
rect 534506 444338 534742 444574
rect 534186 426658 534422 426894
rect 534506 426658 534742 426894
rect 534186 426338 534422 426574
rect 534506 426338 534742 426574
rect 534186 408658 534422 408894
rect 534506 408658 534742 408894
rect 534186 408338 534422 408574
rect 534506 408338 534742 408574
rect 534186 390658 534422 390894
rect 534506 390658 534742 390894
rect 534186 390338 534422 390574
rect 534506 390338 534742 390574
rect 534186 372658 534422 372894
rect 534506 372658 534742 372894
rect 534186 372338 534422 372574
rect 534506 372338 534742 372574
rect 534186 354658 534422 354894
rect 534506 354658 534742 354894
rect 534186 354338 534422 354574
rect 534506 354338 534742 354574
rect 534186 336658 534422 336894
rect 534506 336658 534742 336894
rect 534186 336338 534422 336574
rect 534506 336338 534742 336574
rect 534186 318658 534422 318894
rect 534506 318658 534742 318894
rect 534186 318338 534422 318574
rect 534506 318338 534742 318574
rect 534186 300658 534422 300894
rect 534506 300658 534742 300894
rect 534186 300338 534422 300574
rect 534506 300338 534742 300574
rect 534186 282658 534422 282894
rect 534506 282658 534742 282894
rect 534186 282338 534422 282574
rect 534506 282338 534742 282574
rect 534186 264658 534422 264894
rect 534506 264658 534742 264894
rect 534186 264338 534422 264574
rect 534506 264338 534742 264574
rect 534186 246658 534422 246894
rect 534506 246658 534742 246894
rect 534186 246338 534422 246574
rect 534506 246338 534742 246574
rect 534186 228658 534422 228894
rect 534506 228658 534742 228894
rect 534186 228338 534422 228574
rect 534506 228338 534742 228574
rect 534186 210658 534422 210894
rect 534506 210658 534742 210894
rect 534186 210338 534422 210574
rect 534506 210338 534742 210574
rect 534186 192658 534422 192894
rect 534506 192658 534742 192894
rect 534186 192338 534422 192574
rect 534506 192338 534742 192574
rect 534186 174658 534422 174894
rect 534506 174658 534742 174894
rect 534186 174338 534422 174574
rect 534506 174338 534742 174574
rect 534186 156658 534422 156894
rect 534506 156658 534742 156894
rect 534186 156338 534422 156574
rect 534506 156338 534742 156574
rect 534186 138658 534422 138894
rect 534506 138658 534742 138894
rect 534186 138338 534422 138574
rect 534506 138338 534742 138574
rect 534186 120658 534422 120894
rect 534506 120658 534742 120894
rect 534186 120338 534422 120574
rect 534506 120338 534742 120574
rect 534186 102658 534422 102894
rect 534506 102658 534742 102894
rect 534186 102338 534422 102574
rect 534506 102338 534742 102574
rect 534186 84658 534422 84894
rect 534506 84658 534742 84894
rect 534186 84338 534422 84574
rect 534506 84338 534742 84574
rect 534186 66658 534422 66894
rect 534506 66658 534742 66894
rect 534186 66338 534422 66574
rect 534506 66338 534742 66574
rect 534186 48658 534422 48894
rect 534506 48658 534742 48894
rect 534186 48338 534422 48574
rect 534506 48338 534742 48574
rect 534186 30658 534422 30894
rect 534506 30658 534742 30894
rect 534186 30338 534422 30574
rect 534506 30338 534742 30574
rect 534186 12658 534422 12894
rect 534506 12658 534742 12894
rect 534186 12338 534422 12574
rect 534506 12338 534742 12574
rect 537906 463736 538142 463972
rect 538226 463736 538462 463972
rect 537906 463416 538142 463652
rect 538226 463416 538462 463652
rect 547884 463736 548120 463972
rect 548204 463736 548440 463972
rect 547884 463416 548120 463652
rect 548204 463416 548440 463652
rect 546924 462776 547160 463012
rect 547244 462776 547480 463012
rect 546924 462456 547160 462692
rect 547244 462456 547480 462692
rect 545964 461816 546200 462052
rect 546284 461816 546520 462052
rect 545964 461496 546200 461732
rect 546284 461496 546520 461732
rect 537906 448378 538142 448614
rect 538226 448378 538462 448614
rect 537906 448058 538142 448294
rect 538226 448058 538462 448294
rect 537906 430378 538142 430614
rect 538226 430378 538462 430614
rect 537906 430058 538142 430294
rect 538226 430058 538462 430294
rect 537906 412378 538142 412614
rect 538226 412378 538462 412614
rect 537906 412058 538142 412294
rect 538226 412058 538462 412294
rect 537906 394378 538142 394614
rect 538226 394378 538462 394614
rect 537906 394058 538142 394294
rect 538226 394058 538462 394294
rect 537906 376378 538142 376614
rect 538226 376378 538462 376614
rect 537906 376058 538142 376294
rect 538226 376058 538462 376294
rect 537906 358378 538142 358614
rect 538226 358378 538462 358614
rect 537906 358058 538142 358294
rect 538226 358058 538462 358294
rect 537906 340378 538142 340614
rect 538226 340378 538462 340614
rect 537906 340058 538142 340294
rect 538226 340058 538462 340294
rect 537906 322378 538142 322614
rect 538226 322378 538462 322614
rect 537906 322058 538142 322294
rect 538226 322058 538462 322294
rect 537906 304378 538142 304614
rect 538226 304378 538462 304614
rect 537906 304058 538142 304294
rect 538226 304058 538462 304294
rect 537906 286378 538142 286614
rect 538226 286378 538462 286614
rect 537906 286058 538142 286294
rect 538226 286058 538462 286294
rect 537906 268378 538142 268614
rect 538226 268378 538462 268614
rect 537906 268058 538142 268294
rect 538226 268058 538462 268294
rect 537906 250378 538142 250614
rect 538226 250378 538462 250614
rect 537906 250058 538142 250294
rect 538226 250058 538462 250294
rect 537906 232378 538142 232614
rect 538226 232378 538462 232614
rect 537906 232058 538142 232294
rect 538226 232058 538462 232294
rect 537906 214378 538142 214614
rect 538226 214378 538462 214614
rect 537906 214058 538142 214294
rect 538226 214058 538462 214294
rect 537906 196378 538142 196614
rect 538226 196378 538462 196614
rect 537906 196058 538142 196294
rect 538226 196058 538462 196294
rect 537906 178378 538142 178614
rect 538226 178378 538462 178614
rect 537906 178058 538142 178294
rect 538226 178058 538462 178294
rect 537906 160378 538142 160614
rect 538226 160378 538462 160614
rect 537906 160058 538142 160294
rect 538226 160058 538462 160294
rect 537906 142378 538142 142614
rect 538226 142378 538462 142614
rect 537906 142058 538142 142294
rect 538226 142058 538462 142294
rect 537906 124378 538142 124614
rect 538226 124378 538462 124614
rect 537906 124058 538142 124294
rect 538226 124058 538462 124294
rect 537906 106378 538142 106614
rect 538226 106378 538462 106614
rect 537906 106058 538142 106294
rect 538226 106058 538462 106294
rect 537906 88378 538142 88614
rect 538226 88378 538462 88614
rect 537906 88058 538142 88294
rect 538226 88058 538462 88294
rect 537906 70378 538142 70614
rect 538226 70378 538462 70614
rect 537906 70058 538142 70294
rect 538226 70058 538462 70294
rect 537906 52378 538142 52614
rect 538226 52378 538462 52614
rect 537906 52058 538142 52294
rect 538226 52058 538462 52294
rect 537906 34378 538142 34614
rect 538226 34378 538462 34614
rect 537906 34058 538142 34294
rect 538226 34058 538462 34294
rect 537906 16378 538142 16614
rect 538226 16378 538462 16614
rect 537906 16058 538142 16294
rect 538226 16058 538462 16294
rect 545004 460856 545240 461092
rect 545324 460856 545560 461092
rect 545004 460536 545240 460772
rect 545324 460536 545560 460772
rect 545004 455218 545240 455454
rect 545324 455218 545560 455454
rect 545004 454898 545240 455134
rect 545324 454898 545560 455134
rect 545004 437218 545240 437454
rect 545324 437218 545560 437454
rect 545004 436898 545240 437134
rect 545324 436898 545560 437134
rect 545004 419218 545240 419454
rect 545324 419218 545560 419454
rect 545004 418898 545240 419134
rect 545324 418898 545560 419134
rect 545004 401218 545240 401454
rect 545324 401218 545560 401454
rect 545004 400898 545240 401134
rect 545324 400898 545560 401134
rect 545004 383218 545240 383454
rect 545324 383218 545560 383454
rect 545004 382898 545240 383134
rect 545324 382898 545560 383134
rect 545004 365218 545240 365454
rect 545324 365218 545560 365454
rect 545004 364898 545240 365134
rect 545324 364898 545560 365134
rect 545004 347218 545240 347454
rect 545324 347218 545560 347454
rect 545004 346898 545240 347134
rect 545324 346898 545560 347134
rect 545004 329218 545240 329454
rect 545324 329218 545560 329454
rect 545004 328898 545240 329134
rect 545324 328898 545560 329134
rect 545004 311218 545240 311454
rect 545324 311218 545560 311454
rect 545004 310898 545240 311134
rect 545324 310898 545560 311134
rect 545004 293218 545240 293454
rect 545324 293218 545560 293454
rect 545004 292898 545240 293134
rect 545324 292898 545560 293134
rect 545004 275218 545240 275454
rect 545324 275218 545560 275454
rect 545004 274898 545240 275134
rect 545324 274898 545560 275134
rect 545004 257218 545240 257454
rect 545324 257218 545560 257454
rect 545004 256898 545240 257134
rect 545324 256898 545560 257134
rect 545004 239218 545240 239454
rect 545324 239218 545560 239454
rect 545004 238898 545240 239134
rect 545324 238898 545560 239134
rect 545004 221218 545240 221454
rect 545324 221218 545560 221454
rect 545004 220898 545240 221134
rect 545324 220898 545560 221134
rect 545004 203218 545240 203454
rect 545324 203218 545560 203454
rect 545004 202898 545240 203134
rect 545324 202898 545560 203134
rect 545004 185218 545240 185454
rect 545324 185218 545560 185454
rect 545004 184898 545240 185134
rect 545324 184898 545560 185134
rect 545004 167218 545240 167454
rect 545324 167218 545560 167454
rect 545004 166898 545240 167134
rect 545324 166898 545560 167134
rect 545004 149218 545240 149454
rect 545324 149218 545560 149454
rect 545004 148898 545240 149134
rect 545324 148898 545560 149134
rect 545004 131218 545240 131454
rect 545324 131218 545560 131454
rect 545004 130898 545240 131134
rect 545324 130898 545560 131134
rect 545004 113218 545240 113454
rect 545324 113218 545560 113454
rect 545004 112898 545240 113134
rect 545324 112898 545560 113134
rect 545004 95218 545240 95454
rect 545324 95218 545560 95454
rect 545004 94898 545240 95134
rect 545324 94898 545560 95134
rect 545004 77218 545240 77454
rect 545324 77218 545560 77454
rect 545004 76898 545240 77134
rect 545324 76898 545560 77134
rect 545004 59218 545240 59454
rect 545324 59218 545560 59454
rect 545004 58898 545240 59134
rect 545324 58898 545560 59134
rect 545004 41218 545240 41454
rect 545324 41218 545560 41454
rect 545004 40898 545240 41134
rect 545324 40898 545560 41134
rect 545004 23218 545240 23454
rect 545324 23218 545560 23454
rect 545004 22898 545240 23134
rect 545324 22898 545560 23134
rect 545004 5218 545240 5454
rect 545324 5218 545560 5454
rect 545004 4898 545240 5134
rect 545324 4898 545560 5134
rect 545004 -1092 545240 -856
rect 545324 -1092 545560 -856
rect 545004 -1412 545240 -1176
rect 545324 -1412 545560 -1176
rect 545964 440938 546200 441174
rect 546284 440938 546520 441174
rect 545964 440618 546200 440854
rect 546284 440618 546520 440854
rect 545964 422938 546200 423174
rect 546284 422938 546520 423174
rect 545964 422618 546200 422854
rect 546284 422618 546520 422854
rect 545964 404938 546200 405174
rect 546284 404938 546520 405174
rect 545964 404618 546200 404854
rect 546284 404618 546520 404854
rect 545964 386938 546200 387174
rect 546284 386938 546520 387174
rect 545964 386618 546200 386854
rect 546284 386618 546520 386854
rect 545964 368938 546200 369174
rect 546284 368938 546520 369174
rect 545964 368618 546200 368854
rect 546284 368618 546520 368854
rect 545964 350938 546200 351174
rect 546284 350938 546520 351174
rect 545964 350618 546200 350854
rect 546284 350618 546520 350854
rect 545964 332938 546200 333174
rect 546284 332938 546520 333174
rect 545964 332618 546200 332854
rect 546284 332618 546520 332854
rect 545964 314938 546200 315174
rect 546284 314938 546520 315174
rect 545964 314618 546200 314854
rect 546284 314618 546520 314854
rect 545964 296938 546200 297174
rect 546284 296938 546520 297174
rect 545964 296618 546200 296854
rect 546284 296618 546520 296854
rect 545964 278938 546200 279174
rect 546284 278938 546520 279174
rect 545964 278618 546200 278854
rect 546284 278618 546520 278854
rect 545964 260938 546200 261174
rect 546284 260938 546520 261174
rect 545964 260618 546200 260854
rect 546284 260618 546520 260854
rect 545964 242938 546200 243174
rect 546284 242938 546520 243174
rect 545964 242618 546200 242854
rect 546284 242618 546520 242854
rect 545964 224938 546200 225174
rect 546284 224938 546520 225174
rect 545964 224618 546200 224854
rect 546284 224618 546520 224854
rect 545964 206938 546200 207174
rect 546284 206938 546520 207174
rect 545964 206618 546200 206854
rect 546284 206618 546520 206854
rect 545964 188938 546200 189174
rect 546284 188938 546520 189174
rect 545964 188618 546200 188854
rect 546284 188618 546520 188854
rect 545964 170938 546200 171174
rect 546284 170938 546520 171174
rect 545964 170618 546200 170854
rect 546284 170618 546520 170854
rect 545964 152938 546200 153174
rect 546284 152938 546520 153174
rect 545964 152618 546200 152854
rect 546284 152618 546520 152854
rect 545964 134938 546200 135174
rect 546284 134938 546520 135174
rect 545964 134618 546200 134854
rect 546284 134618 546520 134854
rect 545964 116938 546200 117174
rect 546284 116938 546520 117174
rect 545964 116618 546200 116854
rect 546284 116618 546520 116854
rect 545964 98938 546200 99174
rect 546284 98938 546520 99174
rect 545964 98618 546200 98854
rect 546284 98618 546520 98854
rect 545964 80938 546200 81174
rect 546284 80938 546520 81174
rect 545964 80618 546200 80854
rect 546284 80618 546520 80854
rect 545964 62938 546200 63174
rect 546284 62938 546520 63174
rect 545964 62618 546200 62854
rect 546284 62618 546520 62854
rect 545964 44938 546200 45174
rect 546284 44938 546520 45174
rect 545964 44618 546200 44854
rect 546284 44618 546520 44854
rect 545964 26938 546200 27174
rect 546284 26938 546520 27174
rect 545964 26618 546200 26854
rect 546284 26618 546520 26854
rect 545964 8938 546200 9174
rect 546284 8938 546520 9174
rect 545964 8618 546200 8854
rect 546284 8618 546520 8854
rect 545964 -2052 546200 -1816
rect 546284 -2052 546520 -1816
rect 545964 -2372 546200 -2136
rect 546284 -2372 546520 -2136
rect 546924 444658 547160 444894
rect 547244 444658 547480 444894
rect 546924 444338 547160 444574
rect 547244 444338 547480 444574
rect 546924 426658 547160 426894
rect 547244 426658 547480 426894
rect 546924 426338 547160 426574
rect 547244 426338 547480 426574
rect 546924 408658 547160 408894
rect 547244 408658 547480 408894
rect 546924 408338 547160 408574
rect 547244 408338 547480 408574
rect 546924 390658 547160 390894
rect 547244 390658 547480 390894
rect 546924 390338 547160 390574
rect 547244 390338 547480 390574
rect 546924 372658 547160 372894
rect 547244 372658 547480 372894
rect 546924 372338 547160 372574
rect 547244 372338 547480 372574
rect 546924 354658 547160 354894
rect 547244 354658 547480 354894
rect 546924 354338 547160 354574
rect 547244 354338 547480 354574
rect 546924 336658 547160 336894
rect 547244 336658 547480 336894
rect 546924 336338 547160 336574
rect 547244 336338 547480 336574
rect 546924 318658 547160 318894
rect 547244 318658 547480 318894
rect 546924 318338 547160 318574
rect 547244 318338 547480 318574
rect 546924 300658 547160 300894
rect 547244 300658 547480 300894
rect 546924 300338 547160 300574
rect 547244 300338 547480 300574
rect 546924 282658 547160 282894
rect 547244 282658 547480 282894
rect 546924 282338 547160 282574
rect 547244 282338 547480 282574
rect 546924 264658 547160 264894
rect 547244 264658 547480 264894
rect 546924 264338 547160 264574
rect 547244 264338 547480 264574
rect 546924 246658 547160 246894
rect 547244 246658 547480 246894
rect 546924 246338 547160 246574
rect 547244 246338 547480 246574
rect 546924 228658 547160 228894
rect 547244 228658 547480 228894
rect 546924 228338 547160 228574
rect 547244 228338 547480 228574
rect 546924 210658 547160 210894
rect 547244 210658 547480 210894
rect 546924 210338 547160 210574
rect 547244 210338 547480 210574
rect 546924 192658 547160 192894
rect 547244 192658 547480 192894
rect 546924 192338 547160 192574
rect 547244 192338 547480 192574
rect 546924 174658 547160 174894
rect 547244 174658 547480 174894
rect 546924 174338 547160 174574
rect 547244 174338 547480 174574
rect 546924 156658 547160 156894
rect 547244 156658 547480 156894
rect 546924 156338 547160 156574
rect 547244 156338 547480 156574
rect 546924 138658 547160 138894
rect 547244 138658 547480 138894
rect 546924 138338 547160 138574
rect 547244 138338 547480 138574
rect 546924 120658 547160 120894
rect 547244 120658 547480 120894
rect 546924 120338 547160 120574
rect 547244 120338 547480 120574
rect 546924 102658 547160 102894
rect 547244 102658 547480 102894
rect 546924 102338 547160 102574
rect 547244 102338 547480 102574
rect 546924 84658 547160 84894
rect 547244 84658 547480 84894
rect 546924 84338 547160 84574
rect 547244 84338 547480 84574
rect 546924 66658 547160 66894
rect 547244 66658 547480 66894
rect 546924 66338 547160 66574
rect 547244 66338 547480 66574
rect 546924 48658 547160 48894
rect 547244 48658 547480 48894
rect 546924 48338 547160 48574
rect 547244 48338 547480 48574
rect 546924 30658 547160 30894
rect 547244 30658 547480 30894
rect 546924 30338 547160 30574
rect 547244 30338 547480 30574
rect 546924 12658 547160 12894
rect 547244 12658 547480 12894
rect 546924 12338 547160 12574
rect 547244 12338 547480 12574
rect 498186 -3012 498422 -2776
rect 498506 -3012 498742 -2776
rect 498186 -3332 498422 -3096
rect 498506 -3332 498742 -3096
rect 546924 -3012 547160 -2776
rect 547244 -3012 547480 -2776
rect 546924 -3332 547160 -3096
rect 547244 -3332 547480 -3096
rect 547884 448378 548120 448614
rect 548204 448378 548440 448614
rect 547884 448058 548120 448294
rect 548204 448058 548440 448294
rect 547884 430378 548120 430614
rect 548204 430378 548440 430614
rect 547884 430058 548120 430294
rect 548204 430058 548440 430294
rect 547884 412378 548120 412614
rect 548204 412378 548440 412614
rect 547884 412058 548120 412294
rect 548204 412058 548440 412294
rect 547884 394378 548120 394614
rect 548204 394378 548440 394614
rect 547884 394058 548120 394294
rect 548204 394058 548440 394294
rect 547884 376378 548120 376614
rect 548204 376378 548440 376614
rect 547884 376058 548120 376294
rect 548204 376058 548440 376294
rect 547884 358378 548120 358614
rect 548204 358378 548440 358614
rect 547884 358058 548120 358294
rect 548204 358058 548440 358294
rect 547884 340378 548120 340614
rect 548204 340378 548440 340614
rect 547884 340058 548120 340294
rect 548204 340058 548440 340294
rect 547884 322378 548120 322614
rect 548204 322378 548440 322614
rect 547884 322058 548120 322294
rect 548204 322058 548440 322294
rect 547884 304378 548120 304614
rect 548204 304378 548440 304614
rect 547884 304058 548120 304294
rect 548204 304058 548440 304294
rect 547884 286378 548120 286614
rect 548204 286378 548440 286614
rect 547884 286058 548120 286294
rect 548204 286058 548440 286294
rect 547884 268378 548120 268614
rect 548204 268378 548440 268614
rect 547884 268058 548120 268294
rect 548204 268058 548440 268294
rect 547884 250378 548120 250614
rect 548204 250378 548440 250614
rect 547884 250058 548120 250294
rect 548204 250058 548440 250294
rect 547884 232378 548120 232614
rect 548204 232378 548440 232614
rect 547884 232058 548120 232294
rect 548204 232058 548440 232294
rect 547884 214378 548120 214614
rect 548204 214378 548440 214614
rect 547884 214058 548120 214294
rect 548204 214058 548440 214294
rect 547884 196378 548120 196614
rect 548204 196378 548440 196614
rect 547884 196058 548120 196294
rect 548204 196058 548440 196294
rect 547884 178378 548120 178614
rect 548204 178378 548440 178614
rect 547884 178058 548120 178294
rect 548204 178058 548440 178294
rect 547884 160378 548120 160614
rect 548204 160378 548440 160614
rect 547884 160058 548120 160294
rect 548204 160058 548440 160294
rect 547884 142378 548120 142614
rect 548204 142378 548440 142614
rect 547884 142058 548120 142294
rect 548204 142058 548440 142294
rect 547884 124378 548120 124614
rect 548204 124378 548440 124614
rect 547884 124058 548120 124294
rect 548204 124058 548440 124294
rect 547884 106378 548120 106614
rect 548204 106378 548440 106614
rect 547884 106058 548120 106294
rect 548204 106058 548440 106294
rect 547884 88378 548120 88614
rect 548204 88378 548440 88614
rect 547884 88058 548120 88294
rect 548204 88058 548440 88294
rect 547884 70378 548120 70614
rect 548204 70378 548440 70614
rect 547884 70058 548120 70294
rect 548204 70058 548440 70294
rect 547884 52378 548120 52614
rect 548204 52378 548440 52614
rect 547884 52058 548120 52294
rect 548204 52058 548440 52294
rect 547884 34378 548120 34614
rect 548204 34378 548440 34614
rect 547884 34058 548120 34294
rect 548204 34058 548440 34294
rect 547884 16378 548120 16614
rect 548204 16378 548440 16614
rect 547884 16058 548120 16294
rect 548204 16058 548440 16294
rect 547884 -3972 548120 -3736
rect 548204 -3972 548440 -3736
rect 547884 -4292 548120 -4056
rect 548204 -4292 548440 -4056
<< metal5 >>
rect -4476 463972 548472 464004
rect -4476 463736 -4444 463972
rect -4208 463736 -4124 463972
rect -3888 463736 15906 463972
rect 16142 463736 16226 463972
rect 16462 463736 33906 463972
rect 34142 463736 34226 463972
rect 34462 463736 51906 463972
rect 52142 463736 52226 463972
rect 52462 463736 69906 463972
rect 70142 463736 70226 463972
rect 70462 463736 87906 463972
rect 88142 463736 88226 463972
rect 88462 463736 105906 463972
rect 106142 463736 106226 463972
rect 106462 463736 123906 463972
rect 124142 463736 124226 463972
rect 124462 463736 141906 463972
rect 142142 463736 142226 463972
rect 142462 463736 159906 463972
rect 160142 463736 160226 463972
rect 160462 463736 177906 463972
rect 178142 463736 178226 463972
rect 178462 463736 195906 463972
rect 196142 463736 196226 463972
rect 196462 463736 213906 463972
rect 214142 463736 214226 463972
rect 214462 463736 231906 463972
rect 232142 463736 232226 463972
rect 232462 463736 249906 463972
rect 250142 463736 250226 463972
rect 250462 463736 267906 463972
rect 268142 463736 268226 463972
rect 268462 463736 285906 463972
rect 286142 463736 286226 463972
rect 286462 463736 303906 463972
rect 304142 463736 304226 463972
rect 304462 463736 321906 463972
rect 322142 463736 322226 463972
rect 322462 463736 357906 463972
rect 358142 463736 358226 463972
rect 358462 463736 375906 463972
rect 376142 463736 376226 463972
rect 376462 463736 393906 463972
rect 394142 463736 394226 463972
rect 394462 463736 411906 463972
rect 412142 463736 412226 463972
rect 412462 463736 429906 463972
rect 430142 463736 430226 463972
rect 430462 463736 447906 463972
rect 448142 463736 448226 463972
rect 448462 463736 465906 463972
rect 466142 463736 466226 463972
rect 466462 463736 483906 463972
rect 484142 463736 484226 463972
rect 484462 463736 501906 463972
rect 502142 463736 502226 463972
rect 502462 463736 519906 463972
rect 520142 463736 520226 463972
rect 520462 463736 537906 463972
rect 538142 463736 538226 463972
rect 538462 463736 547884 463972
rect 548120 463736 548204 463972
rect 548440 463736 548472 463972
rect -4476 463652 548472 463736
rect -4476 463416 -4444 463652
rect -4208 463416 -4124 463652
rect -3888 463416 15906 463652
rect 16142 463416 16226 463652
rect 16462 463416 33906 463652
rect 34142 463416 34226 463652
rect 34462 463416 51906 463652
rect 52142 463416 52226 463652
rect 52462 463416 69906 463652
rect 70142 463416 70226 463652
rect 70462 463416 87906 463652
rect 88142 463416 88226 463652
rect 88462 463416 105906 463652
rect 106142 463416 106226 463652
rect 106462 463416 123906 463652
rect 124142 463416 124226 463652
rect 124462 463416 141906 463652
rect 142142 463416 142226 463652
rect 142462 463416 159906 463652
rect 160142 463416 160226 463652
rect 160462 463416 177906 463652
rect 178142 463416 178226 463652
rect 178462 463416 195906 463652
rect 196142 463416 196226 463652
rect 196462 463416 213906 463652
rect 214142 463416 214226 463652
rect 214462 463416 231906 463652
rect 232142 463416 232226 463652
rect 232462 463416 249906 463652
rect 250142 463416 250226 463652
rect 250462 463416 267906 463652
rect 268142 463416 268226 463652
rect 268462 463416 285906 463652
rect 286142 463416 286226 463652
rect 286462 463416 303906 463652
rect 304142 463416 304226 463652
rect 304462 463416 321906 463652
rect 322142 463416 322226 463652
rect 322462 463416 357906 463652
rect 358142 463416 358226 463652
rect 358462 463416 375906 463652
rect 376142 463416 376226 463652
rect 376462 463416 393906 463652
rect 394142 463416 394226 463652
rect 394462 463416 411906 463652
rect 412142 463416 412226 463652
rect 412462 463416 429906 463652
rect 430142 463416 430226 463652
rect 430462 463416 447906 463652
rect 448142 463416 448226 463652
rect 448462 463416 465906 463652
rect 466142 463416 466226 463652
rect 466462 463416 483906 463652
rect 484142 463416 484226 463652
rect 484462 463416 501906 463652
rect 502142 463416 502226 463652
rect 502462 463416 519906 463652
rect 520142 463416 520226 463652
rect 520462 463416 537906 463652
rect 538142 463416 538226 463652
rect 538462 463416 547884 463652
rect 548120 463416 548204 463652
rect 548440 463416 548472 463652
rect -4476 463384 548472 463416
rect -3516 463012 547512 463044
rect -3516 462776 -3484 463012
rect -3248 462776 -3164 463012
rect -2928 462776 12186 463012
rect 12422 462776 12506 463012
rect 12742 462776 30186 463012
rect 30422 462776 30506 463012
rect 30742 462776 48186 463012
rect 48422 462776 48506 463012
rect 48742 462776 66186 463012
rect 66422 462776 66506 463012
rect 66742 462776 84186 463012
rect 84422 462776 84506 463012
rect 84742 462776 102186 463012
rect 102422 462776 102506 463012
rect 102742 462776 120186 463012
rect 120422 462776 120506 463012
rect 120742 462776 138186 463012
rect 138422 462776 138506 463012
rect 138742 462776 156186 463012
rect 156422 462776 156506 463012
rect 156742 462776 174186 463012
rect 174422 462776 174506 463012
rect 174742 462776 192186 463012
rect 192422 462776 192506 463012
rect 192742 462776 210186 463012
rect 210422 462776 210506 463012
rect 210742 462776 228186 463012
rect 228422 462776 228506 463012
rect 228742 462776 246186 463012
rect 246422 462776 246506 463012
rect 246742 462776 264186 463012
rect 264422 462776 264506 463012
rect 264742 462776 282186 463012
rect 282422 462776 282506 463012
rect 282742 462776 300186 463012
rect 300422 462776 300506 463012
rect 300742 462776 318186 463012
rect 318422 462776 318506 463012
rect 318742 462776 354186 463012
rect 354422 462776 354506 463012
rect 354742 462776 372186 463012
rect 372422 462776 372506 463012
rect 372742 462776 390186 463012
rect 390422 462776 390506 463012
rect 390742 462776 408186 463012
rect 408422 462776 408506 463012
rect 408742 462776 426186 463012
rect 426422 462776 426506 463012
rect 426742 462776 444186 463012
rect 444422 462776 444506 463012
rect 444742 462776 462186 463012
rect 462422 462776 462506 463012
rect 462742 462776 480186 463012
rect 480422 462776 480506 463012
rect 480742 462776 498186 463012
rect 498422 462776 498506 463012
rect 498742 462776 516186 463012
rect 516422 462776 516506 463012
rect 516742 462776 534186 463012
rect 534422 462776 534506 463012
rect 534742 462776 546924 463012
rect 547160 462776 547244 463012
rect 547480 462776 547512 463012
rect -3516 462692 547512 462776
rect -3516 462456 -3484 462692
rect -3248 462456 -3164 462692
rect -2928 462456 12186 462692
rect 12422 462456 12506 462692
rect 12742 462456 30186 462692
rect 30422 462456 30506 462692
rect 30742 462456 48186 462692
rect 48422 462456 48506 462692
rect 48742 462456 66186 462692
rect 66422 462456 66506 462692
rect 66742 462456 84186 462692
rect 84422 462456 84506 462692
rect 84742 462456 102186 462692
rect 102422 462456 102506 462692
rect 102742 462456 120186 462692
rect 120422 462456 120506 462692
rect 120742 462456 138186 462692
rect 138422 462456 138506 462692
rect 138742 462456 156186 462692
rect 156422 462456 156506 462692
rect 156742 462456 174186 462692
rect 174422 462456 174506 462692
rect 174742 462456 192186 462692
rect 192422 462456 192506 462692
rect 192742 462456 210186 462692
rect 210422 462456 210506 462692
rect 210742 462456 228186 462692
rect 228422 462456 228506 462692
rect 228742 462456 246186 462692
rect 246422 462456 246506 462692
rect 246742 462456 264186 462692
rect 264422 462456 264506 462692
rect 264742 462456 282186 462692
rect 282422 462456 282506 462692
rect 282742 462456 300186 462692
rect 300422 462456 300506 462692
rect 300742 462456 318186 462692
rect 318422 462456 318506 462692
rect 318742 462456 354186 462692
rect 354422 462456 354506 462692
rect 354742 462456 372186 462692
rect 372422 462456 372506 462692
rect 372742 462456 390186 462692
rect 390422 462456 390506 462692
rect 390742 462456 408186 462692
rect 408422 462456 408506 462692
rect 408742 462456 426186 462692
rect 426422 462456 426506 462692
rect 426742 462456 444186 462692
rect 444422 462456 444506 462692
rect 444742 462456 462186 462692
rect 462422 462456 462506 462692
rect 462742 462456 480186 462692
rect 480422 462456 480506 462692
rect 480742 462456 498186 462692
rect 498422 462456 498506 462692
rect 498742 462456 516186 462692
rect 516422 462456 516506 462692
rect 516742 462456 534186 462692
rect 534422 462456 534506 462692
rect 534742 462456 546924 462692
rect 547160 462456 547244 462692
rect 547480 462456 547512 462692
rect -3516 462424 547512 462456
rect -2556 462052 546552 462084
rect -2556 461816 -2524 462052
rect -2288 461816 -2204 462052
rect -1968 461816 8466 462052
rect 8702 461816 8786 462052
rect 9022 461816 26466 462052
rect 26702 461816 26786 462052
rect 27022 461816 44466 462052
rect 44702 461816 44786 462052
rect 45022 461816 62466 462052
rect 62702 461816 62786 462052
rect 63022 461816 80466 462052
rect 80702 461816 80786 462052
rect 81022 461816 98466 462052
rect 98702 461816 98786 462052
rect 99022 461816 116466 462052
rect 116702 461816 116786 462052
rect 117022 461816 134466 462052
rect 134702 461816 134786 462052
rect 135022 461816 152466 462052
rect 152702 461816 152786 462052
rect 153022 461816 170466 462052
rect 170702 461816 170786 462052
rect 171022 461816 188466 462052
rect 188702 461816 188786 462052
rect 189022 461816 206466 462052
rect 206702 461816 206786 462052
rect 207022 461816 224466 462052
rect 224702 461816 224786 462052
rect 225022 461816 242466 462052
rect 242702 461816 242786 462052
rect 243022 461816 260466 462052
rect 260702 461816 260786 462052
rect 261022 461816 278466 462052
rect 278702 461816 278786 462052
rect 279022 461816 296466 462052
rect 296702 461816 296786 462052
rect 297022 461816 314466 462052
rect 314702 461816 314786 462052
rect 315022 461816 368466 462052
rect 368702 461816 368786 462052
rect 369022 461816 386466 462052
rect 386702 461816 386786 462052
rect 387022 461816 404466 462052
rect 404702 461816 404786 462052
rect 405022 461816 422466 462052
rect 422702 461816 422786 462052
rect 423022 461816 440466 462052
rect 440702 461816 440786 462052
rect 441022 461816 458466 462052
rect 458702 461816 458786 462052
rect 459022 461816 476466 462052
rect 476702 461816 476786 462052
rect 477022 461816 494466 462052
rect 494702 461816 494786 462052
rect 495022 461816 512466 462052
rect 512702 461816 512786 462052
rect 513022 461816 530466 462052
rect 530702 461816 530786 462052
rect 531022 461816 545964 462052
rect 546200 461816 546284 462052
rect 546520 461816 546552 462052
rect -2556 461732 546552 461816
rect -2556 461496 -2524 461732
rect -2288 461496 -2204 461732
rect -1968 461496 8466 461732
rect 8702 461496 8786 461732
rect 9022 461496 26466 461732
rect 26702 461496 26786 461732
rect 27022 461496 44466 461732
rect 44702 461496 44786 461732
rect 45022 461496 62466 461732
rect 62702 461496 62786 461732
rect 63022 461496 80466 461732
rect 80702 461496 80786 461732
rect 81022 461496 98466 461732
rect 98702 461496 98786 461732
rect 99022 461496 116466 461732
rect 116702 461496 116786 461732
rect 117022 461496 134466 461732
rect 134702 461496 134786 461732
rect 135022 461496 152466 461732
rect 152702 461496 152786 461732
rect 153022 461496 170466 461732
rect 170702 461496 170786 461732
rect 171022 461496 188466 461732
rect 188702 461496 188786 461732
rect 189022 461496 206466 461732
rect 206702 461496 206786 461732
rect 207022 461496 224466 461732
rect 224702 461496 224786 461732
rect 225022 461496 242466 461732
rect 242702 461496 242786 461732
rect 243022 461496 260466 461732
rect 260702 461496 260786 461732
rect 261022 461496 278466 461732
rect 278702 461496 278786 461732
rect 279022 461496 296466 461732
rect 296702 461496 296786 461732
rect 297022 461496 314466 461732
rect 314702 461496 314786 461732
rect 315022 461496 368466 461732
rect 368702 461496 368786 461732
rect 369022 461496 386466 461732
rect 386702 461496 386786 461732
rect 387022 461496 404466 461732
rect 404702 461496 404786 461732
rect 405022 461496 422466 461732
rect 422702 461496 422786 461732
rect 423022 461496 440466 461732
rect 440702 461496 440786 461732
rect 441022 461496 458466 461732
rect 458702 461496 458786 461732
rect 459022 461496 476466 461732
rect 476702 461496 476786 461732
rect 477022 461496 494466 461732
rect 494702 461496 494786 461732
rect 495022 461496 512466 461732
rect 512702 461496 512786 461732
rect 513022 461496 530466 461732
rect 530702 461496 530786 461732
rect 531022 461496 545964 461732
rect 546200 461496 546284 461732
rect 546520 461496 546552 461732
rect -2556 461464 546552 461496
rect -1596 461092 545592 461124
rect -1596 460856 -1564 461092
rect -1328 460856 -1244 461092
rect -1008 460856 4746 461092
rect 4982 460856 5066 461092
rect 5302 460856 22746 461092
rect 22982 460856 23066 461092
rect 23302 460856 40746 461092
rect 40982 460856 41066 461092
rect 41302 460856 58746 461092
rect 58982 460856 59066 461092
rect 59302 460856 76746 461092
rect 76982 460856 77066 461092
rect 77302 460856 94746 461092
rect 94982 460856 95066 461092
rect 95302 460856 112746 461092
rect 112982 460856 113066 461092
rect 113302 460856 130746 461092
rect 130982 460856 131066 461092
rect 131302 460856 148746 461092
rect 148982 460856 149066 461092
rect 149302 460856 166746 461092
rect 166982 460856 167066 461092
rect 167302 460856 184746 461092
rect 184982 460856 185066 461092
rect 185302 460856 202746 461092
rect 202982 460856 203066 461092
rect 203302 460856 220746 461092
rect 220982 460856 221066 461092
rect 221302 460856 238746 461092
rect 238982 460856 239066 461092
rect 239302 460856 256746 461092
rect 256982 460856 257066 461092
rect 257302 460856 274746 461092
rect 274982 460856 275066 461092
rect 275302 460856 292746 461092
rect 292982 460856 293066 461092
rect 293302 460856 310746 461092
rect 310982 460856 311066 461092
rect 311302 460856 328746 461092
rect 328982 460856 329066 461092
rect 329302 460856 364746 461092
rect 364982 460856 365066 461092
rect 365302 460856 382746 461092
rect 382982 460856 383066 461092
rect 383302 460856 400746 461092
rect 400982 460856 401066 461092
rect 401302 460856 418746 461092
rect 418982 460856 419066 461092
rect 419302 460856 436746 461092
rect 436982 460856 437066 461092
rect 437302 460856 454746 461092
rect 454982 460856 455066 461092
rect 455302 460856 472746 461092
rect 472982 460856 473066 461092
rect 473302 460856 490746 461092
rect 490982 460856 491066 461092
rect 491302 460856 508746 461092
rect 508982 460856 509066 461092
rect 509302 460856 526746 461092
rect 526982 460856 527066 461092
rect 527302 460856 545004 461092
rect 545240 460856 545324 461092
rect 545560 460856 545592 461092
rect -1596 460772 545592 460856
rect -1596 460536 -1564 460772
rect -1328 460536 -1244 460772
rect -1008 460536 4746 460772
rect 4982 460536 5066 460772
rect 5302 460536 22746 460772
rect 22982 460536 23066 460772
rect 23302 460536 40746 460772
rect 40982 460536 41066 460772
rect 41302 460536 58746 460772
rect 58982 460536 59066 460772
rect 59302 460536 76746 460772
rect 76982 460536 77066 460772
rect 77302 460536 94746 460772
rect 94982 460536 95066 460772
rect 95302 460536 112746 460772
rect 112982 460536 113066 460772
rect 113302 460536 130746 460772
rect 130982 460536 131066 460772
rect 131302 460536 148746 460772
rect 148982 460536 149066 460772
rect 149302 460536 166746 460772
rect 166982 460536 167066 460772
rect 167302 460536 184746 460772
rect 184982 460536 185066 460772
rect 185302 460536 202746 460772
rect 202982 460536 203066 460772
rect 203302 460536 220746 460772
rect 220982 460536 221066 460772
rect 221302 460536 238746 460772
rect 238982 460536 239066 460772
rect 239302 460536 256746 460772
rect 256982 460536 257066 460772
rect 257302 460536 274746 460772
rect 274982 460536 275066 460772
rect 275302 460536 292746 460772
rect 292982 460536 293066 460772
rect 293302 460536 310746 460772
rect 310982 460536 311066 460772
rect 311302 460536 328746 460772
rect 328982 460536 329066 460772
rect 329302 460536 364746 460772
rect 364982 460536 365066 460772
rect 365302 460536 382746 460772
rect 382982 460536 383066 460772
rect 383302 460536 400746 460772
rect 400982 460536 401066 460772
rect 401302 460536 418746 460772
rect 418982 460536 419066 460772
rect 419302 460536 436746 460772
rect 436982 460536 437066 460772
rect 437302 460536 454746 460772
rect 454982 460536 455066 460772
rect 455302 460536 472746 460772
rect 472982 460536 473066 460772
rect 473302 460536 490746 460772
rect 490982 460536 491066 460772
rect 491302 460536 508746 460772
rect 508982 460536 509066 460772
rect 509302 460536 526746 460772
rect 526982 460536 527066 460772
rect 527302 460536 545004 460772
rect 545240 460536 545324 460772
rect 545560 460536 545592 460772
rect -1596 460504 545592 460536
rect -4476 455454 548472 455486
rect -4476 455218 -1564 455454
rect -1328 455218 -1244 455454
rect -1008 455218 4746 455454
rect 4982 455218 5066 455454
rect 5302 455218 22746 455454
rect 22982 455218 23066 455454
rect 23302 455218 40746 455454
rect 40982 455218 41066 455454
rect 41302 455218 58746 455454
rect 58982 455218 59066 455454
rect 59302 455218 76746 455454
rect 76982 455218 77066 455454
rect 77302 455218 94746 455454
rect 94982 455218 95066 455454
rect 95302 455218 112746 455454
rect 112982 455218 113066 455454
rect 113302 455218 130746 455454
rect 130982 455218 131066 455454
rect 131302 455218 148746 455454
rect 148982 455218 149066 455454
rect 149302 455218 166746 455454
rect 166982 455218 167066 455454
rect 167302 455218 184746 455454
rect 184982 455218 185066 455454
rect 185302 455218 202746 455454
rect 202982 455218 203066 455454
rect 203302 455218 220746 455454
rect 220982 455218 221066 455454
rect 221302 455218 238746 455454
rect 238982 455218 239066 455454
rect 239302 455218 256746 455454
rect 256982 455218 257066 455454
rect 257302 455218 274746 455454
rect 274982 455218 275066 455454
rect 275302 455218 292746 455454
rect 292982 455218 293066 455454
rect 293302 455218 310746 455454
rect 310982 455218 311066 455454
rect 311302 455218 328746 455454
rect 328982 455218 329066 455454
rect 329302 455218 346746 455454
rect 346982 455218 347066 455454
rect 347302 455218 364746 455454
rect 364982 455218 365066 455454
rect 365302 455218 382746 455454
rect 382982 455218 383066 455454
rect 383302 455218 400746 455454
rect 400982 455218 401066 455454
rect 401302 455218 418746 455454
rect 418982 455218 419066 455454
rect 419302 455218 436746 455454
rect 436982 455218 437066 455454
rect 437302 455218 454746 455454
rect 454982 455218 455066 455454
rect 455302 455218 472746 455454
rect 472982 455218 473066 455454
rect 473302 455218 490746 455454
rect 490982 455218 491066 455454
rect 491302 455218 508746 455454
rect 508982 455218 509066 455454
rect 509302 455218 526746 455454
rect 526982 455218 527066 455454
rect 527302 455218 545004 455454
rect 545240 455218 545324 455454
rect 545560 455218 548472 455454
rect -4476 455134 548472 455218
rect -4476 454898 -1564 455134
rect -1328 454898 -1244 455134
rect -1008 454898 4746 455134
rect 4982 454898 5066 455134
rect 5302 454898 22746 455134
rect 22982 454898 23066 455134
rect 23302 454898 40746 455134
rect 40982 454898 41066 455134
rect 41302 454898 58746 455134
rect 58982 454898 59066 455134
rect 59302 454898 76746 455134
rect 76982 454898 77066 455134
rect 77302 454898 94746 455134
rect 94982 454898 95066 455134
rect 95302 454898 112746 455134
rect 112982 454898 113066 455134
rect 113302 454898 130746 455134
rect 130982 454898 131066 455134
rect 131302 454898 148746 455134
rect 148982 454898 149066 455134
rect 149302 454898 166746 455134
rect 166982 454898 167066 455134
rect 167302 454898 184746 455134
rect 184982 454898 185066 455134
rect 185302 454898 202746 455134
rect 202982 454898 203066 455134
rect 203302 454898 220746 455134
rect 220982 454898 221066 455134
rect 221302 454898 238746 455134
rect 238982 454898 239066 455134
rect 239302 454898 256746 455134
rect 256982 454898 257066 455134
rect 257302 454898 274746 455134
rect 274982 454898 275066 455134
rect 275302 454898 292746 455134
rect 292982 454898 293066 455134
rect 293302 454898 310746 455134
rect 310982 454898 311066 455134
rect 311302 454898 328746 455134
rect 328982 454898 329066 455134
rect 329302 454898 346746 455134
rect 346982 454898 347066 455134
rect 347302 454898 364746 455134
rect 364982 454898 365066 455134
rect 365302 454898 382746 455134
rect 382982 454898 383066 455134
rect 383302 454898 400746 455134
rect 400982 454898 401066 455134
rect 401302 454898 418746 455134
rect 418982 454898 419066 455134
rect 419302 454898 436746 455134
rect 436982 454898 437066 455134
rect 437302 454898 454746 455134
rect 454982 454898 455066 455134
rect 455302 454898 472746 455134
rect 472982 454898 473066 455134
rect 473302 454898 490746 455134
rect 490982 454898 491066 455134
rect 491302 454898 508746 455134
rect 508982 454898 509066 455134
rect 509302 454898 526746 455134
rect 526982 454898 527066 455134
rect 527302 454898 545004 455134
rect 545240 454898 545324 455134
rect 545560 454898 548472 455134
rect -4476 454866 548472 454898
rect -4476 448614 548472 448646
rect -4476 448378 -4444 448614
rect -4208 448378 -4124 448614
rect -3888 448378 15906 448614
rect 16142 448378 16226 448614
rect 16462 448378 33906 448614
rect 34142 448378 34226 448614
rect 34462 448378 51906 448614
rect 52142 448378 52226 448614
rect 52462 448378 69906 448614
rect 70142 448378 70226 448614
rect 70462 448378 87906 448614
rect 88142 448378 88226 448614
rect 88462 448378 105906 448614
rect 106142 448378 106226 448614
rect 106462 448378 123906 448614
rect 124142 448378 124226 448614
rect 124462 448378 141906 448614
rect 142142 448378 142226 448614
rect 142462 448378 159906 448614
rect 160142 448378 160226 448614
rect 160462 448378 177906 448614
rect 178142 448378 178226 448614
rect 178462 448378 195906 448614
rect 196142 448378 196226 448614
rect 196462 448378 213906 448614
rect 214142 448378 214226 448614
rect 214462 448378 231906 448614
rect 232142 448378 232226 448614
rect 232462 448378 249906 448614
rect 250142 448378 250226 448614
rect 250462 448378 267906 448614
rect 268142 448378 268226 448614
rect 268462 448378 285906 448614
rect 286142 448378 286226 448614
rect 286462 448378 303906 448614
rect 304142 448378 304226 448614
rect 304462 448378 321906 448614
rect 322142 448378 322226 448614
rect 322462 448378 339906 448614
rect 340142 448378 340226 448614
rect 340462 448378 357906 448614
rect 358142 448378 358226 448614
rect 358462 448378 375906 448614
rect 376142 448378 376226 448614
rect 376462 448378 393906 448614
rect 394142 448378 394226 448614
rect 394462 448378 411906 448614
rect 412142 448378 412226 448614
rect 412462 448378 429906 448614
rect 430142 448378 430226 448614
rect 430462 448378 447906 448614
rect 448142 448378 448226 448614
rect 448462 448378 465906 448614
rect 466142 448378 466226 448614
rect 466462 448378 483906 448614
rect 484142 448378 484226 448614
rect 484462 448378 501906 448614
rect 502142 448378 502226 448614
rect 502462 448378 519906 448614
rect 520142 448378 520226 448614
rect 520462 448378 537906 448614
rect 538142 448378 538226 448614
rect 538462 448378 547884 448614
rect 548120 448378 548204 448614
rect 548440 448378 548472 448614
rect -4476 448294 548472 448378
rect -4476 448058 -4444 448294
rect -4208 448058 -4124 448294
rect -3888 448058 15906 448294
rect 16142 448058 16226 448294
rect 16462 448058 33906 448294
rect 34142 448058 34226 448294
rect 34462 448058 51906 448294
rect 52142 448058 52226 448294
rect 52462 448058 69906 448294
rect 70142 448058 70226 448294
rect 70462 448058 87906 448294
rect 88142 448058 88226 448294
rect 88462 448058 105906 448294
rect 106142 448058 106226 448294
rect 106462 448058 123906 448294
rect 124142 448058 124226 448294
rect 124462 448058 141906 448294
rect 142142 448058 142226 448294
rect 142462 448058 159906 448294
rect 160142 448058 160226 448294
rect 160462 448058 177906 448294
rect 178142 448058 178226 448294
rect 178462 448058 195906 448294
rect 196142 448058 196226 448294
rect 196462 448058 213906 448294
rect 214142 448058 214226 448294
rect 214462 448058 231906 448294
rect 232142 448058 232226 448294
rect 232462 448058 249906 448294
rect 250142 448058 250226 448294
rect 250462 448058 267906 448294
rect 268142 448058 268226 448294
rect 268462 448058 285906 448294
rect 286142 448058 286226 448294
rect 286462 448058 303906 448294
rect 304142 448058 304226 448294
rect 304462 448058 321906 448294
rect 322142 448058 322226 448294
rect 322462 448058 339906 448294
rect 340142 448058 340226 448294
rect 340462 448058 357906 448294
rect 358142 448058 358226 448294
rect 358462 448058 375906 448294
rect 376142 448058 376226 448294
rect 376462 448058 393906 448294
rect 394142 448058 394226 448294
rect 394462 448058 411906 448294
rect 412142 448058 412226 448294
rect 412462 448058 429906 448294
rect 430142 448058 430226 448294
rect 430462 448058 447906 448294
rect 448142 448058 448226 448294
rect 448462 448058 465906 448294
rect 466142 448058 466226 448294
rect 466462 448058 483906 448294
rect 484142 448058 484226 448294
rect 484462 448058 501906 448294
rect 502142 448058 502226 448294
rect 502462 448058 519906 448294
rect 520142 448058 520226 448294
rect 520462 448058 537906 448294
rect 538142 448058 538226 448294
rect 538462 448058 547884 448294
rect 548120 448058 548204 448294
rect 548440 448058 548472 448294
rect -4476 448026 548472 448058
rect -4476 444894 548472 444926
rect -4476 444658 -3484 444894
rect -3248 444658 -3164 444894
rect -2928 444658 12186 444894
rect 12422 444658 12506 444894
rect 12742 444658 30186 444894
rect 30422 444658 30506 444894
rect 30742 444658 48186 444894
rect 48422 444658 48506 444894
rect 48742 444658 66186 444894
rect 66422 444658 66506 444894
rect 66742 444658 84186 444894
rect 84422 444658 84506 444894
rect 84742 444658 102186 444894
rect 102422 444658 102506 444894
rect 102742 444658 120186 444894
rect 120422 444658 120506 444894
rect 120742 444658 138186 444894
rect 138422 444658 138506 444894
rect 138742 444658 156186 444894
rect 156422 444658 156506 444894
rect 156742 444658 174186 444894
rect 174422 444658 174506 444894
rect 174742 444658 192186 444894
rect 192422 444658 192506 444894
rect 192742 444658 210186 444894
rect 210422 444658 210506 444894
rect 210742 444658 228186 444894
rect 228422 444658 228506 444894
rect 228742 444658 246186 444894
rect 246422 444658 246506 444894
rect 246742 444658 264186 444894
rect 264422 444658 264506 444894
rect 264742 444658 282186 444894
rect 282422 444658 282506 444894
rect 282742 444658 300186 444894
rect 300422 444658 300506 444894
rect 300742 444658 318186 444894
rect 318422 444658 318506 444894
rect 318742 444658 336186 444894
rect 336422 444658 336506 444894
rect 336742 444658 354186 444894
rect 354422 444658 354506 444894
rect 354742 444658 372186 444894
rect 372422 444658 372506 444894
rect 372742 444658 390186 444894
rect 390422 444658 390506 444894
rect 390742 444658 408186 444894
rect 408422 444658 408506 444894
rect 408742 444658 426186 444894
rect 426422 444658 426506 444894
rect 426742 444658 444186 444894
rect 444422 444658 444506 444894
rect 444742 444658 462186 444894
rect 462422 444658 462506 444894
rect 462742 444658 480186 444894
rect 480422 444658 480506 444894
rect 480742 444658 498186 444894
rect 498422 444658 498506 444894
rect 498742 444658 516186 444894
rect 516422 444658 516506 444894
rect 516742 444658 534186 444894
rect 534422 444658 534506 444894
rect 534742 444658 546924 444894
rect 547160 444658 547244 444894
rect 547480 444658 548472 444894
rect -4476 444574 548472 444658
rect -4476 444338 -3484 444574
rect -3248 444338 -3164 444574
rect -2928 444338 12186 444574
rect 12422 444338 12506 444574
rect 12742 444338 30186 444574
rect 30422 444338 30506 444574
rect 30742 444338 48186 444574
rect 48422 444338 48506 444574
rect 48742 444338 66186 444574
rect 66422 444338 66506 444574
rect 66742 444338 84186 444574
rect 84422 444338 84506 444574
rect 84742 444338 102186 444574
rect 102422 444338 102506 444574
rect 102742 444338 120186 444574
rect 120422 444338 120506 444574
rect 120742 444338 138186 444574
rect 138422 444338 138506 444574
rect 138742 444338 156186 444574
rect 156422 444338 156506 444574
rect 156742 444338 174186 444574
rect 174422 444338 174506 444574
rect 174742 444338 192186 444574
rect 192422 444338 192506 444574
rect 192742 444338 210186 444574
rect 210422 444338 210506 444574
rect 210742 444338 228186 444574
rect 228422 444338 228506 444574
rect 228742 444338 246186 444574
rect 246422 444338 246506 444574
rect 246742 444338 264186 444574
rect 264422 444338 264506 444574
rect 264742 444338 282186 444574
rect 282422 444338 282506 444574
rect 282742 444338 300186 444574
rect 300422 444338 300506 444574
rect 300742 444338 318186 444574
rect 318422 444338 318506 444574
rect 318742 444338 336186 444574
rect 336422 444338 336506 444574
rect 336742 444338 354186 444574
rect 354422 444338 354506 444574
rect 354742 444338 372186 444574
rect 372422 444338 372506 444574
rect 372742 444338 390186 444574
rect 390422 444338 390506 444574
rect 390742 444338 408186 444574
rect 408422 444338 408506 444574
rect 408742 444338 426186 444574
rect 426422 444338 426506 444574
rect 426742 444338 444186 444574
rect 444422 444338 444506 444574
rect 444742 444338 462186 444574
rect 462422 444338 462506 444574
rect 462742 444338 480186 444574
rect 480422 444338 480506 444574
rect 480742 444338 498186 444574
rect 498422 444338 498506 444574
rect 498742 444338 516186 444574
rect 516422 444338 516506 444574
rect 516742 444338 534186 444574
rect 534422 444338 534506 444574
rect 534742 444338 546924 444574
rect 547160 444338 547244 444574
rect 547480 444338 548472 444574
rect -4476 444306 548472 444338
rect -4476 441174 548472 441206
rect -4476 440938 -2524 441174
rect -2288 440938 -2204 441174
rect -1968 440938 8466 441174
rect 8702 440938 8786 441174
rect 9022 440938 26466 441174
rect 26702 440938 26786 441174
rect 27022 440938 44466 441174
rect 44702 440938 44786 441174
rect 45022 440938 62466 441174
rect 62702 440938 62786 441174
rect 63022 440938 80466 441174
rect 80702 440938 80786 441174
rect 81022 440938 98466 441174
rect 98702 440938 98786 441174
rect 99022 440938 116466 441174
rect 116702 440938 116786 441174
rect 117022 440938 134466 441174
rect 134702 440938 134786 441174
rect 135022 440938 152466 441174
rect 152702 440938 152786 441174
rect 153022 440938 170466 441174
rect 170702 440938 170786 441174
rect 171022 440938 188466 441174
rect 188702 440938 188786 441174
rect 189022 440938 206466 441174
rect 206702 440938 206786 441174
rect 207022 440938 224466 441174
rect 224702 440938 224786 441174
rect 225022 440938 242466 441174
rect 242702 440938 242786 441174
rect 243022 440938 260466 441174
rect 260702 440938 260786 441174
rect 261022 440938 278466 441174
rect 278702 440938 278786 441174
rect 279022 440938 296466 441174
rect 296702 440938 296786 441174
rect 297022 440938 314466 441174
rect 314702 440938 314786 441174
rect 315022 440938 332466 441174
rect 332702 440938 332786 441174
rect 333022 440938 350466 441174
rect 350702 440938 350786 441174
rect 351022 440938 368466 441174
rect 368702 440938 368786 441174
rect 369022 440938 386466 441174
rect 386702 440938 386786 441174
rect 387022 440938 404466 441174
rect 404702 440938 404786 441174
rect 405022 440938 422466 441174
rect 422702 440938 422786 441174
rect 423022 440938 440466 441174
rect 440702 440938 440786 441174
rect 441022 440938 458466 441174
rect 458702 440938 458786 441174
rect 459022 440938 476466 441174
rect 476702 440938 476786 441174
rect 477022 440938 494466 441174
rect 494702 440938 494786 441174
rect 495022 440938 512466 441174
rect 512702 440938 512786 441174
rect 513022 440938 530466 441174
rect 530702 440938 530786 441174
rect 531022 440938 545964 441174
rect 546200 440938 546284 441174
rect 546520 440938 548472 441174
rect -4476 440854 548472 440938
rect -4476 440618 -2524 440854
rect -2288 440618 -2204 440854
rect -1968 440618 8466 440854
rect 8702 440618 8786 440854
rect 9022 440618 26466 440854
rect 26702 440618 26786 440854
rect 27022 440618 44466 440854
rect 44702 440618 44786 440854
rect 45022 440618 62466 440854
rect 62702 440618 62786 440854
rect 63022 440618 80466 440854
rect 80702 440618 80786 440854
rect 81022 440618 98466 440854
rect 98702 440618 98786 440854
rect 99022 440618 116466 440854
rect 116702 440618 116786 440854
rect 117022 440618 134466 440854
rect 134702 440618 134786 440854
rect 135022 440618 152466 440854
rect 152702 440618 152786 440854
rect 153022 440618 170466 440854
rect 170702 440618 170786 440854
rect 171022 440618 188466 440854
rect 188702 440618 188786 440854
rect 189022 440618 206466 440854
rect 206702 440618 206786 440854
rect 207022 440618 224466 440854
rect 224702 440618 224786 440854
rect 225022 440618 242466 440854
rect 242702 440618 242786 440854
rect 243022 440618 260466 440854
rect 260702 440618 260786 440854
rect 261022 440618 278466 440854
rect 278702 440618 278786 440854
rect 279022 440618 296466 440854
rect 296702 440618 296786 440854
rect 297022 440618 314466 440854
rect 314702 440618 314786 440854
rect 315022 440618 332466 440854
rect 332702 440618 332786 440854
rect 333022 440618 350466 440854
rect 350702 440618 350786 440854
rect 351022 440618 368466 440854
rect 368702 440618 368786 440854
rect 369022 440618 386466 440854
rect 386702 440618 386786 440854
rect 387022 440618 404466 440854
rect 404702 440618 404786 440854
rect 405022 440618 422466 440854
rect 422702 440618 422786 440854
rect 423022 440618 440466 440854
rect 440702 440618 440786 440854
rect 441022 440618 458466 440854
rect 458702 440618 458786 440854
rect 459022 440618 476466 440854
rect 476702 440618 476786 440854
rect 477022 440618 494466 440854
rect 494702 440618 494786 440854
rect 495022 440618 512466 440854
rect 512702 440618 512786 440854
rect 513022 440618 530466 440854
rect 530702 440618 530786 440854
rect 531022 440618 545964 440854
rect 546200 440618 546284 440854
rect 546520 440618 548472 440854
rect -4476 440586 548472 440618
rect -4476 437454 548472 437486
rect -4476 437218 -1564 437454
rect -1328 437218 -1244 437454
rect -1008 437218 4746 437454
rect 4982 437218 5066 437454
rect 5302 437218 22746 437454
rect 22982 437218 23066 437454
rect 23302 437218 40746 437454
rect 40982 437218 41066 437454
rect 41302 437218 58746 437454
rect 58982 437218 59066 437454
rect 59302 437218 76746 437454
rect 76982 437218 77066 437454
rect 77302 437218 94746 437454
rect 94982 437218 95066 437454
rect 95302 437218 112746 437454
rect 112982 437218 113066 437454
rect 113302 437218 130746 437454
rect 130982 437218 131066 437454
rect 131302 437218 148746 437454
rect 148982 437218 149066 437454
rect 149302 437218 166746 437454
rect 166982 437218 167066 437454
rect 167302 437218 184746 437454
rect 184982 437218 185066 437454
rect 185302 437218 202746 437454
rect 202982 437218 203066 437454
rect 203302 437218 220746 437454
rect 220982 437218 221066 437454
rect 221302 437218 238746 437454
rect 238982 437218 239066 437454
rect 239302 437218 256746 437454
rect 256982 437218 257066 437454
rect 257302 437218 274746 437454
rect 274982 437218 275066 437454
rect 275302 437218 292746 437454
rect 292982 437218 293066 437454
rect 293302 437218 310746 437454
rect 310982 437218 311066 437454
rect 311302 437218 328746 437454
rect 328982 437218 329066 437454
rect 329302 437218 346746 437454
rect 346982 437218 347066 437454
rect 347302 437218 364746 437454
rect 364982 437218 365066 437454
rect 365302 437218 382746 437454
rect 382982 437218 383066 437454
rect 383302 437218 400746 437454
rect 400982 437218 401066 437454
rect 401302 437218 418746 437454
rect 418982 437218 419066 437454
rect 419302 437218 436746 437454
rect 436982 437218 437066 437454
rect 437302 437218 454746 437454
rect 454982 437218 455066 437454
rect 455302 437218 472746 437454
rect 472982 437218 473066 437454
rect 473302 437218 490746 437454
rect 490982 437218 491066 437454
rect 491302 437218 508746 437454
rect 508982 437218 509066 437454
rect 509302 437218 526746 437454
rect 526982 437218 527066 437454
rect 527302 437218 545004 437454
rect 545240 437218 545324 437454
rect 545560 437218 548472 437454
rect -4476 437134 548472 437218
rect -4476 436898 -1564 437134
rect -1328 436898 -1244 437134
rect -1008 436898 4746 437134
rect 4982 436898 5066 437134
rect 5302 436898 22746 437134
rect 22982 436898 23066 437134
rect 23302 436898 40746 437134
rect 40982 436898 41066 437134
rect 41302 436898 58746 437134
rect 58982 436898 59066 437134
rect 59302 436898 76746 437134
rect 76982 436898 77066 437134
rect 77302 436898 94746 437134
rect 94982 436898 95066 437134
rect 95302 436898 112746 437134
rect 112982 436898 113066 437134
rect 113302 436898 130746 437134
rect 130982 436898 131066 437134
rect 131302 436898 148746 437134
rect 148982 436898 149066 437134
rect 149302 436898 166746 437134
rect 166982 436898 167066 437134
rect 167302 436898 184746 437134
rect 184982 436898 185066 437134
rect 185302 436898 202746 437134
rect 202982 436898 203066 437134
rect 203302 436898 220746 437134
rect 220982 436898 221066 437134
rect 221302 436898 238746 437134
rect 238982 436898 239066 437134
rect 239302 436898 256746 437134
rect 256982 436898 257066 437134
rect 257302 436898 274746 437134
rect 274982 436898 275066 437134
rect 275302 436898 292746 437134
rect 292982 436898 293066 437134
rect 293302 436898 310746 437134
rect 310982 436898 311066 437134
rect 311302 436898 328746 437134
rect 328982 436898 329066 437134
rect 329302 436898 346746 437134
rect 346982 436898 347066 437134
rect 347302 436898 364746 437134
rect 364982 436898 365066 437134
rect 365302 436898 382746 437134
rect 382982 436898 383066 437134
rect 383302 436898 400746 437134
rect 400982 436898 401066 437134
rect 401302 436898 418746 437134
rect 418982 436898 419066 437134
rect 419302 436898 436746 437134
rect 436982 436898 437066 437134
rect 437302 436898 454746 437134
rect 454982 436898 455066 437134
rect 455302 436898 472746 437134
rect 472982 436898 473066 437134
rect 473302 436898 490746 437134
rect 490982 436898 491066 437134
rect 491302 436898 508746 437134
rect 508982 436898 509066 437134
rect 509302 436898 526746 437134
rect 526982 436898 527066 437134
rect 527302 436898 545004 437134
rect 545240 436898 545324 437134
rect 545560 436898 548472 437134
rect -4476 436866 548472 436898
rect -4476 430614 548472 430646
rect -4476 430378 -4444 430614
rect -4208 430378 -4124 430614
rect -3888 430378 15906 430614
rect 16142 430378 16226 430614
rect 16462 430378 33906 430614
rect 34142 430378 34226 430614
rect 34462 430378 51906 430614
rect 52142 430378 52226 430614
rect 52462 430378 69906 430614
rect 70142 430378 70226 430614
rect 70462 430378 87906 430614
rect 88142 430378 88226 430614
rect 88462 430378 105906 430614
rect 106142 430378 106226 430614
rect 106462 430378 123906 430614
rect 124142 430378 124226 430614
rect 124462 430378 141906 430614
rect 142142 430378 142226 430614
rect 142462 430378 159906 430614
rect 160142 430378 160226 430614
rect 160462 430378 177906 430614
rect 178142 430378 178226 430614
rect 178462 430378 195906 430614
rect 196142 430378 196226 430614
rect 196462 430378 213906 430614
rect 214142 430378 214226 430614
rect 214462 430378 231906 430614
rect 232142 430378 232226 430614
rect 232462 430378 249906 430614
rect 250142 430378 250226 430614
rect 250462 430378 267906 430614
rect 268142 430378 268226 430614
rect 268462 430378 285906 430614
rect 286142 430378 286226 430614
rect 286462 430378 303906 430614
rect 304142 430378 304226 430614
rect 304462 430378 321906 430614
rect 322142 430378 322226 430614
rect 322462 430378 339906 430614
rect 340142 430378 340226 430614
rect 340462 430378 357906 430614
rect 358142 430378 358226 430614
rect 358462 430378 375906 430614
rect 376142 430378 376226 430614
rect 376462 430378 393906 430614
rect 394142 430378 394226 430614
rect 394462 430378 411906 430614
rect 412142 430378 412226 430614
rect 412462 430378 429906 430614
rect 430142 430378 430226 430614
rect 430462 430378 447906 430614
rect 448142 430378 448226 430614
rect 448462 430378 465906 430614
rect 466142 430378 466226 430614
rect 466462 430378 483906 430614
rect 484142 430378 484226 430614
rect 484462 430378 501906 430614
rect 502142 430378 502226 430614
rect 502462 430378 519906 430614
rect 520142 430378 520226 430614
rect 520462 430378 537906 430614
rect 538142 430378 538226 430614
rect 538462 430378 547884 430614
rect 548120 430378 548204 430614
rect 548440 430378 548472 430614
rect -4476 430294 548472 430378
rect -4476 430058 -4444 430294
rect -4208 430058 -4124 430294
rect -3888 430058 15906 430294
rect 16142 430058 16226 430294
rect 16462 430058 33906 430294
rect 34142 430058 34226 430294
rect 34462 430058 51906 430294
rect 52142 430058 52226 430294
rect 52462 430058 69906 430294
rect 70142 430058 70226 430294
rect 70462 430058 87906 430294
rect 88142 430058 88226 430294
rect 88462 430058 105906 430294
rect 106142 430058 106226 430294
rect 106462 430058 123906 430294
rect 124142 430058 124226 430294
rect 124462 430058 141906 430294
rect 142142 430058 142226 430294
rect 142462 430058 159906 430294
rect 160142 430058 160226 430294
rect 160462 430058 177906 430294
rect 178142 430058 178226 430294
rect 178462 430058 195906 430294
rect 196142 430058 196226 430294
rect 196462 430058 213906 430294
rect 214142 430058 214226 430294
rect 214462 430058 231906 430294
rect 232142 430058 232226 430294
rect 232462 430058 249906 430294
rect 250142 430058 250226 430294
rect 250462 430058 267906 430294
rect 268142 430058 268226 430294
rect 268462 430058 285906 430294
rect 286142 430058 286226 430294
rect 286462 430058 303906 430294
rect 304142 430058 304226 430294
rect 304462 430058 321906 430294
rect 322142 430058 322226 430294
rect 322462 430058 339906 430294
rect 340142 430058 340226 430294
rect 340462 430058 357906 430294
rect 358142 430058 358226 430294
rect 358462 430058 375906 430294
rect 376142 430058 376226 430294
rect 376462 430058 393906 430294
rect 394142 430058 394226 430294
rect 394462 430058 411906 430294
rect 412142 430058 412226 430294
rect 412462 430058 429906 430294
rect 430142 430058 430226 430294
rect 430462 430058 447906 430294
rect 448142 430058 448226 430294
rect 448462 430058 465906 430294
rect 466142 430058 466226 430294
rect 466462 430058 483906 430294
rect 484142 430058 484226 430294
rect 484462 430058 501906 430294
rect 502142 430058 502226 430294
rect 502462 430058 519906 430294
rect 520142 430058 520226 430294
rect 520462 430058 537906 430294
rect 538142 430058 538226 430294
rect 538462 430058 547884 430294
rect 548120 430058 548204 430294
rect 548440 430058 548472 430294
rect -4476 430026 548472 430058
rect -4476 426894 548472 426926
rect -4476 426658 -3484 426894
rect -3248 426658 -3164 426894
rect -2928 426658 12186 426894
rect 12422 426658 12506 426894
rect 12742 426658 30186 426894
rect 30422 426658 30506 426894
rect 30742 426658 48186 426894
rect 48422 426658 48506 426894
rect 48742 426658 66186 426894
rect 66422 426658 66506 426894
rect 66742 426658 84186 426894
rect 84422 426658 84506 426894
rect 84742 426658 102186 426894
rect 102422 426658 102506 426894
rect 102742 426658 120186 426894
rect 120422 426658 120506 426894
rect 120742 426658 138186 426894
rect 138422 426658 138506 426894
rect 138742 426658 156186 426894
rect 156422 426658 156506 426894
rect 156742 426658 174186 426894
rect 174422 426658 174506 426894
rect 174742 426658 192186 426894
rect 192422 426658 192506 426894
rect 192742 426658 210186 426894
rect 210422 426658 210506 426894
rect 210742 426658 228186 426894
rect 228422 426658 228506 426894
rect 228742 426658 246186 426894
rect 246422 426658 246506 426894
rect 246742 426658 264186 426894
rect 264422 426658 264506 426894
rect 264742 426658 282186 426894
rect 282422 426658 282506 426894
rect 282742 426658 300186 426894
rect 300422 426658 300506 426894
rect 300742 426658 318186 426894
rect 318422 426658 318506 426894
rect 318742 426658 336186 426894
rect 336422 426658 336506 426894
rect 336742 426658 354186 426894
rect 354422 426658 354506 426894
rect 354742 426658 372186 426894
rect 372422 426658 372506 426894
rect 372742 426658 390186 426894
rect 390422 426658 390506 426894
rect 390742 426658 408186 426894
rect 408422 426658 408506 426894
rect 408742 426658 426186 426894
rect 426422 426658 426506 426894
rect 426742 426658 444186 426894
rect 444422 426658 444506 426894
rect 444742 426658 462186 426894
rect 462422 426658 462506 426894
rect 462742 426658 480186 426894
rect 480422 426658 480506 426894
rect 480742 426658 498186 426894
rect 498422 426658 498506 426894
rect 498742 426658 516186 426894
rect 516422 426658 516506 426894
rect 516742 426658 534186 426894
rect 534422 426658 534506 426894
rect 534742 426658 546924 426894
rect 547160 426658 547244 426894
rect 547480 426658 548472 426894
rect -4476 426574 548472 426658
rect -4476 426338 -3484 426574
rect -3248 426338 -3164 426574
rect -2928 426338 12186 426574
rect 12422 426338 12506 426574
rect 12742 426338 30186 426574
rect 30422 426338 30506 426574
rect 30742 426338 48186 426574
rect 48422 426338 48506 426574
rect 48742 426338 66186 426574
rect 66422 426338 66506 426574
rect 66742 426338 84186 426574
rect 84422 426338 84506 426574
rect 84742 426338 102186 426574
rect 102422 426338 102506 426574
rect 102742 426338 120186 426574
rect 120422 426338 120506 426574
rect 120742 426338 138186 426574
rect 138422 426338 138506 426574
rect 138742 426338 156186 426574
rect 156422 426338 156506 426574
rect 156742 426338 174186 426574
rect 174422 426338 174506 426574
rect 174742 426338 192186 426574
rect 192422 426338 192506 426574
rect 192742 426338 210186 426574
rect 210422 426338 210506 426574
rect 210742 426338 228186 426574
rect 228422 426338 228506 426574
rect 228742 426338 246186 426574
rect 246422 426338 246506 426574
rect 246742 426338 264186 426574
rect 264422 426338 264506 426574
rect 264742 426338 282186 426574
rect 282422 426338 282506 426574
rect 282742 426338 300186 426574
rect 300422 426338 300506 426574
rect 300742 426338 318186 426574
rect 318422 426338 318506 426574
rect 318742 426338 336186 426574
rect 336422 426338 336506 426574
rect 336742 426338 354186 426574
rect 354422 426338 354506 426574
rect 354742 426338 372186 426574
rect 372422 426338 372506 426574
rect 372742 426338 390186 426574
rect 390422 426338 390506 426574
rect 390742 426338 408186 426574
rect 408422 426338 408506 426574
rect 408742 426338 426186 426574
rect 426422 426338 426506 426574
rect 426742 426338 444186 426574
rect 444422 426338 444506 426574
rect 444742 426338 462186 426574
rect 462422 426338 462506 426574
rect 462742 426338 480186 426574
rect 480422 426338 480506 426574
rect 480742 426338 498186 426574
rect 498422 426338 498506 426574
rect 498742 426338 516186 426574
rect 516422 426338 516506 426574
rect 516742 426338 534186 426574
rect 534422 426338 534506 426574
rect 534742 426338 546924 426574
rect 547160 426338 547244 426574
rect 547480 426338 548472 426574
rect -4476 426306 548472 426338
rect -4476 423174 548472 423206
rect -4476 422938 -2524 423174
rect -2288 422938 -2204 423174
rect -1968 422938 8466 423174
rect 8702 422938 8786 423174
rect 9022 422938 26466 423174
rect 26702 422938 26786 423174
rect 27022 422938 44466 423174
rect 44702 422938 44786 423174
rect 45022 422938 62466 423174
rect 62702 422938 62786 423174
rect 63022 422938 80466 423174
rect 80702 422938 80786 423174
rect 81022 422938 98466 423174
rect 98702 422938 98786 423174
rect 99022 422938 116466 423174
rect 116702 422938 116786 423174
rect 117022 422938 134466 423174
rect 134702 422938 134786 423174
rect 135022 422938 152466 423174
rect 152702 422938 152786 423174
rect 153022 422938 170466 423174
rect 170702 422938 170786 423174
rect 171022 422938 188466 423174
rect 188702 422938 188786 423174
rect 189022 422938 206466 423174
rect 206702 422938 206786 423174
rect 207022 422938 224466 423174
rect 224702 422938 224786 423174
rect 225022 422938 242466 423174
rect 242702 422938 242786 423174
rect 243022 422938 260466 423174
rect 260702 422938 260786 423174
rect 261022 422938 278466 423174
rect 278702 422938 278786 423174
rect 279022 422938 296466 423174
rect 296702 422938 296786 423174
rect 297022 422938 314466 423174
rect 314702 422938 314786 423174
rect 315022 422938 332466 423174
rect 332702 422938 332786 423174
rect 333022 422938 350466 423174
rect 350702 422938 350786 423174
rect 351022 422938 368466 423174
rect 368702 422938 368786 423174
rect 369022 422938 386466 423174
rect 386702 422938 386786 423174
rect 387022 422938 404466 423174
rect 404702 422938 404786 423174
rect 405022 422938 422466 423174
rect 422702 422938 422786 423174
rect 423022 422938 440466 423174
rect 440702 422938 440786 423174
rect 441022 422938 458466 423174
rect 458702 422938 458786 423174
rect 459022 422938 476466 423174
rect 476702 422938 476786 423174
rect 477022 422938 494466 423174
rect 494702 422938 494786 423174
rect 495022 422938 512466 423174
rect 512702 422938 512786 423174
rect 513022 422938 530466 423174
rect 530702 422938 530786 423174
rect 531022 422938 545964 423174
rect 546200 422938 546284 423174
rect 546520 422938 548472 423174
rect -4476 422854 548472 422938
rect -4476 422618 -2524 422854
rect -2288 422618 -2204 422854
rect -1968 422618 8466 422854
rect 8702 422618 8786 422854
rect 9022 422618 26466 422854
rect 26702 422618 26786 422854
rect 27022 422618 44466 422854
rect 44702 422618 44786 422854
rect 45022 422618 62466 422854
rect 62702 422618 62786 422854
rect 63022 422618 80466 422854
rect 80702 422618 80786 422854
rect 81022 422618 98466 422854
rect 98702 422618 98786 422854
rect 99022 422618 116466 422854
rect 116702 422618 116786 422854
rect 117022 422618 134466 422854
rect 134702 422618 134786 422854
rect 135022 422618 152466 422854
rect 152702 422618 152786 422854
rect 153022 422618 170466 422854
rect 170702 422618 170786 422854
rect 171022 422618 188466 422854
rect 188702 422618 188786 422854
rect 189022 422618 206466 422854
rect 206702 422618 206786 422854
rect 207022 422618 224466 422854
rect 224702 422618 224786 422854
rect 225022 422618 242466 422854
rect 242702 422618 242786 422854
rect 243022 422618 260466 422854
rect 260702 422618 260786 422854
rect 261022 422618 278466 422854
rect 278702 422618 278786 422854
rect 279022 422618 296466 422854
rect 296702 422618 296786 422854
rect 297022 422618 314466 422854
rect 314702 422618 314786 422854
rect 315022 422618 332466 422854
rect 332702 422618 332786 422854
rect 333022 422618 350466 422854
rect 350702 422618 350786 422854
rect 351022 422618 368466 422854
rect 368702 422618 368786 422854
rect 369022 422618 386466 422854
rect 386702 422618 386786 422854
rect 387022 422618 404466 422854
rect 404702 422618 404786 422854
rect 405022 422618 422466 422854
rect 422702 422618 422786 422854
rect 423022 422618 440466 422854
rect 440702 422618 440786 422854
rect 441022 422618 458466 422854
rect 458702 422618 458786 422854
rect 459022 422618 476466 422854
rect 476702 422618 476786 422854
rect 477022 422618 494466 422854
rect 494702 422618 494786 422854
rect 495022 422618 512466 422854
rect 512702 422618 512786 422854
rect 513022 422618 530466 422854
rect 530702 422618 530786 422854
rect 531022 422618 545964 422854
rect 546200 422618 546284 422854
rect 546520 422618 548472 422854
rect -4476 422586 548472 422618
rect -4476 419454 548472 419486
rect -4476 419218 -1564 419454
rect -1328 419218 -1244 419454
rect -1008 419218 4746 419454
rect 4982 419218 5066 419454
rect 5302 419218 22746 419454
rect 22982 419218 23066 419454
rect 23302 419218 40746 419454
rect 40982 419218 41066 419454
rect 41302 419218 58746 419454
rect 58982 419218 59066 419454
rect 59302 419218 76746 419454
rect 76982 419218 77066 419454
rect 77302 419218 94746 419454
rect 94982 419218 95066 419454
rect 95302 419218 112746 419454
rect 112982 419218 113066 419454
rect 113302 419218 130746 419454
rect 130982 419218 131066 419454
rect 131302 419218 148746 419454
rect 148982 419218 149066 419454
rect 149302 419218 166746 419454
rect 166982 419218 167066 419454
rect 167302 419218 184746 419454
rect 184982 419218 185066 419454
rect 185302 419218 202746 419454
rect 202982 419218 203066 419454
rect 203302 419218 220746 419454
rect 220982 419218 221066 419454
rect 221302 419218 238746 419454
rect 238982 419218 239066 419454
rect 239302 419218 256746 419454
rect 256982 419218 257066 419454
rect 257302 419218 274746 419454
rect 274982 419218 275066 419454
rect 275302 419218 292746 419454
rect 292982 419218 293066 419454
rect 293302 419218 310746 419454
rect 310982 419218 311066 419454
rect 311302 419218 328746 419454
rect 328982 419218 329066 419454
rect 329302 419218 346746 419454
rect 346982 419218 347066 419454
rect 347302 419218 364746 419454
rect 364982 419218 365066 419454
rect 365302 419218 382746 419454
rect 382982 419218 383066 419454
rect 383302 419218 400746 419454
rect 400982 419218 401066 419454
rect 401302 419218 418746 419454
rect 418982 419218 419066 419454
rect 419302 419218 436746 419454
rect 436982 419218 437066 419454
rect 437302 419218 454746 419454
rect 454982 419218 455066 419454
rect 455302 419218 472746 419454
rect 472982 419218 473066 419454
rect 473302 419218 490746 419454
rect 490982 419218 491066 419454
rect 491302 419218 508746 419454
rect 508982 419218 509066 419454
rect 509302 419218 526746 419454
rect 526982 419218 527066 419454
rect 527302 419218 545004 419454
rect 545240 419218 545324 419454
rect 545560 419218 548472 419454
rect -4476 419134 548472 419218
rect -4476 418898 -1564 419134
rect -1328 418898 -1244 419134
rect -1008 418898 4746 419134
rect 4982 418898 5066 419134
rect 5302 418898 22746 419134
rect 22982 418898 23066 419134
rect 23302 418898 40746 419134
rect 40982 418898 41066 419134
rect 41302 418898 58746 419134
rect 58982 418898 59066 419134
rect 59302 418898 76746 419134
rect 76982 418898 77066 419134
rect 77302 418898 94746 419134
rect 94982 418898 95066 419134
rect 95302 418898 112746 419134
rect 112982 418898 113066 419134
rect 113302 418898 130746 419134
rect 130982 418898 131066 419134
rect 131302 418898 148746 419134
rect 148982 418898 149066 419134
rect 149302 418898 166746 419134
rect 166982 418898 167066 419134
rect 167302 418898 184746 419134
rect 184982 418898 185066 419134
rect 185302 418898 202746 419134
rect 202982 418898 203066 419134
rect 203302 418898 220746 419134
rect 220982 418898 221066 419134
rect 221302 418898 238746 419134
rect 238982 418898 239066 419134
rect 239302 418898 256746 419134
rect 256982 418898 257066 419134
rect 257302 418898 274746 419134
rect 274982 418898 275066 419134
rect 275302 418898 292746 419134
rect 292982 418898 293066 419134
rect 293302 418898 310746 419134
rect 310982 418898 311066 419134
rect 311302 418898 328746 419134
rect 328982 418898 329066 419134
rect 329302 418898 346746 419134
rect 346982 418898 347066 419134
rect 347302 418898 364746 419134
rect 364982 418898 365066 419134
rect 365302 418898 382746 419134
rect 382982 418898 383066 419134
rect 383302 418898 400746 419134
rect 400982 418898 401066 419134
rect 401302 418898 418746 419134
rect 418982 418898 419066 419134
rect 419302 418898 436746 419134
rect 436982 418898 437066 419134
rect 437302 418898 454746 419134
rect 454982 418898 455066 419134
rect 455302 418898 472746 419134
rect 472982 418898 473066 419134
rect 473302 418898 490746 419134
rect 490982 418898 491066 419134
rect 491302 418898 508746 419134
rect 508982 418898 509066 419134
rect 509302 418898 526746 419134
rect 526982 418898 527066 419134
rect 527302 418898 545004 419134
rect 545240 418898 545324 419134
rect 545560 418898 548472 419134
rect -4476 418866 548472 418898
rect -4476 412614 548472 412646
rect -4476 412378 -4444 412614
rect -4208 412378 -4124 412614
rect -3888 412378 15906 412614
rect 16142 412378 16226 412614
rect 16462 412378 33906 412614
rect 34142 412378 34226 412614
rect 34462 412378 51906 412614
rect 52142 412378 52226 412614
rect 52462 412378 69906 412614
rect 70142 412378 70226 412614
rect 70462 412378 87906 412614
rect 88142 412378 88226 412614
rect 88462 412378 105906 412614
rect 106142 412378 106226 412614
rect 106462 412378 123906 412614
rect 124142 412378 124226 412614
rect 124462 412378 141906 412614
rect 142142 412378 142226 412614
rect 142462 412378 159906 412614
rect 160142 412378 160226 412614
rect 160462 412378 177906 412614
rect 178142 412378 178226 412614
rect 178462 412378 195906 412614
rect 196142 412378 196226 412614
rect 196462 412378 213906 412614
rect 214142 412378 214226 412614
rect 214462 412378 231906 412614
rect 232142 412378 232226 412614
rect 232462 412378 249906 412614
rect 250142 412378 250226 412614
rect 250462 412378 267906 412614
rect 268142 412378 268226 412614
rect 268462 412378 285906 412614
rect 286142 412378 286226 412614
rect 286462 412378 303906 412614
rect 304142 412378 304226 412614
rect 304462 412378 321906 412614
rect 322142 412378 322226 412614
rect 322462 412378 339906 412614
rect 340142 412378 340226 412614
rect 340462 412378 357906 412614
rect 358142 412378 358226 412614
rect 358462 412378 375906 412614
rect 376142 412378 376226 412614
rect 376462 412378 393906 412614
rect 394142 412378 394226 412614
rect 394462 412378 411906 412614
rect 412142 412378 412226 412614
rect 412462 412378 429906 412614
rect 430142 412378 430226 412614
rect 430462 412378 447906 412614
rect 448142 412378 448226 412614
rect 448462 412378 465906 412614
rect 466142 412378 466226 412614
rect 466462 412378 483906 412614
rect 484142 412378 484226 412614
rect 484462 412378 501906 412614
rect 502142 412378 502226 412614
rect 502462 412378 519906 412614
rect 520142 412378 520226 412614
rect 520462 412378 537906 412614
rect 538142 412378 538226 412614
rect 538462 412378 547884 412614
rect 548120 412378 548204 412614
rect 548440 412378 548472 412614
rect -4476 412294 548472 412378
rect -4476 412058 -4444 412294
rect -4208 412058 -4124 412294
rect -3888 412058 15906 412294
rect 16142 412058 16226 412294
rect 16462 412058 33906 412294
rect 34142 412058 34226 412294
rect 34462 412058 51906 412294
rect 52142 412058 52226 412294
rect 52462 412058 69906 412294
rect 70142 412058 70226 412294
rect 70462 412058 87906 412294
rect 88142 412058 88226 412294
rect 88462 412058 105906 412294
rect 106142 412058 106226 412294
rect 106462 412058 123906 412294
rect 124142 412058 124226 412294
rect 124462 412058 141906 412294
rect 142142 412058 142226 412294
rect 142462 412058 159906 412294
rect 160142 412058 160226 412294
rect 160462 412058 177906 412294
rect 178142 412058 178226 412294
rect 178462 412058 195906 412294
rect 196142 412058 196226 412294
rect 196462 412058 213906 412294
rect 214142 412058 214226 412294
rect 214462 412058 231906 412294
rect 232142 412058 232226 412294
rect 232462 412058 249906 412294
rect 250142 412058 250226 412294
rect 250462 412058 267906 412294
rect 268142 412058 268226 412294
rect 268462 412058 285906 412294
rect 286142 412058 286226 412294
rect 286462 412058 303906 412294
rect 304142 412058 304226 412294
rect 304462 412058 321906 412294
rect 322142 412058 322226 412294
rect 322462 412058 339906 412294
rect 340142 412058 340226 412294
rect 340462 412058 357906 412294
rect 358142 412058 358226 412294
rect 358462 412058 375906 412294
rect 376142 412058 376226 412294
rect 376462 412058 393906 412294
rect 394142 412058 394226 412294
rect 394462 412058 411906 412294
rect 412142 412058 412226 412294
rect 412462 412058 429906 412294
rect 430142 412058 430226 412294
rect 430462 412058 447906 412294
rect 448142 412058 448226 412294
rect 448462 412058 465906 412294
rect 466142 412058 466226 412294
rect 466462 412058 483906 412294
rect 484142 412058 484226 412294
rect 484462 412058 501906 412294
rect 502142 412058 502226 412294
rect 502462 412058 519906 412294
rect 520142 412058 520226 412294
rect 520462 412058 537906 412294
rect 538142 412058 538226 412294
rect 538462 412058 547884 412294
rect 548120 412058 548204 412294
rect 548440 412058 548472 412294
rect -4476 412026 548472 412058
rect -4476 408894 548472 408926
rect -4476 408658 -3484 408894
rect -3248 408658 -3164 408894
rect -2928 408658 12186 408894
rect 12422 408658 12506 408894
rect 12742 408658 30186 408894
rect 30422 408658 30506 408894
rect 30742 408658 48186 408894
rect 48422 408658 48506 408894
rect 48742 408658 66186 408894
rect 66422 408658 66506 408894
rect 66742 408658 84186 408894
rect 84422 408658 84506 408894
rect 84742 408658 102186 408894
rect 102422 408658 102506 408894
rect 102742 408658 120186 408894
rect 120422 408658 120506 408894
rect 120742 408658 138186 408894
rect 138422 408658 138506 408894
rect 138742 408658 156186 408894
rect 156422 408658 156506 408894
rect 156742 408658 174186 408894
rect 174422 408658 174506 408894
rect 174742 408658 192186 408894
rect 192422 408658 192506 408894
rect 192742 408658 210186 408894
rect 210422 408658 210506 408894
rect 210742 408658 228186 408894
rect 228422 408658 228506 408894
rect 228742 408658 246186 408894
rect 246422 408658 246506 408894
rect 246742 408658 264186 408894
rect 264422 408658 264506 408894
rect 264742 408658 282186 408894
rect 282422 408658 282506 408894
rect 282742 408658 300186 408894
rect 300422 408658 300506 408894
rect 300742 408658 318186 408894
rect 318422 408658 318506 408894
rect 318742 408658 336186 408894
rect 336422 408658 336506 408894
rect 336742 408658 354186 408894
rect 354422 408658 354506 408894
rect 354742 408658 372186 408894
rect 372422 408658 372506 408894
rect 372742 408658 390186 408894
rect 390422 408658 390506 408894
rect 390742 408658 408186 408894
rect 408422 408658 408506 408894
rect 408742 408658 426186 408894
rect 426422 408658 426506 408894
rect 426742 408658 444186 408894
rect 444422 408658 444506 408894
rect 444742 408658 462186 408894
rect 462422 408658 462506 408894
rect 462742 408658 480186 408894
rect 480422 408658 480506 408894
rect 480742 408658 498186 408894
rect 498422 408658 498506 408894
rect 498742 408658 516186 408894
rect 516422 408658 516506 408894
rect 516742 408658 534186 408894
rect 534422 408658 534506 408894
rect 534742 408658 546924 408894
rect 547160 408658 547244 408894
rect 547480 408658 548472 408894
rect -4476 408574 548472 408658
rect -4476 408338 -3484 408574
rect -3248 408338 -3164 408574
rect -2928 408338 12186 408574
rect 12422 408338 12506 408574
rect 12742 408338 30186 408574
rect 30422 408338 30506 408574
rect 30742 408338 48186 408574
rect 48422 408338 48506 408574
rect 48742 408338 66186 408574
rect 66422 408338 66506 408574
rect 66742 408338 84186 408574
rect 84422 408338 84506 408574
rect 84742 408338 102186 408574
rect 102422 408338 102506 408574
rect 102742 408338 120186 408574
rect 120422 408338 120506 408574
rect 120742 408338 138186 408574
rect 138422 408338 138506 408574
rect 138742 408338 156186 408574
rect 156422 408338 156506 408574
rect 156742 408338 174186 408574
rect 174422 408338 174506 408574
rect 174742 408338 192186 408574
rect 192422 408338 192506 408574
rect 192742 408338 210186 408574
rect 210422 408338 210506 408574
rect 210742 408338 228186 408574
rect 228422 408338 228506 408574
rect 228742 408338 246186 408574
rect 246422 408338 246506 408574
rect 246742 408338 264186 408574
rect 264422 408338 264506 408574
rect 264742 408338 282186 408574
rect 282422 408338 282506 408574
rect 282742 408338 300186 408574
rect 300422 408338 300506 408574
rect 300742 408338 318186 408574
rect 318422 408338 318506 408574
rect 318742 408338 336186 408574
rect 336422 408338 336506 408574
rect 336742 408338 354186 408574
rect 354422 408338 354506 408574
rect 354742 408338 372186 408574
rect 372422 408338 372506 408574
rect 372742 408338 390186 408574
rect 390422 408338 390506 408574
rect 390742 408338 408186 408574
rect 408422 408338 408506 408574
rect 408742 408338 426186 408574
rect 426422 408338 426506 408574
rect 426742 408338 444186 408574
rect 444422 408338 444506 408574
rect 444742 408338 462186 408574
rect 462422 408338 462506 408574
rect 462742 408338 480186 408574
rect 480422 408338 480506 408574
rect 480742 408338 498186 408574
rect 498422 408338 498506 408574
rect 498742 408338 516186 408574
rect 516422 408338 516506 408574
rect 516742 408338 534186 408574
rect 534422 408338 534506 408574
rect 534742 408338 546924 408574
rect 547160 408338 547244 408574
rect 547480 408338 548472 408574
rect -4476 408306 548472 408338
rect -4476 405174 548472 405206
rect -4476 404938 -2524 405174
rect -2288 404938 -2204 405174
rect -1968 404938 8466 405174
rect 8702 404938 8786 405174
rect 9022 404938 26466 405174
rect 26702 404938 26786 405174
rect 27022 404938 44466 405174
rect 44702 404938 44786 405174
rect 45022 404938 62466 405174
rect 62702 404938 62786 405174
rect 63022 404938 80466 405174
rect 80702 404938 80786 405174
rect 81022 404938 98466 405174
rect 98702 404938 98786 405174
rect 99022 404938 116466 405174
rect 116702 404938 116786 405174
rect 117022 404938 134466 405174
rect 134702 404938 134786 405174
rect 135022 404938 152466 405174
rect 152702 404938 152786 405174
rect 153022 404938 170466 405174
rect 170702 404938 170786 405174
rect 171022 404938 188466 405174
rect 188702 404938 188786 405174
rect 189022 404938 206466 405174
rect 206702 404938 206786 405174
rect 207022 404938 224466 405174
rect 224702 404938 224786 405174
rect 225022 404938 242466 405174
rect 242702 404938 242786 405174
rect 243022 404938 260466 405174
rect 260702 404938 260786 405174
rect 261022 404938 278466 405174
rect 278702 404938 278786 405174
rect 279022 404938 296466 405174
rect 296702 404938 296786 405174
rect 297022 404938 314466 405174
rect 314702 404938 314786 405174
rect 315022 404938 332466 405174
rect 332702 404938 332786 405174
rect 333022 404938 350466 405174
rect 350702 404938 350786 405174
rect 351022 404938 368466 405174
rect 368702 404938 368786 405174
rect 369022 404938 386466 405174
rect 386702 404938 386786 405174
rect 387022 404938 404466 405174
rect 404702 404938 404786 405174
rect 405022 404938 422466 405174
rect 422702 404938 422786 405174
rect 423022 404938 440466 405174
rect 440702 404938 440786 405174
rect 441022 404938 458466 405174
rect 458702 404938 458786 405174
rect 459022 404938 476466 405174
rect 476702 404938 476786 405174
rect 477022 404938 494466 405174
rect 494702 404938 494786 405174
rect 495022 404938 512466 405174
rect 512702 404938 512786 405174
rect 513022 404938 530466 405174
rect 530702 404938 530786 405174
rect 531022 404938 545964 405174
rect 546200 404938 546284 405174
rect 546520 404938 548472 405174
rect -4476 404854 548472 404938
rect -4476 404618 -2524 404854
rect -2288 404618 -2204 404854
rect -1968 404618 8466 404854
rect 8702 404618 8786 404854
rect 9022 404618 26466 404854
rect 26702 404618 26786 404854
rect 27022 404618 44466 404854
rect 44702 404618 44786 404854
rect 45022 404618 62466 404854
rect 62702 404618 62786 404854
rect 63022 404618 80466 404854
rect 80702 404618 80786 404854
rect 81022 404618 98466 404854
rect 98702 404618 98786 404854
rect 99022 404618 116466 404854
rect 116702 404618 116786 404854
rect 117022 404618 134466 404854
rect 134702 404618 134786 404854
rect 135022 404618 152466 404854
rect 152702 404618 152786 404854
rect 153022 404618 170466 404854
rect 170702 404618 170786 404854
rect 171022 404618 188466 404854
rect 188702 404618 188786 404854
rect 189022 404618 206466 404854
rect 206702 404618 206786 404854
rect 207022 404618 224466 404854
rect 224702 404618 224786 404854
rect 225022 404618 242466 404854
rect 242702 404618 242786 404854
rect 243022 404618 260466 404854
rect 260702 404618 260786 404854
rect 261022 404618 278466 404854
rect 278702 404618 278786 404854
rect 279022 404618 296466 404854
rect 296702 404618 296786 404854
rect 297022 404618 314466 404854
rect 314702 404618 314786 404854
rect 315022 404618 332466 404854
rect 332702 404618 332786 404854
rect 333022 404618 350466 404854
rect 350702 404618 350786 404854
rect 351022 404618 368466 404854
rect 368702 404618 368786 404854
rect 369022 404618 386466 404854
rect 386702 404618 386786 404854
rect 387022 404618 404466 404854
rect 404702 404618 404786 404854
rect 405022 404618 422466 404854
rect 422702 404618 422786 404854
rect 423022 404618 440466 404854
rect 440702 404618 440786 404854
rect 441022 404618 458466 404854
rect 458702 404618 458786 404854
rect 459022 404618 476466 404854
rect 476702 404618 476786 404854
rect 477022 404618 494466 404854
rect 494702 404618 494786 404854
rect 495022 404618 512466 404854
rect 512702 404618 512786 404854
rect 513022 404618 530466 404854
rect 530702 404618 530786 404854
rect 531022 404618 545964 404854
rect 546200 404618 546284 404854
rect 546520 404618 548472 404854
rect -4476 404586 548472 404618
rect -4476 401454 548472 401486
rect -4476 401218 -1564 401454
rect -1328 401218 -1244 401454
rect -1008 401218 4746 401454
rect 4982 401218 5066 401454
rect 5302 401218 22746 401454
rect 22982 401218 23066 401454
rect 23302 401218 40746 401454
rect 40982 401218 41066 401454
rect 41302 401218 58746 401454
rect 58982 401218 59066 401454
rect 59302 401218 76746 401454
rect 76982 401218 77066 401454
rect 77302 401218 94746 401454
rect 94982 401218 95066 401454
rect 95302 401218 112746 401454
rect 112982 401218 113066 401454
rect 113302 401218 130746 401454
rect 130982 401218 131066 401454
rect 131302 401218 148746 401454
rect 148982 401218 149066 401454
rect 149302 401218 166746 401454
rect 166982 401218 167066 401454
rect 167302 401218 184746 401454
rect 184982 401218 185066 401454
rect 185302 401218 202746 401454
rect 202982 401218 203066 401454
rect 203302 401218 220746 401454
rect 220982 401218 221066 401454
rect 221302 401218 238746 401454
rect 238982 401218 239066 401454
rect 239302 401218 256746 401454
rect 256982 401218 257066 401454
rect 257302 401218 274746 401454
rect 274982 401218 275066 401454
rect 275302 401218 292746 401454
rect 292982 401218 293066 401454
rect 293302 401218 310746 401454
rect 310982 401218 311066 401454
rect 311302 401218 328746 401454
rect 328982 401218 329066 401454
rect 329302 401218 346746 401454
rect 346982 401218 347066 401454
rect 347302 401218 364746 401454
rect 364982 401218 365066 401454
rect 365302 401218 382746 401454
rect 382982 401218 383066 401454
rect 383302 401218 400746 401454
rect 400982 401218 401066 401454
rect 401302 401218 418746 401454
rect 418982 401218 419066 401454
rect 419302 401218 436746 401454
rect 436982 401218 437066 401454
rect 437302 401218 454746 401454
rect 454982 401218 455066 401454
rect 455302 401218 472746 401454
rect 472982 401218 473066 401454
rect 473302 401218 490746 401454
rect 490982 401218 491066 401454
rect 491302 401218 508746 401454
rect 508982 401218 509066 401454
rect 509302 401218 526746 401454
rect 526982 401218 527066 401454
rect 527302 401218 545004 401454
rect 545240 401218 545324 401454
rect 545560 401218 548472 401454
rect -4476 401134 548472 401218
rect -4476 400898 -1564 401134
rect -1328 400898 -1244 401134
rect -1008 400898 4746 401134
rect 4982 400898 5066 401134
rect 5302 400898 22746 401134
rect 22982 400898 23066 401134
rect 23302 400898 40746 401134
rect 40982 400898 41066 401134
rect 41302 400898 58746 401134
rect 58982 400898 59066 401134
rect 59302 400898 76746 401134
rect 76982 400898 77066 401134
rect 77302 400898 94746 401134
rect 94982 400898 95066 401134
rect 95302 400898 112746 401134
rect 112982 400898 113066 401134
rect 113302 400898 130746 401134
rect 130982 400898 131066 401134
rect 131302 400898 148746 401134
rect 148982 400898 149066 401134
rect 149302 400898 166746 401134
rect 166982 400898 167066 401134
rect 167302 400898 184746 401134
rect 184982 400898 185066 401134
rect 185302 400898 202746 401134
rect 202982 400898 203066 401134
rect 203302 400898 220746 401134
rect 220982 400898 221066 401134
rect 221302 400898 238746 401134
rect 238982 400898 239066 401134
rect 239302 400898 256746 401134
rect 256982 400898 257066 401134
rect 257302 400898 274746 401134
rect 274982 400898 275066 401134
rect 275302 400898 292746 401134
rect 292982 400898 293066 401134
rect 293302 400898 310746 401134
rect 310982 400898 311066 401134
rect 311302 400898 328746 401134
rect 328982 400898 329066 401134
rect 329302 400898 346746 401134
rect 346982 400898 347066 401134
rect 347302 400898 364746 401134
rect 364982 400898 365066 401134
rect 365302 400898 382746 401134
rect 382982 400898 383066 401134
rect 383302 400898 400746 401134
rect 400982 400898 401066 401134
rect 401302 400898 418746 401134
rect 418982 400898 419066 401134
rect 419302 400898 436746 401134
rect 436982 400898 437066 401134
rect 437302 400898 454746 401134
rect 454982 400898 455066 401134
rect 455302 400898 472746 401134
rect 472982 400898 473066 401134
rect 473302 400898 490746 401134
rect 490982 400898 491066 401134
rect 491302 400898 508746 401134
rect 508982 400898 509066 401134
rect 509302 400898 526746 401134
rect 526982 400898 527066 401134
rect 527302 400898 545004 401134
rect 545240 400898 545324 401134
rect 545560 400898 548472 401134
rect -4476 400866 548472 400898
rect -4476 394614 548472 394646
rect -4476 394378 -4444 394614
rect -4208 394378 -4124 394614
rect -3888 394378 15906 394614
rect 16142 394378 16226 394614
rect 16462 394378 33906 394614
rect 34142 394378 34226 394614
rect 34462 394378 51906 394614
rect 52142 394378 52226 394614
rect 52462 394378 69906 394614
rect 70142 394378 70226 394614
rect 70462 394378 87906 394614
rect 88142 394378 88226 394614
rect 88462 394378 105906 394614
rect 106142 394378 106226 394614
rect 106462 394378 123906 394614
rect 124142 394378 124226 394614
rect 124462 394378 141906 394614
rect 142142 394378 142226 394614
rect 142462 394378 159906 394614
rect 160142 394378 160226 394614
rect 160462 394378 177906 394614
rect 178142 394378 178226 394614
rect 178462 394378 195906 394614
rect 196142 394378 196226 394614
rect 196462 394378 213906 394614
rect 214142 394378 214226 394614
rect 214462 394378 231906 394614
rect 232142 394378 232226 394614
rect 232462 394378 249906 394614
rect 250142 394378 250226 394614
rect 250462 394378 267906 394614
rect 268142 394378 268226 394614
rect 268462 394378 285906 394614
rect 286142 394378 286226 394614
rect 286462 394378 303906 394614
rect 304142 394378 304226 394614
rect 304462 394378 321906 394614
rect 322142 394378 322226 394614
rect 322462 394378 339906 394614
rect 340142 394378 340226 394614
rect 340462 394378 357906 394614
rect 358142 394378 358226 394614
rect 358462 394378 375906 394614
rect 376142 394378 376226 394614
rect 376462 394378 393906 394614
rect 394142 394378 394226 394614
rect 394462 394378 411906 394614
rect 412142 394378 412226 394614
rect 412462 394378 429906 394614
rect 430142 394378 430226 394614
rect 430462 394378 447906 394614
rect 448142 394378 448226 394614
rect 448462 394378 465906 394614
rect 466142 394378 466226 394614
rect 466462 394378 483906 394614
rect 484142 394378 484226 394614
rect 484462 394378 501906 394614
rect 502142 394378 502226 394614
rect 502462 394378 519906 394614
rect 520142 394378 520226 394614
rect 520462 394378 537906 394614
rect 538142 394378 538226 394614
rect 538462 394378 547884 394614
rect 548120 394378 548204 394614
rect 548440 394378 548472 394614
rect -4476 394294 548472 394378
rect -4476 394058 -4444 394294
rect -4208 394058 -4124 394294
rect -3888 394058 15906 394294
rect 16142 394058 16226 394294
rect 16462 394058 33906 394294
rect 34142 394058 34226 394294
rect 34462 394058 51906 394294
rect 52142 394058 52226 394294
rect 52462 394058 69906 394294
rect 70142 394058 70226 394294
rect 70462 394058 87906 394294
rect 88142 394058 88226 394294
rect 88462 394058 105906 394294
rect 106142 394058 106226 394294
rect 106462 394058 123906 394294
rect 124142 394058 124226 394294
rect 124462 394058 141906 394294
rect 142142 394058 142226 394294
rect 142462 394058 159906 394294
rect 160142 394058 160226 394294
rect 160462 394058 177906 394294
rect 178142 394058 178226 394294
rect 178462 394058 195906 394294
rect 196142 394058 196226 394294
rect 196462 394058 213906 394294
rect 214142 394058 214226 394294
rect 214462 394058 231906 394294
rect 232142 394058 232226 394294
rect 232462 394058 249906 394294
rect 250142 394058 250226 394294
rect 250462 394058 267906 394294
rect 268142 394058 268226 394294
rect 268462 394058 285906 394294
rect 286142 394058 286226 394294
rect 286462 394058 303906 394294
rect 304142 394058 304226 394294
rect 304462 394058 321906 394294
rect 322142 394058 322226 394294
rect 322462 394058 339906 394294
rect 340142 394058 340226 394294
rect 340462 394058 357906 394294
rect 358142 394058 358226 394294
rect 358462 394058 375906 394294
rect 376142 394058 376226 394294
rect 376462 394058 393906 394294
rect 394142 394058 394226 394294
rect 394462 394058 411906 394294
rect 412142 394058 412226 394294
rect 412462 394058 429906 394294
rect 430142 394058 430226 394294
rect 430462 394058 447906 394294
rect 448142 394058 448226 394294
rect 448462 394058 465906 394294
rect 466142 394058 466226 394294
rect 466462 394058 483906 394294
rect 484142 394058 484226 394294
rect 484462 394058 501906 394294
rect 502142 394058 502226 394294
rect 502462 394058 519906 394294
rect 520142 394058 520226 394294
rect 520462 394058 537906 394294
rect 538142 394058 538226 394294
rect 538462 394058 547884 394294
rect 548120 394058 548204 394294
rect 548440 394058 548472 394294
rect -4476 394026 548472 394058
rect -4476 390894 548472 390926
rect -4476 390658 -3484 390894
rect -3248 390658 -3164 390894
rect -2928 390658 12186 390894
rect 12422 390658 12506 390894
rect 12742 390658 30186 390894
rect 30422 390658 30506 390894
rect 30742 390658 48186 390894
rect 48422 390658 48506 390894
rect 48742 390658 66186 390894
rect 66422 390658 66506 390894
rect 66742 390658 84186 390894
rect 84422 390658 84506 390894
rect 84742 390658 102186 390894
rect 102422 390658 102506 390894
rect 102742 390658 120186 390894
rect 120422 390658 120506 390894
rect 120742 390658 138186 390894
rect 138422 390658 138506 390894
rect 138742 390658 156186 390894
rect 156422 390658 156506 390894
rect 156742 390658 174186 390894
rect 174422 390658 174506 390894
rect 174742 390658 192186 390894
rect 192422 390658 192506 390894
rect 192742 390658 210186 390894
rect 210422 390658 210506 390894
rect 210742 390658 228186 390894
rect 228422 390658 228506 390894
rect 228742 390658 246186 390894
rect 246422 390658 246506 390894
rect 246742 390658 264186 390894
rect 264422 390658 264506 390894
rect 264742 390658 282186 390894
rect 282422 390658 282506 390894
rect 282742 390658 300186 390894
rect 300422 390658 300506 390894
rect 300742 390658 318186 390894
rect 318422 390658 318506 390894
rect 318742 390658 336186 390894
rect 336422 390658 336506 390894
rect 336742 390658 354186 390894
rect 354422 390658 354506 390894
rect 354742 390658 372186 390894
rect 372422 390658 372506 390894
rect 372742 390658 390186 390894
rect 390422 390658 390506 390894
rect 390742 390658 408186 390894
rect 408422 390658 408506 390894
rect 408742 390658 426186 390894
rect 426422 390658 426506 390894
rect 426742 390658 444186 390894
rect 444422 390658 444506 390894
rect 444742 390658 462186 390894
rect 462422 390658 462506 390894
rect 462742 390658 480186 390894
rect 480422 390658 480506 390894
rect 480742 390658 498186 390894
rect 498422 390658 498506 390894
rect 498742 390658 516186 390894
rect 516422 390658 516506 390894
rect 516742 390658 534186 390894
rect 534422 390658 534506 390894
rect 534742 390658 546924 390894
rect 547160 390658 547244 390894
rect 547480 390658 548472 390894
rect -4476 390574 548472 390658
rect -4476 390338 -3484 390574
rect -3248 390338 -3164 390574
rect -2928 390338 12186 390574
rect 12422 390338 12506 390574
rect 12742 390338 30186 390574
rect 30422 390338 30506 390574
rect 30742 390338 48186 390574
rect 48422 390338 48506 390574
rect 48742 390338 66186 390574
rect 66422 390338 66506 390574
rect 66742 390338 84186 390574
rect 84422 390338 84506 390574
rect 84742 390338 102186 390574
rect 102422 390338 102506 390574
rect 102742 390338 120186 390574
rect 120422 390338 120506 390574
rect 120742 390338 138186 390574
rect 138422 390338 138506 390574
rect 138742 390338 156186 390574
rect 156422 390338 156506 390574
rect 156742 390338 174186 390574
rect 174422 390338 174506 390574
rect 174742 390338 192186 390574
rect 192422 390338 192506 390574
rect 192742 390338 210186 390574
rect 210422 390338 210506 390574
rect 210742 390338 228186 390574
rect 228422 390338 228506 390574
rect 228742 390338 246186 390574
rect 246422 390338 246506 390574
rect 246742 390338 264186 390574
rect 264422 390338 264506 390574
rect 264742 390338 282186 390574
rect 282422 390338 282506 390574
rect 282742 390338 300186 390574
rect 300422 390338 300506 390574
rect 300742 390338 318186 390574
rect 318422 390338 318506 390574
rect 318742 390338 336186 390574
rect 336422 390338 336506 390574
rect 336742 390338 354186 390574
rect 354422 390338 354506 390574
rect 354742 390338 372186 390574
rect 372422 390338 372506 390574
rect 372742 390338 390186 390574
rect 390422 390338 390506 390574
rect 390742 390338 408186 390574
rect 408422 390338 408506 390574
rect 408742 390338 426186 390574
rect 426422 390338 426506 390574
rect 426742 390338 444186 390574
rect 444422 390338 444506 390574
rect 444742 390338 462186 390574
rect 462422 390338 462506 390574
rect 462742 390338 480186 390574
rect 480422 390338 480506 390574
rect 480742 390338 498186 390574
rect 498422 390338 498506 390574
rect 498742 390338 516186 390574
rect 516422 390338 516506 390574
rect 516742 390338 534186 390574
rect 534422 390338 534506 390574
rect 534742 390338 546924 390574
rect 547160 390338 547244 390574
rect 547480 390338 548472 390574
rect -4476 390306 548472 390338
rect -4476 387174 548472 387206
rect -4476 386938 -2524 387174
rect -2288 386938 -2204 387174
rect -1968 386938 8466 387174
rect 8702 386938 8786 387174
rect 9022 386938 26466 387174
rect 26702 386938 26786 387174
rect 27022 386938 44466 387174
rect 44702 386938 44786 387174
rect 45022 386938 62466 387174
rect 62702 386938 62786 387174
rect 63022 386938 80466 387174
rect 80702 386938 80786 387174
rect 81022 386938 98466 387174
rect 98702 386938 98786 387174
rect 99022 386938 116466 387174
rect 116702 386938 116786 387174
rect 117022 386938 134466 387174
rect 134702 386938 134786 387174
rect 135022 386938 152466 387174
rect 152702 386938 152786 387174
rect 153022 386938 170466 387174
rect 170702 386938 170786 387174
rect 171022 386938 188466 387174
rect 188702 386938 188786 387174
rect 189022 386938 206466 387174
rect 206702 386938 206786 387174
rect 207022 386938 224466 387174
rect 224702 386938 224786 387174
rect 225022 386938 242466 387174
rect 242702 386938 242786 387174
rect 243022 386938 260466 387174
rect 260702 386938 260786 387174
rect 261022 386938 278466 387174
rect 278702 386938 278786 387174
rect 279022 386938 296466 387174
rect 296702 386938 296786 387174
rect 297022 386938 314466 387174
rect 314702 386938 314786 387174
rect 315022 386938 332466 387174
rect 332702 386938 332786 387174
rect 333022 386938 350466 387174
rect 350702 386938 350786 387174
rect 351022 386938 368466 387174
rect 368702 386938 368786 387174
rect 369022 386938 386466 387174
rect 386702 386938 386786 387174
rect 387022 386938 404466 387174
rect 404702 386938 404786 387174
rect 405022 386938 422466 387174
rect 422702 386938 422786 387174
rect 423022 386938 440466 387174
rect 440702 386938 440786 387174
rect 441022 386938 458466 387174
rect 458702 386938 458786 387174
rect 459022 386938 476466 387174
rect 476702 386938 476786 387174
rect 477022 386938 494466 387174
rect 494702 386938 494786 387174
rect 495022 386938 512466 387174
rect 512702 386938 512786 387174
rect 513022 386938 530466 387174
rect 530702 386938 530786 387174
rect 531022 386938 545964 387174
rect 546200 386938 546284 387174
rect 546520 386938 548472 387174
rect -4476 386854 548472 386938
rect -4476 386618 -2524 386854
rect -2288 386618 -2204 386854
rect -1968 386618 8466 386854
rect 8702 386618 8786 386854
rect 9022 386618 26466 386854
rect 26702 386618 26786 386854
rect 27022 386618 44466 386854
rect 44702 386618 44786 386854
rect 45022 386618 62466 386854
rect 62702 386618 62786 386854
rect 63022 386618 80466 386854
rect 80702 386618 80786 386854
rect 81022 386618 98466 386854
rect 98702 386618 98786 386854
rect 99022 386618 116466 386854
rect 116702 386618 116786 386854
rect 117022 386618 134466 386854
rect 134702 386618 134786 386854
rect 135022 386618 152466 386854
rect 152702 386618 152786 386854
rect 153022 386618 170466 386854
rect 170702 386618 170786 386854
rect 171022 386618 188466 386854
rect 188702 386618 188786 386854
rect 189022 386618 206466 386854
rect 206702 386618 206786 386854
rect 207022 386618 224466 386854
rect 224702 386618 224786 386854
rect 225022 386618 242466 386854
rect 242702 386618 242786 386854
rect 243022 386618 260466 386854
rect 260702 386618 260786 386854
rect 261022 386618 278466 386854
rect 278702 386618 278786 386854
rect 279022 386618 296466 386854
rect 296702 386618 296786 386854
rect 297022 386618 314466 386854
rect 314702 386618 314786 386854
rect 315022 386618 332466 386854
rect 332702 386618 332786 386854
rect 333022 386618 350466 386854
rect 350702 386618 350786 386854
rect 351022 386618 368466 386854
rect 368702 386618 368786 386854
rect 369022 386618 386466 386854
rect 386702 386618 386786 386854
rect 387022 386618 404466 386854
rect 404702 386618 404786 386854
rect 405022 386618 422466 386854
rect 422702 386618 422786 386854
rect 423022 386618 440466 386854
rect 440702 386618 440786 386854
rect 441022 386618 458466 386854
rect 458702 386618 458786 386854
rect 459022 386618 476466 386854
rect 476702 386618 476786 386854
rect 477022 386618 494466 386854
rect 494702 386618 494786 386854
rect 495022 386618 512466 386854
rect 512702 386618 512786 386854
rect 513022 386618 530466 386854
rect 530702 386618 530786 386854
rect 531022 386618 545964 386854
rect 546200 386618 546284 386854
rect 546520 386618 548472 386854
rect -4476 386586 548472 386618
rect -4476 383454 548472 383486
rect -4476 383218 -1564 383454
rect -1328 383218 -1244 383454
rect -1008 383218 4746 383454
rect 4982 383218 5066 383454
rect 5302 383218 22746 383454
rect 22982 383218 23066 383454
rect 23302 383218 40746 383454
rect 40982 383218 41066 383454
rect 41302 383218 58746 383454
rect 58982 383218 59066 383454
rect 59302 383218 76746 383454
rect 76982 383218 77066 383454
rect 77302 383218 94746 383454
rect 94982 383218 95066 383454
rect 95302 383218 112746 383454
rect 112982 383218 113066 383454
rect 113302 383218 130746 383454
rect 130982 383218 131066 383454
rect 131302 383218 148746 383454
rect 148982 383218 149066 383454
rect 149302 383218 166746 383454
rect 166982 383218 167066 383454
rect 167302 383218 184746 383454
rect 184982 383218 185066 383454
rect 185302 383218 202746 383454
rect 202982 383218 203066 383454
rect 203302 383218 220746 383454
rect 220982 383218 221066 383454
rect 221302 383218 238746 383454
rect 238982 383218 239066 383454
rect 239302 383218 256746 383454
rect 256982 383218 257066 383454
rect 257302 383218 274746 383454
rect 274982 383218 275066 383454
rect 275302 383218 292746 383454
rect 292982 383218 293066 383454
rect 293302 383218 310746 383454
rect 310982 383218 311066 383454
rect 311302 383218 328746 383454
rect 328982 383218 329066 383454
rect 329302 383218 346746 383454
rect 346982 383218 347066 383454
rect 347302 383218 364746 383454
rect 364982 383218 365066 383454
rect 365302 383218 382746 383454
rect 382982 383218 383066 383454
rect 383302 383218 400746 383454
rect 400982 383218 401066 383454
rect 401302 383218 418746 383454
rect 418982 383218 419066 383454
rect 419302 383218 436746 383454
rect 436982 383218 437066 383454
rect 437302 383218 454746 383454
rect 454982 383218 455066 383454
rect 455302 383218 472746 383454
rect 472982 383218 473066 383454
rect 473302 383218 490746 383454
rect 490982 383218 491066 383454
rect 491302 383218 508746 383454
rect 508982 383218 509066 383454
rect 509302 383218 526746 383454
rect 526982 383218 527066 383454
rect 527302 383218 545004 383454
rect 545240 383218 545324 383454
rect 545560 383218 548472 383454
rect -4476 383134 548472 383218
rect -4476 382898 -1564 383134
rect -1328 382898 -1244 383134
rect -1008 382898 4746 383134
rect 4982 382898 5066 383134
rect 5302 382898 22746 383134
rect 22982 382898 23066 383134
rect 23302 382898 40746 383134
rect 40982 382898 41066 383134
rect 41302 382898 58746 383134
rect 58982 382898 59066 383134
rect 59302 382898 76746 383134
rect 76982 382898 77066 383134
rect 77302 382898 94746 383134
rect 94982 382898 95066 383134
rect 95302 382898 112746 383134
rect 112982 382898 113066 383134
rect 113302 382898 130746 383134
rect 130982 382898 131066 383134
rect 131302 382898 148746 383134
rect 148982 382898 149066 383134
rect 149302 382898 166746 383134
rect 166982 382898 167066 383134
rect 167302 382898 184746 383134
rect 184982 382898 185066 383134
rect 185302 382898 202746 383134
rect 202982 382898 203066 383134
rect 203302 382898 220746 383134
rect 220982 382898 221066 383134
rect 221302 382898 238746 383134
rect 238982 382898 239066 383134
rect 239302 382898 256746 383134
rect 256982 382898 257066 383134
rect 257302 382898 274746 383134
rect 274982 382898 275066 383134
rect 275302 382898 292746 383134
rect 292982 382898 293066 383134
rect 293302 382898 310746 383134
rect 310982 382898 311066 383134
rect 311302 382898 328746 383134
rect 328982 382898 329066 383134
rect 329302 382898 346746 383134
rect 346982 382898 347066 383134
rect 347302 382898 364746 383134
rect 364982 382898 365066 383134
rect 365302 382898 382746 383134
rect 382982 382898 383066 383134
rect 383302 382898 400746 383134
rect 400982 382898 401066 383134
rect 401302 382898 418746 383134
rect 418982 382898 419066 383134
rect 419302 382898 436746 383134
rect 436982 382898 437066 383134
rect 437302 382898 454746 383134
rect 454982 382898 455066 383134
rect 455302 382898 472746 383134
rect 472982 382898 473066 383134
rect 473302 382898 490746 383134
rect 490982 382898 491066 383134
rect 491302 382898 508746 383134
rect 508982 382898 509066 383134
rect 509302 382898 526746 383134
rect 526982 382898 527066 383134
rect 527302 382898 545004 383134
rect 545240 382898 545324 383134
rect 545560 382898 548472 383134
rect -4476 382866 548472 382898
rect -4476 376614 548472 376646
rect -4476 376378 -4444 376614
rect -4208 376378 -4124 376614
rect -3888 376378 15906 376614
rect 16142 376378 16226 376614
rect 16462 376378 33906 376614
rect 34142 376378 34226 376614
rect 34462 376378 51906 376614
rect 52142 376378 52226 376614
rect 52462 376378 69906 376614
rect 70142 376378 70226 376614
rect 70462 376378 87906 376614
rect 88142 376378 88226 376614
rect 88462 376378 105906 376614
rect 106142 376378 106226 376614
rect 106462 376378 123906 376614
rect 124142 376378 124226 376614
rect 124462 376378 141906 376614
rect 142142 376378 142226 376614
rect 142462 376378 159906 376614
rect 160142 376378 160226 376614
rect 160462 376378 177906 376614
rect 178142 376378 178226 376614
rect 178462 376378 195906 376614
rect 196142 376378 196226 376614
rect 196462 376378 213906 376614
rect 214142 376378 214226 376614
rect 214462 376378 231906 376614
rect 232142 376378 232226 376614
rect 232462 376378 249906 376614
rect 250142 376378 250226 376614
rect 250462 376378 267906 376614
rect 268142 376378 268226 376614
rect 268462 376378 285906 376614
rect 286142 376378 286226 376614
rect 286462 376378 303906 376614
rect 304142 376378 304226 376614
rect 304462 376378 321906 376614
rect 322142 376378 322226 376614
rect 322462 376378 339906 376614
rect 340142 376378 340226 376614
rect 340462 376378 357906 376614
rect 358142 376378 358226 376614
rect 358462 376378 375906 376614
rect 376142 376378 376226 376614
rect 376462 376378 393906 376614
rect 394142 376378 394226 376614
rect 394462 376378 411906 376614
rect 412142 376378 412226 376614
rect 412462 376378 429906 376614
rect 430142 376378 430226 376614
rect 430462 376378 447906 376614
rect 448142 376378 448226 376614
rect 448462 376378 465906 376614
rect 466142 376378 466226 376614
rect 466462 376378 483906 376614
rect 484142 376378 484226 376614
rect 484462 376378 501906 376614
rect 502142 376378 502226 376614
rect 502462 376378 519906 376614
rect 520142 376378 520226 376614
rect 520462 376378 537906 376614
rect 538142 376378 538226 376614
rect 538462 376378 547884 376614
rect 548120 376378 548204 376614
rect 548440 376378 548472 376614
rect -4476 376294 548472 376378
rect -4476 376058 -4444 376294
rect -4208 376058 -4124 376294
rect -3888 376058 15906 376294
rect 16142 376058 16226 376294
rect 16462 376058 33906 376294
rect 34142 376058 34226 376294
rect 34462 376058 51906 376294
rect 52142 376058 52226 376294
rect 52462 376058 69906 376294
rect 70142 376058 70226 376294
rect 70462 376058 87906 376294
rect 88142 376058 88226 376294
rect 88462 376058 105906 376294
rect 106142 376058 106226 376294
rect 106462 376058 123906 376294
rect 124142 376058 124226 376294
rect 124462 376058 141906 376294
rect 142142 376058 142226 376294
rect 142462 376058 159906 376294
rect 160142 376058 160226 376294
rect 160462 376058 177906 376294
rect 178142 376058 178226 376294
rect 178462 376058 195906 376294
rect 196142 376058 196226 376294
rect 196462 376058 213906 376294
rect 214142 376058 214226 376294
rect 214462 376058 231906 376294
rect 232142 376058 232226 376294
rect 232462 376058 249906 376294
rect 250142 376058 250226 376294
rect 250462 376058 267906 376294
rect 268142 376058 268226 376294
rect 268462 376058 285906 376294
rect 286142 376058 286226 376294
rect 286462 376058 303906 376294
rect 304142 376058 304226 376294
rect 304462 376058 321906 376294
rect 322142 376058 322226 376294
rect 322462 376058 339906 376294
rect 340142 376058 340226 376294
rect 340462 376058 357906 376294
rect 358142 376058 358226 376294
rect 358462 376058 375906 376294
rect 376142 376058 376226 376294
rect 376462 376058 393906 376294
rect 394142 376058 394226 376294
rect 394462 376058 411906 376294
rect 412142 376058 412226 376294
rect 412462 376058 429906 376294
rect 430142 376058 430226 376294
rect 430462 376058 447906 376294
rect 448142 376058 448226 376294
rect 448462 376058 465906 376294
rect 466142 376058 466226 376294
rect 466462 376058 483906 376294
rect 484142 376058 484226 376294
rect 484462 376058 501906 376294
rect 502142 376058 502226 376294
rect 502462 376058 519906 376294
rect 520142 376058 520226 376294
rect 520462 376058 537906 376294
rect 538142 376058 538226 376294
rect 538462 376058 547884 376294
rect 548120 376058 548204 376294
rect 548440 376058 548472 376294
rect -4476 376026 548472 376058
rect -4476 372894 548472 372926
rect -4476 372658 -3484 372894
rect -3248 372658 -3164 372894
rect -2928 372658 12186 372894
rect 12422 372658 12506 372894
rect 12742 372658 30186 372894
rect 30422 372658 30506 372894
rect 30742 372658 48186 372894
rect 48422 372658 48506 372894
rect 48742 372658 66186 372894
rect 66422 372658 66506 372894
rect 66742 372658 84186 372894
rect 84422 372658 84506 372894
rect 84742 372658 102186 372894
rect 102422 372658 102506 372894
rect 102742 372658 120186 372894
rect 120422 372658 120506 372894
rect 120742 372658 138186 372894
rect 138422 372658 138506 372894
rect 138742 372658 156186 372894
rect 156422 372658 156506 372894
rect 156742 372658 174186 372894
rect 174422 372658 174506 372894
rect 174742 372658 192186 372894
rect 192422 372658 192506 372894
rect 192742 372658 210186 372894
rect 210422 372658 210506 372894
rect 210742 372658 228186 372894
rect 228422 372658 228506 372894
rect 228742 372658 246186 372894
rect 246422 372658 246506 372894
rect 246742 372658 264186 372894
rect 264422 372658 264506 372894
rect 264742 372658 282186 372894
rect 282422 372658 282506 372894
rect 282742 372658 300186 372894
rect 300422 372658 300506 372894
rect 300742 372658 318186 372894
rect 318422 372658 318506 372894
rect 318742 372658 336186 372894
rect 336422 372658 336506 372894
rect 336742 372658 354186 372894
rect 354422 372658 354506 372894
rect 354742 372658 372186 372894
rect 372422 372658 372506 372894
rect 372742 372658 390186 372894
rect 390422 372658 390506 372894
rect 390742 372658 408186 372894
rect 408422 372658 408506 372894
rect 408742 372658 426186 372894
rect 426422 372658 426506 372894
rect 426742 372658 444186 372894
rect 444422 372658 444506 372894
rect 444742 372658 462186 372894
rect 462422 372658 462506 372894
rect 462742 372658 480186 372894
rect 480422 372658 480506 372894
rect 480742 372658 498186 372894
rect 498422 372658 498506 372894
rect 498742 372658 516186 372894
rect 516422 372658 516506 372894
rect 516742 372658 534186 372894
rect 534422 372658 534506 372894
rect 534742 372658 546924 372894
rect 547160 372658 547244 372894
rect 547480 372658 548472 372894
rect -4476 372574 548472 372658
rect -4476 372338 -3484 372574
rect -3248 372338 -3164 372574
rect -2928 372338 12186 372574
rect 12422 372338 12506 372574
rect 12742 372338 30186 372574
rect 30422 372338 30506 372574
rect 30742 372338 48186 372574
rect 48422 372338 48506 372574
rect 48742 372338 66186 372574
rect 66422 372338 66506 372574
rect 66742 372338 84186 372574
rect 84422 372338 84506 372574
rect 84742 372338 102186 372574
rect 102422 372338 102506 372574
rect 102742 372338 120186 372574
rect 120422 372338 120506 372574
rect 120742 372338 138186 372574
rect 138422 372338 138506 372574
rect 138742 372338 156186 372574
rect 156422 372338 156506 372574
rect 156742 372338 174186 372574
rect 174422 372338 174506 372574
rect 174742 372338 192186 372574
rect 192422 372338 192506 372574
rect 192742 372338 210186 372574
rect 210422 372338 210506 372574
rect 210742 372338 228186 372574
rect 228422 372338 228506 372574
rect 228742 372338 246186 372574
rect 246422 372338 246506 372574
rect 246742 372338 264186 372574
rect 264422 372338 264506 372574
rect 264742 372338 282186 372574
rect 282422 372338 282506 372574
rect 282742 372338 300186 372574
rect 300422 372338 300506 372574
rect 300742 372338 318186 372574
rect 318422 372338 318506 372574
rect 318742 372338 336186 372574
rect 336422 372338 336506 372574
rect 336742 372338 354186 372574
rect 354422 372338 354506 372574
rect 354742 372338 372186 372574
rect 372422 372338 372506 372574
rect 372742 372338 390186 372574
rect 390422 372338 390506 372574
rect 390742 372338 408186 372574
rect 408422 372338 408506 372574
rect 408742 372338 426186 372574
rect 426422 372338 426506 372574
rect 426742 372338 444186 372574
rect 444422 372338 444506 372574
rect 444742 372338 462186 372574
rect 462422 372338 462506 372574
rect 462742 372338 480186 372574
rect 480422 372338 480506 372574
rect 480742 372338 498186 372574
rect 498422 372338 498506 372574
rect 498742 372338 516186 372574
rect 516422 372338 516506 372574
rect 516742 372338 534186 372574
rect 534422 372338 534506 372574
rect 534742 372338 546924 372574
rect 547160 372338 547244 372574
rect 547480 372338 548472 372574
rect -4476 372306 548472 372338
rect -4476 369174 548472 369206
rect -4476 368938 -2524 369174
rect -2288 368938 -2204 369174
rect -1968 368938 8466 369174
rect 8702 368938 8786 369174
rect 9022 368938 26466 369174
rect 26702 368938 26786 369174
rect 27022 368938 44466 369174
rect 44702 368938 44786 369174
rect 45022 368938 62466 369174
rect 62702 368938 62786 369174
rect 63022 368938 80466 369174
rect 80702 368938 80786 369174
rect 81022 368938 98466 369174
rect 98702 368938 98786 369174
rect 99022 368938 116466 369174
rect 116702 368938 116786 369174
rect 117022 368938 134466 369174
rect 134702 368938 134786 369174
rect 135022 368938 152466 369174
rect 152702 368938 152786 369174
rect 153022 368938 170466 369174
rect 170702 368938 170786 369174
rect 171022 368938 188466 369174
rect 188702 368938 188786 369174
rect 189022 368938 206466 369174
rect 206702 368938 206786 369174
rect 207022 368938 224466 369174
rect 224702 368938 224786 369174
rect 225022 368938 242466 369174
rect 242702 368938 242786 369174
rect 243022 368938 260466 369174
rect 260702 368938 260786 369174
rect 261022 368938 278466 369174
rect 278702 368938 278786 369174
rect 279022 368938 296466 369174
rect 296702 368938 296786 369174
rect 297022 368938 314466 369174
rect 314702 368938 314786 369174
rect 315022 368938 332466 369174
rect 332702 368938 332786 369174
rect 333022 368938 350466 369174
rect 350702 368938 350786 369174
rect 351022 368938 368466 369174
rect 368702 368938 368786 369174
rect 369022 368938 386466 369174
rect 386702 368938 386786 369174
rect 387022 368938 404466 369174
rect 404702 368938 404786 369174
rect 405022 368938 422466 369174
rect 422702 368938 422786 369174
rect 423022 368938 440466 369174
rect 440702 368938 440786 369174
rect 441022 368938 458466 369174
rect 458702 368938 458786 369174
rect 459022 368938 476466 369174
rect 476702 368938 476786 369174
rect 477022 368938 494466 369174
rect 494702 368938 494786 369174
rect 495022 368938 512466 369174
rect 512702 368938 512786 369174
rect 513022 368938 530466 369174
rect 530702 368938 530786 369174
rect 531022 368938 545964 369174
rect 546200 368938 546284 369174
rect 546520 368938 548472 369174
rect -4476 368854 548472 368938
rect -4476 368618 -2524 368854
rect -2288 368618 -2204 368854
rect -1968 368618 8466 368854
rect 8702 368618 8786 368854
rect 9022 368618 26466 368854
rect 26702 368618 26786 368854
rect 27022 368618 44466 368854
rect 44702 368618 44786 368854
rect 45022 368618 62466 368854
rect 62702 368618 62786 368854
rect 63022 368618 80466 368854
rect 80702 368618 80786 368854
rect 81022 368618 98466 368854
rect 98702 368618 98786 368854
rect 99022 368618 116466 368854
rect 116702 368618 116786 368854
rect 117022 368618 134466 368854
rect 134702 368618 134786 368854
rect 135022 368618 152466 368854
rect 152702 368618 152786 368854
rect 153022 368618 170466 368854
rect 170702 368618 170786 368854
rect 171022 368618 188466 368854
rect 188702 368618 188786 368854
rect 189022 368618 206466 368854
rect 206702 368618 206786 368854
rect 207022 368618 224466 368854
rect 224702 368618 224786 368854
rect 225022 368618 242466 368854
rect 242702 368618 242786 368854
rect 243022 368618 260466 368854
rect 260702 368618 260786 368854
rect 261022 368618 278466 368854
rect 278702 368618 278786 368854
rect 279022 368618 296466 368854
rect 296702 368618 296786 368854
rect 297022 368618 314466 368854
rect 314702 368618 314786 368854
rect 315022 368618 332466 368854
rect 332702 368618 332786 368854
rect 333022 368618 350466 368854
rect 350702 368618 350786 368854
rect 351022 368618 368466 368854
rect 368702 368618 368786 368854
rect 369022 368618 386466 368854
rect 386702 368618 386786 368854
rect 387022 368618 404466 368854
rect 404702 368618 404786 368854
rect 405022 368618 422466 368854
rect 422702 368618 422786 368854
rect 423022 368618 440466 368854
rect 440702 368618 440786 368854
rect 441022 368618 458466 368854
rect 458702 368618 458786 368854
rect 459022 368618 476466 368854
rect 476702 368618 476786 368854
rect 477022 368618 494466 368854
rect 494702 368618 494786 368854
rect 495022 368618 512466 368854
rect 512702 368618 512786 368854
rect 513022 368618 530466 368854
rect 530702 368618 530786 368854
rect 531022 368618 545964 368854
rect 546200 368618 546284 368854
rect 546520 368618 548472 368854
rect -4476 368586 548472 368618
rect -4476 365454 548472 365486
rect -4476 365218 -1564 365454
rect -1328 365218 -1244 365454
rect -1008 365218 4746 365454
rect 4982 365218 5066 365454
rect 5302 365218 22746 365454
rect 22982 365218 23066 365454
rect 23302 365218 40746 365454
rect 40982 365218 41066 365454
rect 41302 365218 58746 365454
rect 58982 365218 59066 365454
rect 59302 365218 76746 365454
rect 76982 365218 77066 365454
rect 77302 365218 94746 365454
rect 94982 365218 95066 365454
rect 95302 365218 112746 365454
rect 112982 365218 113066 365454
rect 113302 365218 130746 365454
rect 130982 365218 131066 365454
rect 131302 365218 148746 365454
rect 148982 365218 149066 365454
rect 149302 365218 166746 365454
rect 166982 365218 167066 365454
rect 167302 365218 184746 365454
rect 184982 365218 185066 365454
rect 185302 365218 202746 365454
rect 202982 365218 203066 365454
rect 203302 365218 220746 365454
rect 220982 365218 221066 365454
rect 221302 365218 238746 365454
rect 238982 365218 239066 365454
rect 239302 365218 256746 365454
rect 256982 365218 257066 365454
rect 257302 365218 274746 365454
rect 274982 365218 275066 365454
rect 275302 365218 292746 365454
rect 292982 365218 293066 365454
rect 293302 365218 310746 365454
rect 310982 365218 311066 365454
rect 311302 365218 328746 365454
rect 328982 365218 329066 365454
rect 329302 365218 346746 365454
rect 346982 365218 347066 365454
rect 347302 365218 364746 365454
rect 364982 365218 365066 365454
rect 365302 365218 382746 365454
rect 382982 365218 383066 365454
rect 383302 365218 400746 365454
rect 400982 365218 401066 365454
rect 401302 365218 418746 365454
rect 418982 365218 419066 365454
rect 419302 365218 436746 365454
rect 436982 365218 437066 365454
rect 437302 365218 454746 365454
rect 454982 365218 455066 365454
rect 455302 365218 472746 365454
rect 472982 365218 473066 365454
rect 473302 365218 490746 365454
rect 490982 365218 491066 365454
rect 491302 365218 508746 365454
rect 508982 365218 509066 365454
rect 509302 365218 526746 365454
rect 526982 365218 527066 365454
rect 527302 365218 545004 365454
rect 545240 365218 545324 365454
rect 545560 365218 548472 365454
rect -4476 365134 548472 365218
rect -4476 364898 -1564 365134
rect -1328 364898 -1244 365134
rect -1008 364898 4746 365134
rect 4982 364898 5066 365134
rect 5302 364898 22746 365134
rect 22982 364898 23066 365134
rect 23302 364898 40746 365134
rect 40982 364898 41066 365134
rect 41302 364898 58746 365134
rect 58982 364898 59066 365134
rect 59302 364898 76746 365134
rect 76982 364898 77066 365134
rect 77302 364898 94746 365134
rect 94982 364898 95066 365134
rect 95302 364898 112746 365134
rect 112982 364898 113066 365134
rect 113302 364898 130746 365134
rect 130982 364898 131066 365134
rect 131302 364898 148746 365134
rect 148982 364898 149066 365134
rect 149302 364898 166746 365134
rect 166982 364898 167066 365134
rect 167302 364898 184746 365134
rect 184982 364898 185066 365134
rect 185302 364898 202746 365134
rect 202982 364898 203066 365134
rect 203302 364898 220746 365134
rect 220982 364898 221066 365134
rect 221302 364898 238746 365134
rect 238982 364898 239066 365134
rect 239302 364898 256746 365134
rect 256982 364898 257066 365134
rect 257302 364898 274746 365134
rect 274982 364898 275066 365134
rect 275302 364898 292746 365134
rect 292982 364898 293066 365134
rect 293302 364898 310746 365134
rect 310982 364898 311066 365134
rect 311302 364898 328746 365134
rect 328982 364898 329066 365134
rect 329302 364898 346746 365134
rect 346982 364898 347066 365134
rect 347302 364898 364746 365134
rect 364982 364898 365066 365134
rect 365302 364898 382746 365134
rect 382982 364898 383066 365134
rect 383302 364898 400746 365134
rect 400982 364898 401066 365134
rect 401302 364898 418746 365134
rect 418982 364898 419066 365134
rect 419302 364898 436746 365134
rect 436982 364898 437066 365134
rect 437302 364898 454746 365134
rect 454982 364898 455066 365134
rect 455302 364898 472746 365134
rect 472982 364898 473066 365134
rect 473302 364898 490746 365134
rect 490982 364898 491066 365134
rect 491302 364898 508746 365134
rect 508982 364898 509066 365134
rect 509302 364898 526746 365134
rect 526982 364898 527066 365134
rect 527302 364898 545004 365134
rect 545240 364898 545324 365134
rect 545560 364898 548472 365134
rect -4476 364866 548472 364898
rect -4476 358614 548472 358646
rect -4476 358378 -4444 358614
rect -4208 358378 -4124 358614
rect -3888 358378 15906 358614
rect 16142 358378 16226 358614
rect 16462 358378 33906 358614
rect 34142 358378 34226 358614
rect 34462 358378 51906 358614
rect 52142 358378 52226 358614
rect 52462 358378 69906 358614
rect 70142 358378 70226 358614
rect 70462 358378 87906 358614
rect 88142 358378 88226 358614
rect 88462 358378 105906 358614
rect 106142 358378 106226 358614
rect 106462 358378 123906 358614
rect 124142 358378 124226 358614
rect 124462 358378 141906 358614
rect 142142 358378 142226 358614
rect 142462 358378 159906 358614
rect 160142 358378 160226 358614
rect 160462 358378 177906 358614
rect 178142 358378 178226 358614
rect 178462 358378 195906 358614
rect 196142 358378 196226 358614
rect 196462 358378 213906 358614
rect 214142 358378 214226 358614
rect 214462 358378 231906 358614
rect 232142 358378 232226 358614
rect 232462 358378 249906 358614
rect 250142 358378 250226 358614
rect 250462 358378 267906 358614
rect 268142 358378 268226 358614
rect 268462 358378 285906 358614
rect 286142 358378 286226 358614
rect 286462 358378 303906 358614
rect 304142 358378 304226 358614
rect 304462 358378 321906 358614
rect 322142 358378 322226 358614
rect 322462 358378 339906 358614
rect 340142 358378 340226 358614
rect 340462 358378 357906 358614
rect 358142 358378 358226 358614
rect 358462 358378 375906 358614
rect 376142 358378 376226 358614
rect 376462 358378 393906 358614
rect 394142 358378 394226 358614
rect 394462 358378 411906 358614
rect 412142 358378 412226 358614
rect 412462 358378 429906 358614
rect 430142 358378 430226 358614
rect 430462 358378 447906 358614
rect 448142 358378 448226 358614
rect 448462 358378 465906 358614
rect 466142 358378 466226 358614
rect 466462 358378 483906 358614
rect 484142 358378 484226 358614
rect 484462 358378 501906 358614
rect 502142 358378 502226 358614
rect 502462 358378 519906 358614
rect 520142 358378 520226 358614
rect 520462 358378 537906 358614
rect 538142 358378 538226 358614
rect 538462 358378 547884 358614
rect 548120 358378 548204 358614
rect 548440 358378 548472 358614
rect -4476 358294 548472 358378
rect -4476 358058 -4444 358294
rect -4208 358058 -4124 358294
rect -3888 358058 15906 358294
rect 16142 358058 16226 358294
rect 16462 358058 33906 358294
rect 34142 358058 34226 358294
rect 34462 358058 51906 358294
rect 52142 358058 52226 358294
rect 52462 358058 69906 358294
rect 70142 358058 70226 358294
rect 70462 358058 87906 358294
rect 88142 358058 88226 358294
rect 88462 358058 105906 358294
rect 106142 358058 106226 358294
rect 106462 358058 123906 358294
rect 124142 358058 124226 358294
rect 124462 358058 141906 358294
rect 142142 358058 142226 358294
rect 142462 358058 159906 358294
rect 160142 358058 160226 358294
rect 160462 358058 177906 358294
rect 178142 358058 178226 358294
rect 178462 358058 195906 358294
rect 196142 358058 196226 358294
rect 196462 358058 213906 358294
rect 214142 358058 214226 358294
rect 214462 358058 231906 358294
rect 232142 358058 232226 358294
rect 232462 358058 249906 358294
rect 250142 358058 250226 358294
rect 250462 358058 267906 358294
rect 268142 358058 268226 358294
rect 268462 358058 285906 358294
rect 286142 358058 286226 358294
rect 286462 358058 303906 358294
rect 304142 358058 304226 358294
rect 304462 358058 321906 358294
rect 322142 358058 322226 358294
rect 322462 358058 339906 358294
rect 340142 358058 340226 358294
rect 340462 358058 357906 358294
rect 358142 358058 358226 358294
rect 358462 358058 375906 358294
rect 376142 358058 376226 358294
rect 376462 358058 393906 358294
rect 394142 358058 394226 358294
rect 394462 358058 411906 358294
rect 412142 358058 412226 358294
rect 412462 358058 429906 358294
rect 430142 358058 430226 358294
rect 430462 358058 447906 358294
rect 448142 358058 448226 358294
rect 448462 358058 465906 358294
rect 466142 358058 466226 358294
rect 466462 358058 483906 358294
rect 484142 358058 484226 358294
rect 484462 358058 501906 358294
rect 502142 358058 502226 358294
rect 502462 358058 519906 358294
rect 520142 358058 520226 358294
rect 520462 358058 537906 358294
rect 538142 358058 538226 358294
rect 538462 358058 547884 358294
rect 548120 358058 548204 358294
rect 548440 358058 548472 358294
rect -4476 358026 548472 358058
rect -4476 354894 548472 354926
rect -4476 354658 -3484 354894
rect -3248 354658 -3164 354894
rect -2928 354658 12186 354894
rect 12422 354658 12506 354894
rect 12742 354658 30186 354894
rect 30422 354658 30506 354894
rect 30742 354658 48186 354894
rect 48422 354658 48506 354894
rect 48742 354658 66186 354894
rect 66422 354658 66506 354894
rect 66742 354658 84186 354894
rect 84422 354658 84506 354894
rect 84742 354658 102186 354894
rect 102422 354658 102506 354894
rect 102742 354658 120186 354894
rect 120422 354658 120506 354894
rect 120742 354658 138186 354894
rect 138422 354658 138506 354894
rect 138742 354658 156186 354894
rect 156422 354658 156506 354894
rect 156742 354658 174186 354894
rect 174422 354658 174506 354894
rect 174742 354658 192186 354894
rect 192422 354658 192506 354894
rect 192742 354658 210186 354894
rect 210422 354658 210506 354894
rect 210742 354658 228186 354894
rect 228422 354658 228506 354894
rect 228742 354658 246186 354894
rect 246422 354658 246506 354894
rect 246742 354658 264186 354894
rect 264422 354658 264506 354894
rect 264742 354658 282186 354894
rect 282422 354658 282506 354894
rect 282742 354658 300186 354894
rect 300422 354658 300506 354894
rect 300742 354658 318186 354894
rect 318422 354658 318506 354894
rect 318742 354658 336186 354894
rect 336422 354658 336506 354894
rect 336742 354658 354186 354894
rect 354422 354658 354506 354894
rect 354742 354658 372186 354894
rect 372422 354658 372506 354894
rect 372742 354658 390186 354894
rect 390422 354658 390506 354894
rect 390742 354658 408186 354894
rect 408422 354658 408506 354894
rect 408742 354658 426186 354894
rect 426422 354658 426506 354894
rect 426742 354658 444186 354894
rect 444422 354658 444506 354894
rect 444742 354658 462186 354894
rect 462422 354658 462506 354894
rect 462742 354658 480186 354894
rect 480422 354658 480506 354894
rect 480742 354658 498186 354894
rect 498422 354658 498506 354894
rect 498742 354658 516186 354894
rect 516422 354658 516506 354894
rect 516742 354658 534186 354894
rect 534422 354658 534506 354894
rect 534742 354658 546924 354894
rect 547160 354658 547244 354894
rect 547480 354658 548472 354894
rect -4476 354574 548472 354658
rect -4476 354338 -3484 354574
rect -3248 354338 -3164 354574
rect -2928 354338 12186 354574
rect 12422 354338 12506 354574
rect 12742 354338 30186 354574
rect 30422 354338 30506 354574
rect 30742 354338 48186 354574
rect 48422 354338 48506 354574
rect 48742 354338 66186 354574
rect 66422 354338 66506 354574
rect 66742 354338 84186 354574
rect 84422 354338 84506 354574
rect 84742 354338 102186 354574
rect 102422 354338 102506 354574
rect 102742 354338 120186 354574
rect 120422 354338 120506 354574
rect 120742 354338 138186 354574
rect 138422 354338 138506 354574
rect 138742 354338 156186 354574
rect 156422 354338 156506 354574
rect 156742 354338 174186 354574
rect 174422 354338 174506 354574
rect 174742 354338 192186 354574
rect 192422 354338 192506 354574
rect 192742 354338 210186 354574
rect 210422 354338 210506 354574
rect 210742 354338 228186 354574
rect 228422 354338 228506 354574
rect 228742 354338 246186 354574
rect 246422 354338 246506 354574
rect 246742 354338 264186 354574
rect 264422 354338 264506 354574
rect 264742 354338 282186 354574
rect 282422 354338 282506 354574
rect 282742 354338 300186 354574
rect 300422 354338 300506 354574
rect 300742 354338 318186 354574
rect 318422 354338 318506 354574
rect 318742 354338 336186 354574
rect 336422 354338 336506 354574
rect 336742 354338 354186 354574
rect 354422 354338 354506 354574
rect 354742 354338 372186 354574
rect 372422 354338 372506 354574
rect 372742 354338 390186 354574
rect 390422 354338 390506 354574
rect 390742 354338 408186 354574
rect 408422 354338 408506 354574
rect 408742 354338 426186 354574
rect 426422 354338 426506 354574
rect 426742 354338 444186 354574
rect 444422 354338 444506 354574
rect 444742 354338 462186 354574
rect 462422 354338 462506 354574
rect 462742 354338 480186 354574
rect 480422 354338 480506 354574
rect 480742 354338 498186 354574
rect 498422 354338 498506 354574
rect 498742 354338 516186 354574
rect 516422 354338 516506 354574
rect 516742 354338 534186 354574
rect 534422 354338 534506 354574
rect 534742 354338 546924 354574
rect 547160 354338 547244 354574
rect 547480 354338 548472 354574
rect -4476 354306 548472 354338
rect -4476 351174 548472 351206
rect -4476 350938 -2524 351174
rect -2288 350938 -2204 351174
rect -1968 350938 8466 351174
rect 8702 350938 8786 351174
rect 9022 350938 26466 351174
rect 26702 350938 26786 351174
rect 27022 350938 44466 351174
rect 44702 350938 44786 351174
rect 45022 350938 62466 351174
rect 62702 350938 62786 351174
rect 63022 350938 80466 351174
rect 80702 350938 80786 351174
rect 81022 350938 98466 351174
rect 98702 350938 98786 351174
rect 99022 350938 116466 351174
rect 116702 350938 116786 351174
rect 117022 350938 134466 351174
rect 134702 350938 134786 351174
rect 135022 350938 152466 351174
rect 152702 350938 152786 351174
rect 153022 350938 170466 351174
rect 170702 350938 170786 351174
rect 171022 350938 188466 351174
rect 188702 350938 188786 351174
rect 189022 350938 206466 351174
rect 206702 350938 206786 351174
rect 207022 350938 224466 351174
rect 224702 350938 224786 351174
rect 225022 350938 242466 351174
rect 242702 350938 242786 351174
rect 243022 350938 260466 351174
rect 260702 350938 260786 351174
rect 261022 350938 278466 351174
rect 278702 350938 278786 351174
rect 279022 350938 296466 351174
rect 296702 350938 296786 351174
rect 297022 350938 314466 351174
rect 314702 350938 314786 351174
rect 315022 350938 332466 351174
rect 332702 350938 332786 351174
rect 333022 350938 350466 351174
rect 350702 350938 350786 351174
rect 351022 350938 368466 351174
rect 368702 350938 368786 351174
rect 369022 350938 386466 351174
rect 386702 350938 386786 351174
rect 387022 350938 404466 351174
rect 404702 350938 404786 351174
rect 405022 350938 422466 351174
rect 422702 350938 422786 351174
rect 423022 350938 440466 351174
rect 440702 350938 440786 351174
rect 441022 350938 458466 351174
rect 458702 350938 458786 351174
rect 459022 350938 476466 351174
rect 476702 350938 476786 351174
rect 477022 350938 494466 351174
rect 494702 350938 494786 351174
rect 495022 350938 512466 351174
rect 512702 350938 512786 351174
rect 513022 350938 530466 351174
rect 530702 350938 530786 351174
rect 531022 350938 545964 351174
rect 546200 350938 546284 351174
rect 546520 350938 548472 351174
rect -4476 350854 548472 350938
rect -4476 350618 -2524 350854
rect -2288 350618 -2204 350854
rect -1968 350618 8466 350854
rect 8702 350618 8786 350854
rect 9022 350618 26466 350854
rect 26702 350618 26786 350854
rect 27022 350618 44466 350854
rect 44702 350618 44786 350854
rect 45022 350618 62466 350854
rect 62702 350618 62786 350854
rect 63022 350618 80466 350854
rect 80702 350618 80786 350854
rect 81022 350618 98466 350854
rect 98702 350618 98786 350854
rect 99022 350618 116466 350854
rect 116702 350618 116786 350854
rect 117022 350618 134466 350854
rect 134702 350618 134786 350854
rect 135022 350618 152466 350854
rect 152702 350618 152786 350854
rect 153022 350618 170466 350854
rect 170702 350618 170786 350854
rect 171022 350618 188466 350854
rect 188702 350618 188786 350854
rect 189022 350618 206466 350854
rect 206702 350618 206786 350854
rect 207022 350618 224466 350854
rect 224702 350618 224786 350854
rect 225022 350618 242466 350854
rect 242702 350618 242786 350854
rect 243022 350618 260466 350854
rect 260702 350618 260786 350854
rect 261022 350618 278466 350854
rect 278702 350618 278786 350854
rect 279022 350618 296466 350854
rect 296702 350618 296786 350854
rect 297022 350618 314466 350854
rect 314702 350618 314786 350854
rect 315022 350618 332466 350854
rect 332702 350618 332786 350854
rect 333022 350618 350466 350854
rect 350702 350618 350786 350854
rect 351022 350618 368466 350854
rect 368702 350618 368786 350854
rect 369022 350618 386466 350854
rect 386702 350618 386786 350854
rect 387022 350618 404466 350854
rect 404702 350618 404786 350854
rect 405022 350618 422466 350854
rect 422702 350618 422786 350854
rect 423022 350618 440466 350854
rect 440702 350618 440786 350854
rect 441022 350618 458466 350854
rect 458702 350618 458786 350854
rect 459022 350618 476466 350854
rect 476702 350618 476786 350854
rect 477022 350618 494466 350854
rect 494702 350618 494786 350854
rect 495022 350618 512466 350854
rect 512702 350618 512786 350854
rect 513022 350618 530466 350854
rect 530702 350618 530786 350854
rect 531022 350618 545964 350854
rect 546200 350618 546284 350854
rect 546520 350618 548472 350854
rect -4476 350586 548472 350618
rect -4476 347454 548472 347486
rect -4476 347218 -1564 347454
rect -1328 347218 -1244 347454
rect -1008 347218 4746 347454
rect 4982 347218 5066 347454
rect 5302 347218 22746 347454
rect 22982 347218 23066 347454
rect 23302 347218 40746 347454
rect 40982 347218 41066 347454
rect 41302 347218 58746 347454
rect 58982 347218 59066 347454
rect 59302 347218 76746 347454
rect 76982 347218 77066 347454
rect 77302 347218 94746 347454
rect 94982 347218 95066 347454
rect 95302 347218 112746 347454
rect 112982 347218 113066 347454
rect 113302 347218 130746 347454
rect 130982 347218 131066 347454
rect 131302 347218 148746 347454
rect 148982 347218 149066 347454
rect 149302 347218 166746 347454
rect 166982 347218 167066 347454
rect 167302 347218 184746 347454
rect 184982 347218 185066 347454
rect 185302 347218 202746 347454
rect 202982 347218 203066 347454
rect 203302 347218 220746 347454
rect 220982 347218 221066 347454
rect 221302 347218 238746 347454
rect 238982 347218 239066 347454
rect 239302 347218 256746 347454
rect 256982 347218 257066 347454
rect 257302 347218 274746 347454
rect 274982 347218 275066 347454
rect 275302 347218 292746 347454
rect 292982 347218 293066 347454
rect 293302 347218 310746 347454
rect 310982 347218 311066 347454
rect 311302 347218 328746 347454
rect 328982 347218 329066 347454
rect 329302 347218 346746 347454
rect 346982 347218 347066 347454
rect 347302 347218 364746 347454
rect 364982 347218 365066 347454
rect 365302 347218 382746 347454
rect 382982 347218 383066 347454
rect 383302 347218 400746 347454
rect 400982 347218 401066 347454
rect 401302 347218 418746 347454
rect 418982 347218 419066 347454
rect 419302 347218 436746 347454
rect 436982 347218 437066 347454
rect 437302 347218 454746 347454
rect 454982 347218 455066 347454
rect 455302 347218 472746 347454
rect 472982 347218 473066 347454
rect 473302 347218 490746 347454
rect 490982 347218 491066 347454
rect 491302 347218 508746 347454
rect 508982 347218 509066 347454
rect 509302 347218 526746 347454
rect 526982 347218 527066 347454
rect 527302 347218 545004 347454
rect 545240 347218 545324 347454
rect 545560 347218 548472 347454
rect -4476 347134 548472 347218
rect -4476 346898 -1564 347134
rect -1328 346898 -1244 347134
rect -1008 346898 4746 347134
rect 4982 346898 5066 347134
rect 5302 346898 22746 347134
rect 22982 346898 23066 347134
rect 23302 346898 40746 347134
rect 40982 346898 41066 347134
rect 41302 346898 58746 347134
rect 58982 346898 59066 347134
rect 59302 346898 76746 347134
rect 76982 346898 77066 347134
rect 77302 346898 94746 347134
rect 94982 346898 95066 347134
rect 95302 346898 112746 347134
rect 112982 346898 113066 347134
rect 113302 346898 130746 347134
rect 130982 346898 131066 347134
rect 131302 346898 148746 347134
rect 148982 346898 149066 347134
rect 149302 346898 166746 347134
rect 166982 346898 167066 347134
rect 167302 346898 184746 347134
rect 184982 346898 185066 347134
rect 185302 346898 202746 347134
rect 202982 346898 203066 347134
rect 203302 346898 220746 347134
rect 220982 346898 221066 347134
rect 221302 346898 238746 347134
rect 238982 346898 239066 347134
rect 239302 346898 256746 347134
rect 256982 346898 257066 347134
rect 257302 346898 274746 347134
rect 274982 346898 275066 347134
rect 275302 346898 292746 347134
rect 292982 346898 293066 347134
rect 293302 346898 310746 347134
rect 310982 346898 311066 347134
rect 311302 346898 328746 347134
rect 328982 346898 329066 347134
rect 329302 346898 346746 347134
rect 346982 346898 347066 347134
rect 347302 346898 364746 347134
rect 364982 346898 365066 347134
rect 365302 346898 382746 347134
rect 382982 346898 383066 347134
rect 383302 346898 400746 347134
rect 400982 346898 401066 347134
rect 401302 346898 418746 347134
rect 418982 346898 419066 347134
rect 419302 346898 436746 347134
rect 436982 346898 437066 347134
rect 437302 346898 454746 347134
rect 454982 346898 455066 347134
rect 455302 346898 472746 347134
rect 472982 346898 473066 347134
rect 473302 346898 490746 347134
rect 490982 346898 491066 347134
rect 491302 346898 508746 347134
rect 508982 346898 509066 347134
rect 509302 346898 526746 347134
rect 526982 346898 527066 347134
rect 527302 346898 545004 347134
rect 545240 346898 545324 347134
rect 545560 346898 548472 347134
rect -4476 346866 548472 346898
rect -4476 340614 548472 340646
rect -4476 340378 -4444 340614
rect -4208 340378 -4124 340614
rect -3888 340378 15906 340614
rect 16142 340378 16226 340614
rect 16462 340378 33906 340614
rect 34142 340378 34226 340614
rect 34462 340378 51906 340614
rect 52142 340378 52226 340614
rect 52462 340378 69906 340614
rect 70142 340378 70226 340614
rect 70462 340378 87906 340614
rect 88142 340378 88226 340614
rect 88462 340378 105906 340614
rect 106142 340378 106226 340614
rect 106462 340378 123906 340614
rect 124142 340378 124226 340614
rect 124462 340378 141906 340614
rect 142142 340378 142226 340614
rect 142462 340378 159906 340614
rect 160142 340378 160226 340614
rect 160462 340378 177906 340614
rect 178142 340378 178226 340614
rect 178462 340378 195906 340614
rect 196142 340378 196226 340614
rect 196462 340378 213906 340614
rect 214142 340378 214226 340614
rect 214462 340378 231906 340614
rect 232142 340378 232226 340614
rect 232462 340378 249906 340614
rect 250142 340378 250226 340614
rect 250462 340378 267906 340614
rect 268142 340378 268226 340614
rect 268462 340378 285906 340614
rect 286142 340378 286226 340614
rect 286462 340378 303906 340614
rect 304142 340378 304226 340614
rect 304462 340378 321906 340614
rect 322142 340378 322226 340614
rect 322462 340378 339906 340614
rect 340142 340378 340226 340614
rect 340462 340378 357906 340614
rect 358142 340378 358226 340614
rect 358462 340378 375906 340614
rect 376142 340378 376226 340614
rect 376462 340378 393906 340614
rect 394142 340378 394226 340614
rect 394462 340378 411906 340614
rect 412142 340378 412226 340614
rect 412462 340378 429906 340614
rect 430142 340378 430226 340614
rect 430462 340378 447906 340614
rect 448142 340378 448226 340614
rect 448462 340378 465906 340614
rect 466142 340378 466226 340614
rect 466462 340378 483906 340614
rect 484142 340378 484226 340614
rect 484462 340378 501906 340614
rect 502142 340378 502226 340614
rect 502462 340378 519906 340614
rect 520142 340378 520226 340614
rect 520462 340378 537906 340614
rect 538142 340378 538226 340614
rect 538462 340378 547884 340614
rect 548120 340378 548204 340614
rect 548440 340378 548472 340614
rect -4476 340294 548472 340378
rect -4476 340058 -4444 340294
rect -4208 340058 -4124 340294
rect -3888 340058 15906 340294
rect 16142 340058 16226 340294
rect 16462 340058 33906 340294
rect 34142 340058 34226 340294
rect 34462 340058 51906 340294
rect 52142 340058 52226 340294
rect 52462 340058 69906 340294
rect 70142 340058 70226 340294
rect 70462 340058 87906 340294
rect 88142 340058 88226 340294
rect 88462 340058 105906 340294
rect 106142 340058 106226 340294
rect 106462 340058 123906 340294
rect 124142 340058 124226 340294
rect 124462 340058 141906 340294
rect 142142 340058 142226 340294
rect 142462 340058 159906 340294
rect 160142 340058 160226 340294
rect 160462 340058 177906 340294
rect 178142 340058 178226 340294
rect 178462 340058 195906 340294
rect 196142 340058 196226 340294
rect 196462 340058 213906 340294
rect 214142 340058 214226 340294
rect 214462 340058 231906 340294
rect 232142 340058 232226 340294
rect 232462 340058 249906 340294
rect 250142 340058 250226 340294
rect 250462 340058 267906 340294
rect 268142 340058 268226 340294
rect 268462 340058 285906 340294
rect 286142 340058 286226 340294
rect 286462 340058 303906 340294
rect 304142 340058 304226 340294
rect 304462 340058 321906 340294
rect 322142 340058 322226 340294
rect 322462 340058 339906 340294
rect 340142 340058 340226 340294
rect 340462 340058 357906 340294
rect 358142 340058 358226 340294
rect 358462 340058 375906 340294
rect 376142 340058 376226 340294
rect 376462 340058 393906 340294
rect 394142 340058 394226 340294
rect 394462 340058 411906 340294
rect 412142 340058 412226 340294
rect 412462 340058 429906 340294
rect 430142 340058 430226 340294
rect 430462 340058 447906 340294
rect 448142 340058 448226 340294
rect 448462 340058 465906 340294
rect 466142 340058 466226 340294
rect 466462 340058 483906 340294
rect 484142 340058 484226 340294
rect 484462 340058 501906 340294
rect 502142 340058 502226 340294
rect 502462 340058 519906 340294
rect 520142 340058 520226 340294
rect 520462 340058 537906 340294
rect 538142 340058 538226 340294
rect 538462 340058 547884 340294
rect 548120 340058 548204 340294
rect 548440 340058 548472 340294
rect -4476 340026 548472 340058
rect -4476 336894 548472 336926
rect -4476 336658 -3484 336894
rect -3248 336658 -3164 336894
rect -2928 336658 12186 336894
rect 12422 336658 12506 336894
rect 12742 336658 30186 336894
rect 30422 336658 30506 336894
rect 30742 336658 48186 336894
rect 48422 336658 48506 336894
rect 48742 336658 66186 336894
rect 66422 336658 66506 336894
rect 66742 336658 84186 336894
rect 84422 336658 84506 336894
rect 84742 336658 102186 336894
rect 102422 336658 102506 336894
rect 102742 336658 120186 336894
rect 120422 336658 120506 336894
rect 120742 336658 138186 336894
rect 138422 336658 138506 336894
rect 138742 336658 156186 336894
rect 156422 336658 156506 336894
rect 156742 336658 174186 336894
rect 174422 336658 174506 336894
rect 174742 336658 192186 336894
rect 192422 336658 192506 336894
rect 192742 336658 210186 336894
rect 210422 336658 210506 336894
rect 210742 336658 228186 336894
rect 228422 336658 228506 336894
rect 228742 336658 246186 336894
rect 246422 336658 246506 336894
rect 246742 336658 264186 336894
rect 264422 336658 264506 336894
rect 264742 336658 282186 336894
rect 282422 336658 282506 336894
rect 282742 336658 300186 336894
rect 300422 336658 300506 336894
rect 300742 336658 318186 336894
rect 318422 336658 318506 336894
rect 318742 336658 336186 336894
rect 336422 336658 336506 336894
rect 336742 336658 354186 336894
rect 354422 336658 354506 336894
rect 354742 336658 372186 336894
rect 372422 336658 372506 336894
rect 372742 336658 390186 336894
rect 390422 336658 390506 336894
rect 390742 336658 408186 336894
rect 408422 336658 408506 336894
rect 408742 336658 426186 336894
rect 426422 336658 426506 336894
rect 426742 336658 444186 336894
rect 444422 336658 444506 336894
rect 444742 336658 462186 336894
rect 462422 336658 462506 336894
rect 462742 336658 480186 336894
rect 480422 336658 480506 336894
rect 480742 336658 498186 336894
rect 498422 336658 498506 336894
rect 498742 336658 516186 336894
rect 516422 336658 516506 336894
rect 516742 336658 534186 336894
rect 534422 336658 534506 336894
rect 534742 336658 546924 336894
rect 547160 336658 547244 336894
rect 547480 336658 548472 336894
rect -4476 336574 548472 336658
rect -4476 336338 -3484 336574
rect -3248 336338 -3164 336574
rect -2928 336338 12186 336574
rect 12422 336338 12506 336574
rect 12742 336338 30186 336574
rect 30422 336338 30506 336574
rect 30742 336338 48186 336574
rect 48422 336338 48506 336574
rect 48742 336338 66186 336574
rect 66422 336338 66506 336574
rect 66742 336338 84186 336574
rect 84422 336338 84506 336574
rect 84742 336338 102186 336574
rect 102422 336338 102506 336574
rect 102742 336338 120186 336574
rect 120422 336338 120506 336574
rect 120742 336338 138186 336574
rect 138422 336338 138506 336574
rect 138742 336338 156186 336574
rect 156422 336338 156506 336574
rect 156742 336338 174186 336574
rect 174422 336338 174506 336574
rect 174742 336338 192186 336574
rect 192422 336338 192506 336574
rect 192742 336338 210186 336574
rect 210422 336338 210506 336574
rect 210742 336338 228186 336574
rect 228422 336338 228506 336574
rect 228742 336338 246186 336574
rect 246422 336338 246506 336574
rect 246742 336338 264186 336574
rect 264422 336338 264506 336574
rect 264742 336338 282186 336574
rect 282422 336338 282506 336574
rect 282742 336338 300186 336574
rect 300422 336338 300506 336574
rect 300742 336338 318186 336574
rect 318422 336338 318506 336574
rect 318742 336338 336186 336574
rect 336422 336338 336506 336574
rect 336742 336338 354186 336574
rect 354422 336338 354506 336574
rect 354742 336338 372186 336574
rect 372422 336338 372506 336574
rect 372742 336338 390186 336574
rect 390422 336338 390506 336574
rect 390742 336338 408186 336574
rect 408422 336338 408506 336574
rect 408742 336338 426186 336574
rect 426422 336338 426506 336574
rect 426742 336338 444186 336574
rect 444422 336338 444506 336574
rect 444742 336338 462186 336574
rect 462422 336338 462506 336574
rect 462742 336338 480186 336574
rect 480422 336338 480506 336574
rect 480742 336338 498186 336574
rect 498422 336338 498506 336574
rect 498742 336338 516186 336574
rect 516422 336338 516506 336574
rect 516742 336338 534186 336574
rect 534422 336338 534506 336574
rect 534742 336338 546924 336574
rect 547160 336338 547244 336574
rect 547480 336338 548472 336574
rect -4476 336306 548472 336338
rect -4476 333174 548472 333206
rect -4476 332938 -2524 333174
rect -2288 332938 -2204 333174
rect -1968 332938 8466 333174
rect 8702 332938 8786 333174
rect 9022 332938 26466 333174
rect 26702 332938 26786 333174
rect 27022 332938 44466 333174
rect 44702 332938 44786 333174
rect 45022 332938 62466 333174
rect 62702 332938 62786 333174
rect 63022 332938 80466 333174
rect 80702 332938 80786 333174
rect 81022 332938 98466 333174
rect 98702 332938 98786 333174
rect 99022 332938 116466 333174
rect 116702 332938 116786 333174
rect 117022 332938 134466 333174
rect 134702 332938 134786 333174
rect 135022 332938 152466 333174
rect 152702 332938 152786 333174
rect 153022 332938 170466 333174
rect 170702 332938 170786 333174
rect 171022 332938 188466 333174
rect 188702 332938 188786 333174
rect 189022 332938 206466 333174
rect 206702 332938 206786 333174
rect 207022 332938 224466 333174
rect 224702 332938 224786 333174
rect 225022 332938 242466 333174
rect 242702 332938 242786 333174
rect 243022 332938 260466 333174
rect 260702 332938 260786 333174
rect 261022 332938 278466 333174
rect 278702 332938 278786 333174
rect 279022 332938 296466 333174
rect 296702 332938 296786 333174
rect 297022 332938 314466 333174
rect 314702 332938 314786 333174
rect 315022 332938 332466 333174
rect 332702 332938 332786 333174
rect 333022 332938 350466 333174
rect 350702 332938 350786 333174
rect 351022 332938 368466 333174
rect 368702 332938 368786 333174
rect 369022 332938 386466 333174
rect 386702 332938 386786 333174
rect 387022 332938 404466 333174
rect 404702 332938 404786 333174
rect 405022 332938 422466 333174
rect 422702 332938 422786 333174
rect 423022 332938 440466 333174
rect 440702 332938 440786 333174
rect 441022 332938 458466 333174
rect 458702 332938 458786 333174
rect 459022 332938 476466 333174
rect 476702 332938 476786 333174
rect 477022 332938 494466 333174
rect 494702 332938 494786 333174
rect 495022 332938 512466 333174
rect 512702 332938 512786 333174
rect 513022 332938 530466 333174
rect 530702 332938 530786 333174
rect 531022 332938 545964 333174
rect 546200 332938 546284 333174
rect 546520 332938 548472 333174
rect -4476 332854 548472 332938
rect -4476 332618 -2524 332854
rect -2288 332618 -2204 332854
rect -1968 332618 8466 332854
rect 8702 332618 8786 332854
rect 9022 332618 26466 332854
rect 26702 332618 26786 332854
rect 27022 332618 44466 332854
rect 44702 332618 44786 332854
rect 45022 332618 62466 332854
rect 62702 332618 62786 332854
rect 63022 332618 80466 332854
rect 80702 332618 80786 332854
rect 81022 332618 98466 332854
rect 98702 332618 98786 332854
rect 99022 332618 116466 332854
rect 116702 332618 116786 332854
rect 117022 332618 134466 332854
rect 134702 332618 134786 332854
rect 135022 332618 152466 332854
rect 152702 332618 152786 332854
rect 153022 332618 170466 332854
rect 170702 332618 170786 332854
rect 171022 332618 188466 332854
rect 188702 332618 188786 332854
rect 189022 332618 206466 332854
rect 206702 332618 206786 332854
rect 207022 332618 224466 332854
rect 224702 332618 224786 332854
rect 225022 332618 242466 332854
rect 242702 332618 242786 332854
rect 243022 332618 260466 332854
rect 260702 332618 260786 332854
rect 261022 332618 278466 332854
rect 278702 332618 278786 332854
rect 279022 332618 296466 332854
rect 296702 332618 296786 332854
rect 297022 332618 314466 332854
rect 314702 332618 314786 332854
rect 315022 332618 332466 332854
rect 332702 332618 332786 332854
rect 333022 332618 350466 332854
rect 350702 332618 350786 332854
rect 351022 332618 368466 332854
rect 368702 332618 368786 332854
rect 369022 332618 386466 332854
rect 386702 332618 386786 332854
rect 387022 332618 404466 332854
rect 404702 332618 404786 332854
rect 405022 332618 422466 332854
rect 422702 332618 422786 332854
rect 423022 332618 440466 332854
rect 440702 332618 440786 332854
rect 441022 332618 458466 332854
rect 458702 332618 458786 332854
rect 459022 332618 476466 332854
rect 476702 332618 476786 332854
rect 477022 332618 494466 332854
rect 494702 332618 494786 332854
rect 495022 332618 512466 332854
rect 512702 332618 512786 332854
rect 513022 332618 530466 332854
rect 530702 332618 530786 332854
rect 531022 332618 545964 332854
rect 546200 332618 546284 332854
rect 546520 332618 548472 332854
rect -4476 332586 548472 332618
rect -4476 329454 548472 329486
rect -4476 329218 -1564 329454
rect -1328 329218 -1244 329454
rect -1008 329218 4746 329454
rect 4982 329218 5066 329454
rect 5302 329218 22746 329454
rect 22982 329218 23066 329454
rect 23302 329218 40746 329454
rect 40982 329218 41066 329454
rect 41302 329218 58746 329454
rect 58982 329218 59066 329454
rect 59302 329218 76746 329454
rect 76982 329218 77066 329454
rect 77302 329218 94746 329454
rect 94982 329218 95066 329454
rect 95302 329218 112746 329454
rect 112982 329218 113066 329454
rect 113302 329218 130746 329454
rect 130982 329218 131066 329454
rect 131302 329218 148746 329454
rect 148982 329218 149066 329454
rect 149302 329218 166746 329454
rect 166982 329218 167066 329454
rect 167302 329218 184746 329454
rect 184982 329218 185066 329454
rect 185302 329218 202746 329454
rect 202982 329218 203066 329454
rect 203302 329218 220746 329454
rect 220982 329218 221066 329454
rect 221302 329218 238746 329454
rect 238982 329218 239066 329454
rect 239302 329218 256746 329454
rect 256982 329218 257066 329454
rect 257302 329218 274746 329454
rect 274982 329218 275066 329454
rect 275302 329218 292746 329454
rect 292982 329218 293066 329454
rect 293302 329218 310746 329454
rect 310982 329218 311066 329454
rect 311302 329218 328746 329454
rect 328982 329218 329066 329454
rect 329302 329218 346746 329454
rect 346982 329218 347066 329454
rect 347302 329218 364746 329454
rect 364982 329218 365066 329454
rect 365302 329218 382746 329454
rect 382982 329218 383066 329454
rect 383302 329218 400746 329454
rect 400982 329218 401066 329454
rect 401302 329218 418746 329454
rect 418982 329218 419066 329454
rect 419302 329218 436746 329454
rect 436982 329218 437066 329454
rect 437302 329218 454746 329454
rect 454982 329218 455066 329454
rect 455302 329218 472746 329454
rect 472982 329218 473066 329454
rect 473302 329218 490746 329454
rect 490982 329218 491066 329454
rect 491302 329218 508746 329454
rect 508982 329218 509066 329454
rect 509302 329218 526746 329454
rect 526982 329218 527066 329454
rect 527302 329218 545004 329454
rect 545240 329218 545324 329454
rect 545560 329218 548472 329454
rect -4476 329134 548472 329218
rect -4476 328898 -1564 329134
rect -1328 328898 -1244 329134
rect -1008 328898 4746 329134
rect 4982 328898 5066 329134
rect 5302 328898 22746 329134
rect 22982 328898 23066 329134
rect 23302 328898 40746 329134
rect 40982 328898 41066 329134
rect 41302 328898 58746 329134
rect 58982 328898 59066 329134
rect 59302 328898 76746 329134
rect 76982 328898 77066 329134
rect 77302 328898 94746 329134
rect 94982 328898 95066 329134
rect 95302 328898 112746 329134
rect 112982 328898 113066 329134
rect 113302 328898 130746 329134
rect 130982 328898 131066 329134
rect 131302 328898 148746 329134
rect 148982 328898 149066 329134
rect 149302 328898 166746 329134
rect 166982 328898 167066 329134
rect 167302 328898 184746 329134
rect 184982 328898 185066 329134
rect 185302 328898 202746 329134
rect 202982 328898 203066 329134
rect 203302 328898 220746 329134
rect 220982 328898 221066 329134
rect 221302 328898 238746 329134
rect 238982 328898 239066 329134
rect 239302 328898 256746 329134
rect 256982 328898 257066 329134
rect 257302 328898 274746 329134
rect 274982 328898 275066 329134
rect 275302 328898 292746 329134
rect 292982 328898 293066 329134
rect 293302 328898 310746 329134
rect 310982 328898 311066 329134
rect 311302 328898 328746 329134
rect 328982 328898 329066 329134
rect 329302 328898 346746 329134
rect 346982 328898 347066 329134
rect 347302 328898 364746 329134
rect 364982 328898 365066 329134
rect 365302 328898 382746 329134
rect 382982 328898 383066 329134
rect 383302 328898 400746 329134
rect 400982 328898 401066 329134
rect 401302 328898 418746 329134
rect 418982 328898 419066 329134
rect 419302 328898 436746 329134
rect 436982 328898 437066 329134
rect 437302 328898 454746 329134
rect 454982 328898 455066 329134
rect 455302 328898 472746 329134
rect 472982 328898 473066 329134
rect 473302 328898 490746 329134
rect 490982 328898 491066 329134
rect 491302 328898 508746 329134
rect 508982 328898 509066 329134
rect 509302 328898 526746 329134
rect 526982 328898 527066 329134
rect 527302 328898 545004 329134
rect 545240 328898 545324 329134
rect 545560 328898 548472 329134
rect -4476 328866 548472 328898
rect -4476 322614 548472 322646
rect -4476 322378 -4444 322614
rect -4208 322378 -4124 322614
rect -3888 322378 15906 322614
rect 16142 322378 16226 322614
rect 16462 322378 33906 322614
rect 34142 322378 34226 322614
rect 34462 322378 51906 322614
rect 52142 322378 52226 322614
rect 52462 322378 69906 322614
rect 70142 322378 70226 322614
rect 70462 322378 87906 322614
rect 88142 322378 88226 322614
rect 88462 322378 105906 322614
rect 106142 322378 106226 322614
rect 106462 322378 123906 322614
rect 124142 322378 124226 322614
rect 124462 322378 141906 322614
rect 142142 322378 142226 322614
rect 142462 322378 159906 322614
rect 160142 322378 160226 322614
rect 160462 322378 177906 322614
rect 178142 322378 178226 322614
rect 178462 322378 195906 322614
rect 196142 322378 196226 322614
rect 196462 322378 213906 322614
rect 214142 322378 214226 322614
rect 214462 322378 231906 322614
rect 232142 322378 232226 322614
rect 232462 322378 249906 322614
rect 250142 322378 250226 322614
rect 250462 322378 267906 322614
rect 268142 322378 268226 322614
rect 268462 322378 285906 322614
rect 286142 322378 286226 322614
rect 286462 322378 303906 322614
rect 304142 322378 304226 322614
rect 304462 322378 321906 322614
rect 322142 322378 322226 322614
rect 322462 322378 339906 322614
rect 340142 322378 340226 322614
rect 340462 322378 357906 322614
rect 358142 322378 358226 322614
rect 358462 322378 375906 322614
rect 376142 322378 376226 322614
rect 376462 322378 393906 322614
rect 394142 322378 394226 322614
rect 394462 322378 411906 322614
rect 412142 322378 412226 322614
rect 412462 322378 429906 322614
rect 430142 322378 430226 322614
rect 430462 322378 447906 322614
rect 448142 322378 448226 322614
rect 448462 322378 465906 322614
rect 466142 322378 466226 322614
rect 466462 322378 483906 322614
rect 484142 322378 484226 322614
rect 484462 322378 501906 322614
rect 502142 322378 502226 322614
rect 502462 322378 519906 322614
rect 520142 322378 520226 322614
rect 520462 322378 537906 322614
rect 538142 322378 538226 322614
rect 538462 322378 547884 322614
rect 548120 322378 548204 322614
rect 548440 322378 548472 322614
rect -4476 322294 548472 322378
rect -4476 322058 -4444 322294
rect -4208 322058 -4124 322294
rect -3888 322058 15906 322294
rect 16142 322058 16226 322294
rect 16462 322058 33906 322294
rect 34142 322058 34226 322294
rect 34462 322058 51906 322294
rect 52142 322058 52226 322294
rect 52462 322058 69906 322294
rect 70142 322058 70226 322294
rect 70462 322058 87906 322294
rect 88142 322058 88226 322294
rect 88462 322058 105906 322294
rect 106142 322058 106226 322294
rect 106462 322058 123906 322294
rect 124142 322058 124226 322294
rect 124462 322058 141906 322294
rect 142142 322058 142226 322294
rect 142462 322058 159906 322294
rect 160142 322058 160226 322294
rect 160462 322058 177906 322294
rect 178142 322058 178226 322294
rect 178462 322058 195906 322294
rect 196142 322058 196226 322294
rect 196462 322058 213906 322294
rect 214142 322058 214226 322294
rect 214462 322058 231906 322294
rect 232142 322058 232226 322294
rect 232462 322058 249906 322294
rect 250142 322058 250226 322294
rect 250462 322058 267906 322294
rect 268142 322058 268226 322294
rect 268462 322058 285906 322294
rect 286142 322058 286226 322294
rect 286462 322058 303906 322294
rect 304142 322058 304226 322294
rect 304462 322058 321906 322294
rect 322142 322058 322226 322294
rect 322462 322058 339906 322294
rect 340142 322058 340226 322294
rect 340462 322058 357906 322294
rect 358142 322058 358226 322294
rect 358462 322058 375906 322294
rect 376142 322058 376226 322294
rect 376462 322058 393906 322294
rect 394142 322058 394226 322294
rect 394462 322058 411906 322294
rect 412142 322058 412226 322294
rect 412462 322058 429906 322294
rect 430142 322058 430226 322294
rect 430462 322058 447906 322294
rect 448142 322058 448226 322294
rect 448462 322058 465906 322294
rect 466142 322058 466226 322294
rect 466462 322058 483906 322294
rect 484142 322058 484226 322294
rect 484462 322058 501906 322294
rect 502142 322058 502226 322294
rect 502462 322058 519906 322294
rect 520142 322058 520226 322294
rect 520462 322058 537906 322294
rect 538142 322058 538226 322294
rect 538462 322058 547884 322294
rect 548120 322058 548204 322294
rect 548440 322058 548472 322294
rect -4476 322026 548472 322058
rect -4476 318894 548472 318926
rect -4476 318658 -3484 318894
rect -3248 318658 -3164 318894
rect -2928 318658 12186 318894
rect 12422 318658 12506 318894
rect 12742 318658 30186 318894
rect 30422 318658 30506 318894
rect 30742 318658 48186 318894
rect 48422 318658 48506 318894
rect 48742 318658 66186 318894
rect 66422 318658 66506 318894
rect 66742 318658 84186 318894
rect 84422 318658 84506 318894
rect 84742 318658 102186 318894
rect 102422 318658 102506 318894
rect 102742 318658 120186 318894
rect 120422 318658 120506 318894
rect 120742 318658 138186 318894
rect 138422 318658 138506 318894
rect 138742 318658 156186 318894
rect 156422 318658 156506 318894
rect 156742 318658 174186 318894
rect 174422 318658 174506 318894
rect 174742 318658 192186 318894
rect 192422 318658 192506 318894
rect 192742 318658 210186 318894
rect 210422 318658 210506 318894
rect 210742 318658 228186 318894
rect 228422 318658 228506 318894
rect 228742 318658 246186 318894
rect 246422 318658 246506 318894
rect 246742 318658 264186 318894
rect 264422 318658 264506 318894
rect 264742 318658 282186 318894
rect 282422 318658 282506 318894
rect 282742 318658 300186 318894
rect 300422 318658 300506 318894
rect 300742 318658 318186 318894
rect 318422 318658 318506 318894
rect 318742 318658 336186 318894
rect 336422 318658 336506 318894
rect 336742 318658 354186 318894
rect 354422 318658 354506 318894
rect 354742 318658 372186 318894
rect 372422 318658 372506 318894
rect 372742 318658 390186 318894
rect 390422 318658 390506 318894
rect 390742 318658 408186 318894
rect 408422 318658 408506 318894
rect 408742 318658 426186 318894
rect 426422 318658 426506 318894
rect 426742 318658 444186 318894
rect 444422 318658 444506 318894
rect 444742 318658 462186 318894
rect 462422 318658 462506 318894
rect 462742 318658 480186 318894
rect 480422 318658 480506 318894
rect 480742 318658 498186 318894
rect 498422 318658 498506 318894
rect 498742 318658 516186 318894
rect 516422 318658 516506 318894
rect 516742 318658 534186 318894
rect 534422 318658 534506 318894
rect 534742 318658 546924 318894
rect 547160 318658 547244 318894
rect 547480 318658 548472 318894
rect -4476 318574 548472 318658
rect -4476 318338 -3484 318574
rect -3248 318338 -3164 318574
rect -2928 318338 12186 318574
rect 12422 318338 12506 318574
rect 12742 318338 30186 318574
rect 30422 318338 30506 318574
rect 30742 318338 48186 318574
rect 48422 318338 48506 318574
rect 48742 318338 66186 318574
rect 66422 318338 66506 318574
rect 66742 318338 84186 318574
rect 84422 318338 84506 318574
rect 84742 318338 102186 318574
rect 102422 318338 102506 318574
rect 102742 318338 120186 318574
rect 120422 318338 120506 318574
rect 120742 318338 138186 318574
rect 138422 318338 138506 318574
rect 138742 318338 156186 318574
rect 156422 318338 156506 318574
rect 156742 318338 174186 318574
rect 174422 318338 174506 318574
rect 174742 318338 192186 318574
rect 192422 318338 192506 318574
rect 192742 318338 210186 318574
rect 210422 318338 210506 318574
rect 210742 318338 228186 318574
rect 228422 318338 228506 318574
rect 228742 318338 246186 318574
rect 246422 318338 246506 318574
rect 246742 318338 264186 318574
rect 264422 318338 264506 318574
rect 264742 318338 282186 318574
rect 282422 318338 282506 318574
rect 282742 318338 300186 318574
rect 300422 318338 300506 318574
rect 300742 318338 318186 318574
rect 318422 318338 318506 318574
rect 318742 318338 336186 318574
rect 336422 318338 336506 318574
rect 336742 318338 354186 318574
rect 354422 318338 354506 318574
rect 354742 318338 372186 318574
rect 372422 318338 372506 318574
rect 372742 318338 390186 318574
rect 390422 318338 390506 318574
rect 390742 318338 408186 318574
rect 408422 318338 408506 318574
rect 408742 318338 426186 318574
rect 426422 318338 426506 318574
rect 426742 318338 444186 318574
rect 444422 318338 444506 318574
rect 444742 318338 462186 318574
rect 462422 318338 462506 318574
rect 462742 318338 480186 318574
rect 480422 318338 480506 318574
rect 480742 318338 498186 318574
rect 498422 318338 498506 318574
rect 498742 318338 516186 318574
rect 516422 318338 516506 318574
rect 516742 318338 534186 318574
rect 534422 318338 534506 318574
rect 534742 318338 546924 318574
rect 547160 318338 547244 318574
rect 547480 318338 548472 318574
rect -4476 318306 548472 318338
rect -4476 315174 548472 315206
rect -4476 314938 -2524 315174
rect -2288 314938 -2204 315174
rect -1968 314938 8466 315174
rect 8702 314938 8786 315174
rect 9022 314938 26466 315174
rect 26702 314938 26786 315174
rect 27022 314938 44466 315174
rect 44702 314938 44786 315174
rect 45022 314938 62466 315174
rect 62702 314938 62786 315174
rect 63022 314938 80466 315174
rect 80702 314938 80786 315174
rect 81022 314938 98466 315174
rect 98702 314938 98786 315174
rect 99022 314938 116466 315174
rect 116702 314938 116786 315174
rect 117022 314938 134466 315174
rect 134702 314938 134786 315174
rect 135022 314938 152466 315174
rect 152702 314938 152786 315174
rect 153022 314938 170466 315174
rect 170702 314938 170786 315174
rect 171022 314938 188466 315174
rect 188702 314938 188786 315174
rect 189022 314938 206466 315174
rect 206702 314938 206786 315174
rect 207022 314938 224466 315174
rect 224702 314938 224786 315174
rect 225022 314938 242466 315174
rect 242702 314938 242786 315174
rect 243022 314938 260466 315174
rect 260702 314938 260786 315174
rect 261022 314938 278466 315174
rect 278702 314938 278786 315174
rect 279022 314938 296466 315174
rect 296702 314938 296786 315174
rect 297022 314938 314466 315174
rect 314702 314938 314786 315174
rect 315022 314938 332466 315174
rect 332702 314938 332786 315174
rect 333022 314938 350466 315174
rect 350702 314938 350786 315174
rect 351022 314938 368466 315174
rect 368702 314938 368786 315174
rect 369022 314938 386466 315174
rect 386702 314938 386786 315174
rect 387022 314938 404466 315174
rect 404702 314938 404786 315174
rect 405022 314938 422466 315174
rect 422702 314938 422786 315174
rect 423022 314938 440466 315174
rect 440702 314938 440786 315174
rect 441022 314938 458466 315174
rect 458702 314938 458786 315174
rect 459022 314938 476466 315174
rect 476702 314938 476786 315174
rect 477022 314938 494466 315174
rect 494702 314938 494786 315174
rect 495022 314938 512466 315174
rect 512702 314938 512786 315174
rect 513022 314938 530466 315174
rect 530702 314938 530786 315174
rect 531022 314938 545964 315174
rect 546200 314938 546284 315174
rect 546520 314938 548472 315174
rect -4476 314854 548472 314938
rect -4476 314618 -2524 314854
rect -2288 314618 -2204 314854
rect -1968 314618 8466 314854
rect 8702 314618 8786 314854
rect 9022 314618 26466 314854
rect 26702 314618 26786 314854
rect 27022 314618 44466 314854
rect 44702 314618 44786 314854
rect 45022 314618 62466 314854
rect 62702 314618 62786 314854
rect 63022 314618 80466 314854
rect 80702 314618 80786 314854
rect 81022 314618 98466 314854
rect 98702 314618 98786 314854
rect 99022 314618 116466 314854
rect 116702 314618 116786 314854
rect 117022 314618 134466 314854
rect 134702 314618 134786 314854
rect 135022 314618 152466 314854
rect 152702 314618 152786 314854
rect 153022 314618 170466 314854
rect 170702 314618 170786 314854
rect 171022 314618 188466 314854
rect 188702 314618 188786 314854
rect 189022 314618 206466 314854
rect 206702 314618 206786 314854
rect 207022 314618 224466 314854
rect 224702 314618 224786 314854
rect 225022 314618 242466 314854
rect 242702 314618 242786 314854
rect 243022 314618 260466 314854
rect 260702 314618 260786 314854
rect 261022 314618 278466 314854
rect 278702 314618 278786 314854
rect 279022 314618 296466 314854
rect 296702 314618 296786 314854
rect 297022 314618 314466 314854
rect 314702 314618 314786 314854
rect 315022 314618 332466 314854
rect 332702 314618 332786 314854
rect 333022 314618 350466 314854
rect 350702 314618 350786 314854
rect 351022 314618 368466 314854
rect 368702 314618 368786 314854
rect 369022 314618 386466 314854
rect 386702 314618 386786 314854
rect 387022 314618 404466 314854
rect 404702 314618 404786 314854
rect 405022 314618 422466 314854
rect 422702 314618 422786 314854
rect 423022 314618 440466 314854
rect 440702 314618 440786 314854
rect 441022 314618 458466 314854
rect 458702 314618 458786 314854
rect 459022 314618 476466 314854
rect 476702 314618 476786 314854
rect 477022 314618 494466 314854
rect 494702 314618 494786 314854
rect 495022 314618 512466 314854
rect 512702 314618 512786 314854
rect 513022 314618 530466 314854
rect 530702 314618 530786 314854
rect 531022 314618 545964 314854
rect 546200 314618 546284 314854
rect 546520 314618 548472 314854
rect -4476 314586 548472 314618
rect -4476 311454 548472 311486
rect -4476 311218 -1564 311454
rect -1328 311218 -1244 311454
rect -1008 311218 4746 311454
rect 4982 311218 5066 311454
rect 5302 311218 22746 311454
rect 22982 311218 23066 311454
rect 23302 311218 40746 311454
rect 40982 311218 41066 311454
rect 41302 311218 58746 311454
rect 58982 311218 59066 311454
rect 59302 311218 76746 311454
rect 76982 311218 77066 311454
rect 77302 311218 94746 311454
rect 94982 311218 95066 311454
rect 95302 311218 112746 311454
rect 112982 311218 113066 311454
rect 113302 311218 130746 311454
rect 130982 311218 131066 311454
rect 131302 311218 148746 311454
rect 148982 311218 149066 311454
rect 149302 311218 166746 311454
rect 166982 311218 167066 311454
rect 167302 311218 184746 311454
rect 184982 311218 185066 311454
rect 185302 311218 202746 311454
rect 202982 311218 203066 311454
rect 203302 311218 220746 311454
rect 220982 311218 221066 311454
rect 221302 311218 238746 311454
rect 238982 311218 239066 311454
rect 239302 311218 256746 311454
rect 256982 311218 257066 311454
rect 257302 311218 274746 311454
rect 274982 311218 275066 311454
rect 275302 311218 292746 311454
rect 292982 311218 293066 311454
rect 293302 311218 310746 311454
rect 310982 311218 311066 311454
rect 311302 311218 328746 311454
rect 328982 311218 329066 311454
rect 329302 311218 346746 311454
rect 346982 311218 347066 311454
rect 347302 311218 364746 311454
rect 364982 311218 365066 311454
rect 365302 311218 382746 311454
rect 382982 311218 383066 311454
rect 383302 311218 400746 311454
rect 400982 311218 401066 311454
rect 401302 311218 418746 311454
rect 418982 311218 419066 311454
rect 419302 311218 436746 311454
rect 436982 311218 437066 311454
rect 437302 311218 454746 311454
rect 454982 311218 455066 311454
rect 455302 311218 472746 311454
rect 472982 311218 473066 311454
rect 473302 311218 490746 311454
rect 490982 311218 491066 311454
rect 491302 311218 508746 311454
rect 508982 311218 509066 311454
rect 509302 311218 526746 311454
rect 526982 311218 527066 311454
rect 527302 311218 545004 311454
rect 545240 311218 545324 311454
rect 545560 311218 548472 311454
rect -4476 311134 548472 311218
rect -4476 310898 -1564 311134
rect -1328 310898 -1244 311134
rect -1008 310898 4746 311134
rect 4982 310898 5066 311134
rect 5302 310898 22746 311134
rect 22982 310898 23066 311134
rect 23302 310898 40746 311134
rect 40982 310898 41066 311134
rect 41302 310898 58746 311134
rect 58982 310898 59066 311134
rect 59302 310898 76746 311134
rect 76982 310898 77066 311134
rect 77302 310898 94746 311134
rect 94982 310898 95066 311134
rect 95302 310898 112746 311134
rect 112982 310898 113066 311134
rect 113302 310898 130746 311134
rect 130982 310898 131066 311134
rect 131302 310898 148746 311134
rect 148982 310898 149066 311134
rect 149302 310898 166746 311134
rect 166982 310898 167066 311134
rect 167302 310898 184746 311134
rect 184982 310898 185066 311134
rect 185302 310898 202746 311134
rect 202982 310898 203066 311134
rect 203302 310898 220746 311134
rect 220982 310898 221066 311134
rect 221302 310898 238746 311134
rect 238982 310898 239066 311134
rect 239302 310898 256746 311134
rect 256982 310898 257066 311134
rect 257302 310898 274746 311134
rect 274982 310898 275066 311134
rect 275302 310898 292746 311134
rect 292982 310898 293066 311134
rect 293302 310898 310746 311134
rect 310982 310898 311066 311134
rect 311302 310898 328746 311134
rect 328982 310898 329066 311134
rect 329302 310898 346746 311134
rect 346982 310898 347066 311134
rect 347302 310898 364746 311134
rect 364982 310898 365066 311134
rect 365302 310898 382746 311134
rect 382982 310898 383066 311134
rect 383302 310898 400746 311134
rect 400982 310898 401066 311134
rect 401302 310898 418746 311134
rect 418982 310898 419066 311134
rect 419302 310898 436746 311134
rect 436982 310898 437066 311134
rect 437302 310898 454746 311134
rect 454982 310898 455066 311134
rect 455302 310898 472746 311134
rect 472982 310898 473066 311134
rect 473302 310898 490746 311134
rect 490982 310898 491066 311134
rect 491302 310898 508746 311134
rect 508982 310898 509066 311134
rect 509302 310898 526746 311134
rect 526982 310898 527066 311134
rect 527302 310898 545004 311134
rect 545240 310898 545324 311134
rect 545560 310898 548472 311134
rect -4476 310866 548472 310898
rect -4476 304614 548472 304646
rect -4476 304378 -4444 304614
rect -4208 304378 -4124 304614
rect -3888 304378 15906 304614
rect 16142 304378 16226 304614
rect 16462 304378 33906 304614
rect 34142 304378 34226 304614
rect 34462 304378 51906 304614
rect 52142 304378 52226 304614
rect 52462 304378 69906 304614
rect 70142 304378 70226 304614
rect 70462 304378 87906 304614
rect 88142 304378 88226 304614
rect 88462 304378 105906 304614
rect 106142 304378 106226 304614
rect 106462 304378 123906 304614
rect 124142 304378 124226 304614
rect 124462 304378 141906 304614
rect 142142 304378 142226 304614
rect 142462 304378 159906 304614
rect 160142 304378 160226 304614
rect 160462 304378 177906 304614
rect 178142 304378 178226 304614
rect 178462 304378 195906 304614
rect 196142 304378 196226 304614
rect 196462 304378 213906 304614
rect 214142 304378 214226 304614
rect 214462 304378 231906 304614
rect 232142 304378 232226 304614
rect 232462 304378 249906 304614
rect 250142 304378 250226 304614
rect 250462 304378 267906 304614
rect 268142 304378 268226 304614
rect 268462 304378 285906 304614
rect 286142 304378 286226 304614
rect 286462 304378 303906 304614
rect 304142 304378 304226 304614
rect 304462 304378 321906 304614
rect 322142 304378 322226 304614
rect 322462 304378 339906 304614
rect 340142 304378 340226 304614
rect 340462 304378 357906 304614
rect 358142 304378 358226 304614
rect 358462 304378 375906 304614
rect 376142 304378 376226 304614
rect 376462 304378 393906 304614
rect 394142 304378 394226 304614
rect 394462 304378 411906 304614
rect 412142 304378 412226 304614
rect 412462 304378 429906 304614
rect 430142 304378 430226 304614
rect 430462 304378 447906 304614
rect 448142 304378 448226 304614
rect 448462 304378 465906 304614
rect 466142 304378 466226 304614
rect 466462 304378 483906 304614
rect 484142 304378 484226 304614
rect 484462 304378 501906 304614
rect 502142 304378 502226 304614
rect 502462 304378 519906 304614
rect 520142 304378 520226 304614
rect 520462 304378 537906 304614
rect 538142 304378 538226 304614
rect 538462 304378 547884 304614
rect 548120 304378 548204 304614
rect 548440 304378 548472 304614
rect -4476 304294 548472 304378
rect -4476 304058 -4444 304294
rect -4208 304058 -4124 304294
rect -3888 304058 15906 304294
rect 16142 304058 16226 304294
rect 16462 304058 33906 304294
rect 34142 304058 34226 304294
rect 34462 304058 51906 304294
rect 52142 304058 52226 304294
rect 52462 304058 69906 304294
rect 70142 304058 70226 304294
rect 70462 304058 87906 304294
rect 88142 304058 88226 304294
rect 88462 304058 105906 304294
rect 106142 304058 106226 304294
rect 106462 304058 123906 304294
rect 124142 304058 124226 304294
rect 124462 304058 141906 304294
rect 142142 304058 142226 304294
rect 142462 304058 159906 304294
rect 160142 304058 160226 304294
rect 160462 304058 177906 304294
rect 178142 304058 178226 304294
rect 178462 304058 195906 304294
rect 196142 304058 196226 304294
rect 196462 304058 213906 304294
rect 214142 304058 214226 304294
rect 214462 304058 231906 304294
rect 232142 304058 232226 304294
rect 232462 304058 249906 304294
rect 250142 304058 250226 304294
rect 250462 304058 267906 304294
rect 268142 304058 268226 304294
rect 268462 304058 285906 304294
rect 286142 304058 286226 304294
rect 286462 304058 303906 304294
rect 304142 304058 304226 304294
rect 304462 304058 321906 304294
rect 322142 304058 322226 304294
rect 322462 304058 339906 304294
rect 340142 304058 340226 304294
rect 340462 304058 357906 304294
rect 358142 304058 358226 304294
rect 358462 304058 375906 304294
rect 376142 304058 376226 304294
rect 376462 304058 393906 304294
rect 394142 304058 394226 304294
rect 394462 304058 411906 304294
rect 412142 304058 412226 304294
rect 412462 304058 429906 304294
rect 430142 304058 430226 304294
rect 430462 304058 447906 304294
rect 448142 304058 448226 304294
rect 448462 304058 465906 304294
rect 466142 304058 466226 304294
rect 466462 304058 483906 304294
rect 484142 304058 484226 304294
rect 484462 304058 501906 304294
rect 502142 304058 502226 304294
rect 502462 304058 519906 304294
rect 520142 304058 520226 304294
rect 520462 304058 537906 304294
rect 538142 304058 538226 304294
rect 538462 304058 547884 304294
rect 548120 304058 548204 304294
rect 548440 304058 548472 304294
rect -4476 304026 548472 304058
rect -4476 300894 548472 300926
rect -4476 300658 -3484 300894
rect -3248 300658 -3164 300894
rect -2928 300658 12186 300894
rect 12422 300658 12506 300894
rect 12742 300658 30186 300894
rect 30422 300658 30506 300894
rect 30742 300658 48186 300894
rect 48422 300658 48506 300894
rect 48742 300658 66186 300894
rect 66422 300658 66506 300894
rect 66742 300658 84186 300894
rect 84422 300658 84506 300894
rect 84742 300658 102186 300894
rect 102422 300658 102506 300894
rect 102742 300658 120186 300894
rect 120422 300658 120506 300894
rect 120742 300658 138186 300894
rect 138422 300658 138506 300894
rect 138742 300658 156186 300894
rect 156422 300658 156506 300894
rect 156742 300658 174186 300894
rect 174422 300658 174506 300894
rect 174742 300658 192186 300894
rect 192422 300658 192506 300894
rect 192742 300658 210186 300894
rect 210422 300658 210506 300894
rect 210742 300658 228186 300894
rect 228422 300658 228506 300894
rect 228742 300658 246186 300894
rect 246422 300658 246506 300894
rect 246742 300658 264186 300894
rect 264422 300658 264506 300894
rect 264742 300658 282186 300894
rect 282422 300658 282506 300894
rect 282742 300658 300186 300894
rect 300422 300658 300506 300894
rect 300742 300658 318186 300894
rect 318422 300658 318506 300894
rect 318742 300658 336186 300894
rect 336422 300658 336506 300894
rect 336742 300658 354186 300894
rect 354422 300658 354506 300894
rect 354742 300658 372186 300894
rect 372422 300658 372506 300894
rect 372742 300658 390186 300894
rect 390422 300658 390506 300894
rect 390742 300658 408186 300894
rect 408422 300658 408506 300894
rect 408742 300658 426186 300894
rect 426422 300658 426506 300894
rect 426742 300658 444186 300894
rect 444422 300658 444506 300894
rect 444742 300658 462186 300894
rect 462422 300658 462506 300894
rect 462742 300658 480186 300894
rect 480422 300658 480506 300894
rect 480742 300658 498186 300894
rect 498422 300658 498506 300894
rect 498742 300658 516186 300894
rect 516422 300658 516506 300894
rect 516742 300658 534186 300894
rect 534422 300658 534506 300894
rect 534742 300658 546924 300894
rect 547160 300658 547244 300894
rect 547480 300658 548472 300894
rect -4476 300574 548472 300658
rect -4476 300338 -3484 300574
rect -3248 300338 -3164 300574
rect -2928 300338 12186 300574
rect 12422 300338 12506 300574
rect 12742 300338 30186 300574
rect 30422 300338 30506 300574
rect 30742 300338 48186 300574
rect 48422 300338 48506 300574
rect 48742 300338 66186 300574
rect 66422 300338 66506 300574
rect 66742 300338 84186 300574
rect 84422 300338 84506 300574
rect 84742 300338 102186 300574
rect 102422 300338 102506 300574
rect 102742 300338 120186 300574
rect 120422 300338 120506 300574
rect 120742 300338 138186 300574
rect 138422 300338 138506 300574
rect 138742 300338 156186 300574
rect 156422 300338 156506 300574
rect 156742 300338 174186 300574
rect 174422 300338 174506 300574
rect 174742 300338 192186 300574
rect 192422 300338 192506 300574
rect 192742 300338 210186 300574
rect 210422 300338 210506 300574
rect 210742 300338 228186 300574
rect 228422 300338 228506 300574
rect 228742 300338 246186 300574
rect 246422 300338 246506 300574
rect 246742 300338 264186 300574
rect 264422 300338 264506 300574
rect 264742 300338 282186 300574
rect 282422 300338 282506 300574
rect 282742 300338 300186 300574
rect 300422 300338 300506 300574
rect 300742 300338 318186 300574
rect 318422 300338 318506 300574
rect 318742 300338 336186 300574
rect 336422 300338 336506 300574
rect 336742 300338 354186 300574
rect 354422 300338 354506 300574
rect 354742 300338 372186 300574
rect 372422 300338 372506 300574
rect 372742 300338 390186 300574
rect 390422 300338 390506 300574
rect 390742 300338 408186 300574
rect 408422 300338 408506 300574
rect 408742 300338 426186 300574
rect 426422 300338 426506 300574
rect 426742 300338 444186 300574
rect 444422 300338 444506 300574
rect 444742 300338 462186 300574
rect 462422 300338 462506 300574
rect 462742 300338 480186 300574
rect 480422 300338 480506 300574
rect 480742 300338 498186 300574
rect 498422 300338 498506 300574
rect 498742 300338 516186 300574
rect 516422 300338 516506 300574
rect 516742 300338 534186 300574
rect 534422 300338 534506 300574
rect 534742 300338 546924 300574
rect 547160 300338 547244 300574
rect 547480 300338 548472 300574
rect -4476 300306 548472 300338
rect -4476 297174 548472 297206
rect -4476 296938 -2524 297174
rect -2288 296938 -2204 297174
rect -1968 296938 8466 297174
rect 8702 296938 8786 297174
rect 9022 296938 26466 297174
rect 26702 296938 26786 297174
rect 27022 296938 44466 297174
rect 44702 296938 44786 297174
rect 45022 296938 62466 297174
rect 62702 296938 62786 297174
rect 63022 296938 80466 297174
rect 80702 296938 80786 297174
rect 81022 296938 98466 297174
rect 98702 296938 98786 297174
rect 99022 296938 116466 297174
rect 116702 296938 116786 297174
rect 117022 296938 134466 297174
rect 134702 296938 134786 297174
rect 135022 296938 152466 297174
rect 152702 296938 152786 297174
rect 153022 296938 170466 297174
rect 170702 296938 170786 297174
rect 171022 296938 188466 297174
rect 188702 296938 188786 297174
rect 189022 296938 206466 297174
rect 206702 296938 206786 297174
rect 207022 296938 224466 297174
rect 224702 296938 224786 297174
rect 225022 296938 242466 297174
rect 242702 296938 242786 297174
rect 243022 296938 260466 297174
rect 260702 296938 260786 297174
rect 261022 296938 278466 297174
rect 278702 296938 278786 297174
rect 279022 296938 296466 297174
rect 296702 296938 296786 297174
rect 297022 296938 314466 297174
rect 314702 296938 314786 297174
rect 315022 296938 332466 297174
rect 332702 296938 332786 297174
rect 333022 296938 350466 297174
rect 350702 296938 350786 297174
rect 351022 296938 368466 297174
rect 368702 296938 368786 297174
rect 369022 296938 386466 297174
rect 386702 296938 386786 297174
rect 387022 296938 404466 297174
rect 404702 296938 404786 297174
rect 405022 296938 422466 297174
rect 422702 296938 422786 297174
rect 423022 296938 440466 297174
rect 440702 296938 440786 297174
rect 441022 296938 458466 297174
rect 458702 296938 458786 297174
rect 459022 296938 476466 297174
rect 476702 296938 476786 297174
rect 477022 296938 494466 297174
rect 494702 296938 494786 297174
rect 495022 296938 512466 297174
rect 512702 296938 512786 297174
rect 513022 296938 530466 297174
rect 530702 296938 530786 297174
rect 531022 296938 545964 297174
rect 546200 296938 546284 297174
rect 546520 296938 548472 297174
rect -4476 296854 548472 296938
rect -4476 296618 -2524 296854
rect -2288 296618 -2204 296854
rect -1968 296618 8466 296854
rect 8702 296618 8786 296854
rect 9022 296618 26466 296854
rect 26702 296618 26786 296854
rect 27022 296618 44466 296854
rect 44702 296618 44786 296854
rect 45022 296618 62466 296854
rect 62702 296618 62786 296854
rect 63022 296618 80466 296854
rect 80702 296618 80786 296854
rect 81022 296618 98466 296854
rect 98702 296618 98786 296854
rect 99022 296618 116466 296854
rect 116702 296618 116786 296854
rect 117022 296618 134466 296854
rect 134702 296618 134786 296854
rect 135022 296618 152466 296854
rect 152702 296618 152786 296854
rect 153022 296618 170466 296854
rect 170702 296618 170786 296854
rect 171022 296618 188466 296854
rect 188702 296618 188786 296854
rect 189022 296618 206466 296854
rect 206702 296618 206786 296854
rect 207022 296618 224466 296854
rect 224702 296618 224786 296854
rect 225022 296618 242466 296854
rect 242702 296618 242786 296854
rect 243022 296618 260466 296854
rect 260702 296618 260786 296854
rect 261022 296618 278466 296854
rect 278702 296618 278786 296854
rect 279022 296618 296466 296854
rect 296702 296618 296786 296854
rect 297022 296618 314466 296854
rect 314702 296618 314786 296854
rect 315022 296618 332466 296854
rect 332702 296618 332786 296854
rect 333022 296618 350466 296854
rect 350702 296618 350786 296854
rect 351022 296618 368466 296854
rect 368702 296618 368786 296854
rect 369022 296618 386466 296854
rect 386702 296618 386786 296854
rect 387022 296618 404466 296854
rect 404702 296618 404786 296854
rect 405022 296618 422466 296854
rect 422702 296618 422786 296854
rect 423022 296618 440466 296854
rect 440702 296618 440786 296854
rect 441022 296618 458466 296854
rect 458702 296618 458786 296854
rect 459022 296618 476466 296854
rect 476702 296618 476786 296854
rect 477022 296618 494466 296854
rect 494702 296618 494786 296854
rect 495022 296618 512466 296854
rect 512702 296618 512786 296854
rect 513022 296618 530466 296854
rect 530702 296618 530786 296854
rect 531022 296618 545964 296854
rect 546200 296618 546284 296854
rect 546520 296618 548472 296854
rect -4476 296586 548472 296618
rect -4476 293454 548472 293486
rect -4476 293218 -1564 293454
rect -1328 293218 -1244 293454
rect -1008 293218 4746 293454
rect 4982 293218 5066 293454
rect 5302 293218 22746 293454
rect 22982 293218 23066 293454
rect 23302 293218 40746 293454
rect 40982 293218 41066 293454
rect 41302 293218 58746 293454
rect 58982 293218 59066 293454
rect 59302 293218 76746 293454
rect 76982 293218 77066 293454
rect 77302 293218 94746 293454
rect 94982 293218 95066 293454
rect 95302 293218 112746 293454
rect 112982 293218 113066 293454
rect 113302 293218 130746 293454
rect 130982 293218 131066 293454
rect 131302 293218 148746 293454
rect 148982 293218 149066 293454
rect 149302 293218 166746 293454
rect 166982 293218 167066 293454
rect 167302 293218 184746 293454
rect 184982 293218 185066 293454
rect 185302 293218 202746 293454
rect 202982 293218 203066 293454
rect 203302 293218 220746 293454
rect 220982 293218 221066 293454
rect 221302 293218 238746 293454
rect 238982 293218 239066 293454
rect 239302 293218 256746 293454
rect 256982 293218 257066 293454
rect 257302 293218 274746 293454
rect 274982 293218 275066 293454
rect 275302 293218 292746 293454
rect 292982 293218 293066 293454
rect 293302 293218 310746 293454
rect 310982 293218 311066 293454
rect 311302 293218 328746 293454
rect 328982 293218 329066 293454
rect 329302 293218 346746 293454
rect 346982 293218 347066 293454
rect 347302 293218 364746 293454
rect 364982 293218 365066 293454
rect 365302 293218 382746 293454
rect 382982 293218 383066 293454
rect 383302 293218 400746 293454
rect 400982 293218 401066 293454
rect 401302 293218 418746 293454
rect 418982 293218 419066 293454
rect 419302 293218 436746 293454
rect 436982 293218 437066 293454
rect 437302 293218 454746 293454
rect 454982 293218 455066 293454
rect 455302 293218 472746 293454
rect 472982 293218 473066 293454
rect 473302 293218 490746 293454
rect 490982 293218 491066 293454
rect 491302 293218 508746 293454
rect 508982 293218 509066 293454
rect 509302 293218 526746 293454
rect 526982 293218 527066 293454
rect 527302 293218 545004 293454
rect 545240 293218 545324 293454
rect 545560 293218 548472 293454
rect -4476 293134 548472 293218
rect -4476 292898 -1564 293134
rect -1328 292898 -1244 293134
rect -1008 292898 4746 293134
rect 4982 292898 5066 293134
rect 5302 292898 22746 293134
rect 22982 292898 23066 293134
rect 23302 292898 40746 293134
rect 40982 292898 41066 293134
rect 41302 292898 58746 293134
rect 58982 292898 59066 293134
rect 59302 292898 76746 293134
rect 76982 292898 77066 293134
rect 77302 292898 94746 293134
rect 94982 292898 95066 293134
rect 95302 292898 112746 293134
rect 112982 292898 113066 293134
rect 113302 292898 130746 293134
rect 130982 292898 131066 293134
rect 131302 292898 148746 293134
rect 148982 292898 149066 293134
rect 149302 292898 166746 293134
rect 166982 292898 167066 293134
rect 167302 292898 184746 293134
rect 184982 292898 185066 293134
rect 185302 292898 202746 293134
rect 202982 292898 203066 293134
rect 203302 292898 220746 293134
rect 220982 292898 221066 293134
rect 221302 292898 238746 293134
rect 238982 292898 239066 293134
rect 239302 292898 256746 293134
rect 256982 292898 257066 293134
rect 257302 292898 274746 293134
rect 274982 292898 275066 293134
rect 275302 292898 292746 293134
rect 292982 292898 293066 293134
rect 293302 292898 310746 293134
rect 310982 292898 311066 293134
rect 311302 292898 328746 293134
rect 328982 292898 329066 293134
rect 329302 292898 346746 293134
rect 346982 292898 347066 293134
rect 347302 292898 364746 293134
rect 364982 292898 365066 293134
rect 365302 292898 382746 293134
rect 382982 292898 383066 293134
rect 383302 292898 400746 293134
rect 400982 292898 401066 293134
rect 401302 292898 418746 293134
rect 418982 292898 419066 293134
rect 419302 292898 436746 293134
rect 436982 292898 437066 293134
rect 437302 292898 454746 293134
rect 454982 292898 455066 293134
rect 455302 292898 472746 293134
rect 472982 292898 473066 293134
rect 473302 292898 490746 293134
rect 490982 292898 491066 293134
rect 491302 292898 508746 293134
rect 508982 292898 509066 293134
rect 509302 292898 526746 293134
rect 526982 292898 527066 293134
rect 527302 292898 545004 293134
rect 545240 292898 545324 293134
rect 545560 292898 548472 293134
rect -4476 292866 548472 292898
rect -4476 286614 548472 286646
rect -4476 286378 -4444 286614
rect -4208 286378 -4124 286614
rect -3888 286378 15906 286614
rect 16142 286378 16226 286614
rect 16462 286378 33906 286614
rect 34142 286378 34226 286614
rect 34462 286378 51906 286614
rect 52142 286378 52226 286614
rect 52462 286378 69906 286614
rect 70142 286378 70226 286614
rect 70462 286378 87906 286614
rect 88142 286378 88226 286614
rect 88462 286378 105906 286614
rect 106142 286378 106226 286614
rect 106462 286378 123906 286614
rect 124142 286378 124226 286614
rect 124462 286378 141906 286614
rect 142142 286378 142226 286614
rect 142462 286378 159906 286614
rect 160142 286378 160226 286614
rect 160462 286378 177906 286614
rect 178142 286378 178226 286614
rect 178462 286378 195906 286614
rect 196142 286378 196226 286614
rect 196462 286378 213906 286614
rect 214142 286378 214226 286614
rect 214462 286378 231906 286614
rect 232142 286378 232226 286614
rect 232462 286378 249906 286614
rect 250142 286378 250226 286614
rect 250462 286378 267906 286614
rect 268142 286378 268226 286614
rect 268462 286378 285906 286614
rect 286142 286378 286226 286614
rect 286462 286378 303906 286614
rect 304142 286378 304226 286614
rect 304462 286378 321906 286614
rect 322142 286378 322226 286614
rect 322462 286378 339906 286614
rect 340142 286378 340226 286614
rect 340462 286378 357906 286614
rect 358142 286378 358226 286614
rect 358462 286378 375906 286614
rect 376142 286378 376226 286614
rect 376462 286378 393906 286614
rect 394142 286378 394226 286614
rect 394462 286378 411906 286614
rect 412142 286378 412226 286614
rect 412462 286378 429906 286614
rect 430142 286378 430226 286614
rect 430462 286378 447906 286614
rect 448142 286378 448226 286614
rect 448462 286378 465906 286614
rect 466142 286378 466226 286614
rect 466462 286378 483906 286614
rect 484142 286378 484226 286614
rect 484462 286378 501906 286614
rect 502142 286378 502226 286614
rect 502462 286378 519906 286614
rect 520142 286378 520226 286614
rect 520462 286378 537906 286614
rect 538142 286378 538226 286614
rect 538462 286378 547884 286614
rect 548120 286378 548204 286614
rect 548440 286378 548472 286614
rect -4476 286294 548472 286378
rect -4476 286058 -4444 286294
rect -4208 286058 -4124 286294
rect -3888 286058 15906 286294
rect 16142 286058 16226 286294
rect 16462 286058 33906 286294
rect 34142 286058 34226 286294
rect 34462 286058 51906 286294
rect 52142 286058 52226 286294
rect 52462 286058 69906 286294
rect 70142 286058 70226 286294
rect 70462 286058 87906 286294
rect 88142 286058 88226 286294
rect 88462 286058 105906 286294
rect 106142 286058 106226 286294
rect 106462 286058 123906 286294
rect 124142 286058 124226 286294
rect 124462 286058 141906 286294
rect 142142 286058 142226 286294
rect 142462 286058 159906 286294
rect 160142 286058 160226 286294
rect 160462 286058 177906 286294
rect 178142 286058 178226 286294
rect 178462 286058 195906 286294
rect 196142 286058 196226 286294
rect 196462 286058 213906 286294
rect 214142 286058 214226 286294
rect 214462 286058 231906 286294
rect 232142 286058 232226 286294
rect 232462 286058 249906 286294
rect 250142 286058 250226 286294
rect 250462 286058 267906 286294
rect 268142 286058 268226 286294
rect 268462 286058 285906 286294
rect 286142 286058 286226 286294
rect 286462 286058 303906 286294
rect 304142 286058 304226 286294
rect 304462 286058 321906 286294
rect 322142 286058 322226 286294
rect 322462 286058 339906 286294
rect 340142 286058 340226 286294
rect 340462 286058 357906 286294
rect 358142 286058 358226 286294
rect 358462 286058 375906 286294
rect 376142 286058 376226 286294
rect 376462 286058 393906 286294
rect 394142 286058 394226 286294
rect 394462 286058 411906 286294
rect 412142 286058 412226 286294
rect 412462 286058 429906 286294
rect 430142 286058 430226 286294
rect 430462 286058 447906 286294
rect 448142 286058 448226 286294
rect 448462 286058 465906 286294
rect 466142 286058 466226 286294
rect 466462 286058 483906 286294
rect 484142 286058 484226 286294
rect 484462 286058 501906 286294
rect 502142 286058 502226 286294
rect 502462 286058 519906 286294
rect 520142 286058 520226 286294
rect 520462 286058 537906 286294
rect 538142 286058 538226 286294
rect 538462 286058 547884 286294
rect 548120 286058 548204 286294
rect 548440 286058 548472 286294
rect -4476 286026 548472 286058
rect -4476 282894 548472 282926
rect -4476 282658 -3484 282894
rect -3248 282658 -3164 282894
rect -2928 282658 12186 282894
rect 12422 282658 12506 282894
rect 12742 282658 30186 282894
rect 30422 282658 30506 282894
rect 30742 282658 48186 282894
rect 48422 282658 48506 282894
rect 48742 282658 66186 282894
rect 66422 282658 66506 282894
rect 66742 282658 84186 282894
rect 84422 282658 84506 282894
rect 84742 282658 102186 282894
rect 102422 282658 102506 282894
rect 102742 282658 120186 282894
rect 120422 282658 120506 282894
rect 120742 282658 138186 282894
rect 138422 282658 138506 282894
rect 138742 282658 156186 282894
rect 156422 282658 156506 282894
rect 156742 282658 174186 282894
rect 174422 282658 174506 282894
rect 174742 282658 192186 282894
rect 192422 282658 192506 282894
rect 192742 282658 210186 282894
rect 210422 282658 210506 282894
rect 210742 282658 228186 282894
rect 228422 282658 228506 282894
rect 228742 282658 246186 282894
rect 246422 282658 246506 282894
rect 246742 282658 264186 282894
rect 264422 282658 264506 282894
rect 264742 282658 282186 282894
rect 282422 282658 282506 282894
rect 282742 282658 300186 282894
rect 300422 282658 300506 282894
rect 300742 282658 318186 282894
rect 318422 282658 318506 282894
rect 318742 282658 336186 282894
rect 336422 282658 336506 282894
rect 336742 282658 354186 282894
rect 354422 282658 354506 282894
rect 354742 282658 372186 282894
rect 372422 282658 372506 282894
rect 372742 282658 390186 282894
rect 390422 282658 390506 282894
rect 390742 282658 408186 282894
rect 408422 282658 408506 282894
rect 408742 282658 426186 282894
rect 426422 282658 426506 282894
rect 426742 282658 444186 282894
rect 444422 282658 444506 282894
rect 444742 282658 462186 282894
rect 462422 282658 462506 282894
rect 462742 282658 480186 282894
rect 480422 282658 480506 282894
rect 480742 282658 498186 282894
rect 498422 282658 498506 282894
rect 498742 282658 516186 282894
rect 516422 282658 516506 282894
rect 516742 282658 534186 282894
rect 534422 282658 534506 282894
rect 534742 282658 546924 282894
rect 547160 282658 547244 282894
rect 547480 282658 548472 282894
rect -4476 282574 548472 282658
rect -4476 282338 -3484 282574
rect -3248 282338 -3164 282574
rect -2928 282338 12186 282574
rect 12422 282338 12506 282574
rect 12742 282338 30186 282574
rect 30422 282338 30506 282574
rect 30742 282338 48186 282574
rect 48422 282338 48506 282574
rect 48742 282338 66186 282574
rect 66422 282338 66506 282574
rect 66742 282338 84186 282574
rect 84422 282338 84506 282574
rect 84742 282338 102186 282574
rect 102422 282338 102506 282574
rect 102742 282338 120186 282574
rect 120422 282338 120506 282574
rect 120742 282338 138186 282574
rect 138422 282338 138506 282574
rect 138742 282338 156186 282574
rect 156422 282338 156506 282574
rect 156742 282338 174186 282574
rect 174422 282338 174506 282574
rect 174742 282338 192186 282574
rect 192422 282338 192506 282574
rect 192742 282338 210186 282574
rect 210422 282338 210506 282574
rect 210742 282338 228186 282574
rect 228422 282338 228506 282574
rect 228742 282338 246186 282574
rect 246422 282338 246506 282574
rect 246742 282338 264186 282574
rect 264422 282338 264506 282574
rect 264742 282338 282186 282574
rect 282422 282338 282506 282574
rect 282742 282338 300186 282574
rect 300422 282338 300506 282574
rect 300742 282338 318186 282574
rect 318422 282338 318506 282574
rect 318742 282338 336186 282574
rect 336422 282338 336506 282574
rect 336742 282338 354186 282574
rect 354422 282338 354506 282574
rect 354742 282338 372186 282574
rect 372422 282338 372506 282574
rect 372742 282338 390186 282574
rect 390422 282338 390506 282574
rect 390742 282338 408186 282574
rect 408422 282338 408506 282574
rect 408742 282338 426186 282574
rect 426422 282338 426506 282574
rect 426742 282338 444186 282574
rect 444422 282338 444506 282574
rect 444742 282338 462186 282574
rect 462422 282338 462506 282574
rect 462742 282338 480186 282574
rect 480422 282338 480506 282574
rect 480742 282338 498186 282574
rect 498422 282338 498506 282574
rect 498742 282338 516186 282574
rect 516422 282338 516506 282574
rect 516742 282338 534186 282574
rect 534422 282338 534506 282574
rect 534742 282338 546924 282574
rect 547160 282338 547244 282574
rect 547480 282338 548472 282574
rect -4476 282306 548472 282338
rect -4476 279174 548472 279206
rect -4476 278938 -2524 279174
rect -2288 278938 -2204 279174
rect -1968 278938 8466 279174
rect 8702 278938 8786 279174
rect 9022 278938 26466 279174
rect 26702 278938 26786 279174
rect 27022 278938 44466 279174
rect 44702 278938 44786 279174
rect 45022 278938 62466 279174
rect 62702 278938 62786 279174
rect 63022 278938 80466 279174
rect 80702 278938 80786 279174
rect 81022 278938 98466 279174
rect 98702 278938 98786 279174
rect 99022 278938 116466 279174
rect 116702 278938 116786 279174
rect 117022 278938 134466 279174
rect 134702 278938 134786 279174
rect 135022 278938 152466 279174
rect 152702 278938 152786 279174
rect 153022 278938 170466 279174
rect 170702 278938 170786 279174
rect 171022 278938 188466 279174
rect 188702 278938 188786 279174
rect 189022 278938 206466 279174
rect 206702 278938 206786 279174
rect 207022 278938 224466 279174
rect 224702 278938 224786 279174
rect 225022 278938 242466 279174
rect 242702 278938 242786 279174
rect 243022 278938 260466 279174
rect 260702 278938 260786 279174
rect 261022 278938 278466 279174
rect 278702 278938 278786 279174
rect 279022 278938 296466 279174
rect 296702 278938 296786 279174
rect 297022 278938 314466 279174
rect 314702 278938 314786 279174
rect 315022 278938 332466 279174
rect 332702 278938 332786 279174
rect 333022 278938 350466 279174
rect 350702 278938 350786 279174
rect 351022 278938 368466 279174
rect 368702 278938 368786 279174
rect 369022 278938 386466 279174
rect 386702 278938 386786 279174
rect 387022 278938 404466 279174
rect 404702 278938 404786 279174
rect 405022 278938 422466 279174
rect 422702 278938 422786 279174
rect 423022 278938 440466 279174
rect 440702 278938 440786 279174
rect 441022 278938 458466 279174
rect 458702 278938 458786 279174
rect 459022 278938 476466 279174
rect 476702 278938 476786 279174
rect 477022 278938 494466 279174
rect 494702 278938 494786 279174
rect 495022 278938 512466 279174
rect 512702 278938 512786 279174
rect 513022 278938 530466 279174
rect 530702 278938 530786 279174
rect 531022 278938 545964 279174
rect 546200 278938 546284 279174
rect 546520 278938 548472 279174
rect -4476 278854 548472 278938
rect -4476 278618 -2524 278854
rect -2288 278618 -2204 278854
rect -1968 278618 8466 278854
rect 8702 278618 8786 278854
rect 9022 278618 26466 278854
rect 26702 278618 26786 278854
rect 27022 278618 44466 278854
rect 44702 278618 44786 278854
rect 45022 278618 62466 278854
rect 62702 278618 62786 278854
rect 63022 278618 80466 278854
rect 80702 278618 80786 278854
rect 81022 278618 98466 278854
rect 98702 278618 98786 278854
rect 99022 278618 116466 278854
rect 116702 278618 116786 278854
rect 117022 278618 134466 278854
rect 134702 278618 134786 278854
rect 135022 278618 152466 278854
rect 152702 278618 152786 278854
rect 153022 278618 170466 278854
rect 170702 278618 170786 278854
rect 171022 278618 188466 278854
rect 188702 278618 188786 278854
rect 189022 278618 206466 278854
rect 206702 278618 206786 278854
rect 207022 278618 224466 278854
rect 224702 278618 224786 278854
rect 225022 278618 242466 278854
rect 242702 278618 242786 278854
rect 243022 278618 260466 278854
rect 260702 278618 260786 278854
rect 261022 278618 278466 278854
rect 278702 278618 278786 278854
rect 279022 278618 296466 278854
rect 296702 278618 296786 278854
rect 297022 278618 314466 278854
rect 314702 278618 314786 278854
rect 315022 278618 332466 278854
rect 332702 278618 332786 278854
rect 333022 278618 350466 278854
rect 350702 278618 350786 278854
rect 351022 278618 368466 278854
rect 368702 278618 368786 278854
rect 369022 278618 386466 278854
rect 386702 278618 386786 278854
rect 387022 278618 404466 278854
rect 404702 278618 404786 278854
rect 405022 278618 422466 278854
rect 422702 278618 422786 278854
rect 423022 278618 440466 278854
rect 440702 278618 440786 278854
rect 441022 278618 458466 278854
rect 458702 278618 458786 278854
rect 459022 278618 476466 278854
rect 476702 278618 476786 278854
rect 477022 278618 494466 278854
rect 494702 278618 494786 278854
rect 495022 278618 512466 278854
rect 512702 278618 512786 278854
rect 513022 278618 530466 278854
rect 530702 278618 530786 278854
rect 531022 278618 545964 278854
rect 546200 278618 546284 278854
rect 546520 278618 548472 278854
rect -4476 278586 548472 278618
rect -4476 275454 548472 275486
rect -4476 275218 -1564 275454
rect -1328 275218 -1244 275454
rect -1008 275218 4746 275454
rect 4982 275218 5066 275454
rect 5302 275218 22746 275454
rect 22982 275218 23066 275454
rect 23302 275218 40746 275454
rect 40982 275218 41066 275454
rect 41302 275218 58746 275454
rect 58982 275218 59066 275454
rect 59302 275218 76746 275454
rect 76982 275218 77066 275454
rect 77302 275218 94746 275454
rect 94982 275218 95066 275454
rect 95302 275218 112746 275454
rect 112982 275218 113066 275454
rect 113302 275218 130746 275454
rect 130982 275218 131066 275454
rect 131302 275218 148746 275454
rect 148982 275218 149066 275454
rect 149302 275218 166746 275454
rect 166982 275218 167066 275454
rect 167302 275218 184746 275454
rect 184982 275218 185066 275454
rect 185302 275218 202746 275454
rect 202982 275218 203066 275454
rect 203302 275218 220746 275454
rect 220982 275218 221066 275454
rect 221302 275218 238746 275454
rect 238982 275218 239066 275454
rect 239302 275218 256746 275454
rect 256982 275218 257066 275454
rect 257302 275218 274746 275454
rect 274982 275218 275066 275454
rect 275302 275218 292746 275454
rect 292982 275218 293066 275454
rect 293302 275218 310746 275454
rect 310982 275218 311066 275454
rect 311302 275218 328746 275454
rect 328982 275218 329066 275454
rect 329302 275218 346746 275454
rect 346982 275218 347066 275454
rect 347302 275218 364746 275454
rect 364982 275218 365066 275454
rect 365302 275218 382746 275454
rect 382982 275218 383066 275454
rect 383302 275218 400746 275454
rect 400982 275218 401066 275454
rect 401302 275218 418746 275454
rect 418982 275218 419066 275454
rect 419302 275218 436746 275454
rect 436982 275218 437066 275454
rect 437302 275218 454746 275454
rect 454982 275218 455066 275454
rect 455302 275218 472746 275454
rect 472982 275218 473066 275454
rect 473302 275218 490746 275454
rect 490982 275218 491066 275454
rect 491302 275218 508746 275454
rect 508982 275218 509066 275454
rect 509302 275218 526746 275454
rect 526982 275218 527066 275454
rect 527302 275218 545004 275454
rect 545240 275218 545324 275454
rect 545560 275218 548472 275454
rect -4476 275134 548472 275218
rect -4476 274898 -1564 275134
rect -1328 274898 -1244 275134
rect -1008 274898 4746 275134
rect 4982 274898 5066 275134
rect 5302 274898 22746 275134
rect 22982 274898 23066 275134
rect 23302 274898 40746 275134
rect 40982 274898 41066 275134
rect 41302 274898 58746 275134
rect 58982 274898 59066 275134
rect 59302 274898 76746 275134
rect 76982 274898 77066 275134
rect 77302 274898 94746 275134
rect 94982 274898 95066 275134
rect 95302 274898 112746 275134
rect 112982 274898 113066 275134
rect 113302 274898 130746 275134
rect 130982 274898 131066 275134
rect 131302 274898 148746 275134
rect 148982 274898 149066 275134
rect 149302 274898 166746 275134
rect 166982 274898 167066 275134
rect 167302 274898 184746 275134
rect 184982 274898 185066 275134
rect 185302 274898 202746 275134
rect 202982 274898 203066 275134
rect 203302 274898 220746 275134
rect 220982 274898 221066 275134
rect 221302 274898 238746 275134
rect 238982 274898 239066 275134
rect 239302 274898 256746 275134
rect 256982 274898 257066 275134
rect 257302 274898 274746 275134
rect 274982 274898 275066 275134
rect 275302 274898 292746 275134
rect 292982 274898 293066 275134
rect 293302 274898 310746 275134
rect 310982 274898 311066 275134
rect 311302 274898 328746 275134
rect 328982 274898 329066 275134
rect 329302 274898 346746 275134
rect 346982 274898 347066 275134
rect 347302 274898 364746 275134
rect 364982 274898 365066 275134
rect 365302 274898 382746 275134
rect 382982 274898 383066 275134
rect 383302 274898 400746 275134
rect 400982 274898 401066 275134
rect 401302 274898 418746 275134
rect 418982 274898 419066 275134
rect 419302 274898 436746 275134
rect 436982 274898 437066 275134
rect 437302 274898 454746 275134
rect 454982 274898 455066 275134
rect 455302 274898 472746 275134
rect 472982 274898 473066 275134
rect 473302 274898 490746 275134
rect 490982 274898 491066 275134
rect 491302 274898 508746 275134
rect 508982 274898 509066 275134
rect 509302 274898 526746 275134
rect 526982 274898 527066 275134
rect 527302 274898 545004 275134
rect 545240 274898 545324 275134
rect 545560 274898 548472 275134
rect -4476 274866 548472 274898
rect -4476 268614 548472 268646
rect -4476 268378 -4444 268614
rect -4208 268378 -4124 268614
rect -3888 268378 15906 268614
rect 16142 268378 16226 268614
rect 16462 268378 33906 268614
rect 34142 268378 34226 268614
rect 34462 268378 51906 268614
rect 52142 268378 52226 268614
rect 52462 268378 69906 268614
rect 70142 268378 70226 268614
rect 70462 268378 87906 268614
rect 88142 268378 88226 268614
rect 88462 268378 105906 268614
rect 106142 268378 106226 268614
rect 106462 268378 123906 268614
rect 124142 268378 124226 268614
rect 124462 268378 141906 268614
rect 142142 268378 142226 268614
rect 142462 268378 159906 268614
rect 160142 268378 160226 268614
rect 160462 268378 177906 268614
rect 178142 268378 178226 268614
rect 178462 268378 195906 268614
rect 196142 268378 196226 268614
rect 196462 268378 213906 268614
rect 214142 268378 214226 268614
rect 214462 268378 231906 268614
rect 232142 268378 232226 268614
rect 232462 268378 249906 268614
rect 250142 268378 250226 268614
rect 250462 268378 267906 268614
rect 268142 268378 268226 268614
rect 268462 268378 285906 268614
rect 286142 268378 286226 268614
rect 286462 268378 303906 268614
rect 304142 268378 304226 268614
rect 304462 268378 321906 268614
rect 322142 268378 322226 268614
rect 322462 268378 339906 268614
rect 340142 268378 340226 268614
rect 340462 268378 357906 268614
rect 358142 268378 358226 268614
rect 358462 268378 375906 268614
rect 376142 268378 376226 268614
rect 376462 268378 393906 268614
rect 394142 268378 394226 268614
rect 394462 268378 411906 268614
rect 412142 268378 412226 268614
rect 412462 268378 429906 268614
rect 430142 268378 430226 268614
rect 430462 268378 447906 268614
rect 448142 268378 448226 268614
rect 448462 268378 465906 268614
rect 466142 268378 466226 268614
rect 466462 268378 483906 268614
rect 484142 268378 484226 268614
rect 484462 268378 501906 268614
rect 502142 268378 502226 268614
rect 502462 268378 519906 268614
rect 520142 268378 520226 268614
rect 520462 268378 537906 268614
rect 538142 268378 538226 268614
rect 538462 268378 547884 268614
rect 548120 268378 548204 268614
rect 548440 268378 548472 268614
rect -4476 268294 548472 268378
rect -4476 268058 -4444 268294
rect -4208 268058 -4124 268294
rect -3888 268058 15906 268294
rect 16142 268058 16226 268294
rect 16462 268058 33906 268294
rect 34142 268058 34226 268294
rect 34462 268058 51906 268294
rect 52142 268058 52226 268294
rect 52462 268058 69906 268294
rect 70142 268058 70226 268294
rect 70462 268058 87906 268294
rect 88142 268058 88226 268294
rect 88462 268058 105906 268294
rect 106142 268058 106226 268294
rect 106462 268058 123906 268294
rect 124142 268058 124226 268294
rect 124462 268058 141906 268294
rect 142142 268058 142226 268294
rect 142462 268058 159906 268294
rect 160142 268058 160226 268294
rect 160462 268058 177906 268294
rect 178142 268058 178226 268294
rect 178462 268058 195906 268294
rect 196142 268058 196226 268294
rect 196462 268058 213906 268294
rect 214142 268058 214226 268294
rect 214462 268058 231906 268294
rect 232142 268058 232226 268294
rect 232462 268058 249906 268294
rect 250142 268058 250226 268294
rect 250462 268058 267906 268294
rect 268142 268058 268226 268294
rect 268462 268058 285906 268294
rect 286142 268058 286226 268294
rect 286462 268058 303906 268294
rect 304142 268058 304226 268294
rect 304462 268058 321906 268294
rect 322142 268058 322226 268294
rect 322462 268058 339906 268294
rect 340142 268058 340226 268294
rect 340462 268058 357906 268294
rect 358142 268058 358226 268294
rect 358462 268058 375906 268294
rect 376142 268058 376226 268294
rect 376462 268058 393906 268294
rect 394142 268058 394226 268294
rect 394462 268058 411906 268294
rect 412142 268058 412226 268294
rect 412462 268058 429906 268294
rect 430142 268058 430226 268294
rect 430462 268058 447906 268294
rect 448142 268058 448226 268294
rect 448462 268058 465906 268294
rect 466142 268058 466226 268294
rect 466462 268058 483906 268294
rect 484142 268058 484226 268294
rect 484462 268058 501906 268294
rect 502142 268058 502226 268294
rect 502462 268058 519906 268294
rect 520142 268058 520226 268294
rect 520462 268058 537906 268294
rect 538142 268058 538226 268294
rect 538462 268058 547884 268294
rect 548120 268058 548204 268294
rect 548440 268058 548472 268294
rect -4476 268026 548472 268058
rect -4476 264894 548472 264926
rect -4476 264658 -3484 264894
rect -3248 264658 -3164 264894
rect -2928 264658 12186 264894
rect 12422 264658 12506 264894
rect 12742 264658 30186 264894
rect 30422 264658 30506 264894
rect 30742 264658 48186 264894
rect 48422 264658 48506 264894
rect 48742 264658 66186 264894
rect 66422 264658 66506 264894
rect 66742 264658 84186 264894
rect 84422 264658 84506 264894
rect 84742 264658 102186 264894
rect 102422 264658 102506 264894
rect 102742 264658 120186 264894
rect 120422 264658 120506 264894
rect 120742 264658 138186 264894
rect 138422 264658 138506 264894
rect 138742 264658 156186 264894
rect 156422 264658 156506 264894
rect 156742 264658 174186 264894
rect 174422 264658 174506 264894
rect 174742 264658 192186 264894
rect 192422 264658 192506 264894
rect 192742 264658 210186 264894
rect 210422 264658 210506 264894
rect 210742 264658 228186 264894
rect 228422 264658 228506 264894
rect 228742 264658 246186 264894
rect 246422 264658 246506 264894
rect 246742 264658 264186 264894
rect 264422 264658 264506 264894
rect 264742 264658 282186 264894
rect 282422 264658 282506 264894
rect 282742 264658 300186 264894
rect 300422 264658 300506 264894
rect 300742 264658 318186 264894
rect 318422 264658 318506 264894
rect 318742 264658 336186 264894
rect 336422 264658 336506 264894
rect 336742 264658 354186 264894
rect 354422 264658 354506 264894
rect 354742 264658 372186 264894
rect 372422 264658 372506 264894
rect 372742 264658 390186 264894
rect 390422 264658 390506 264894
rect 390742 264658 408186 264894
rect 408422 264658 408506 264894
rect 408742 264658 426186 264894
rect 426422 264658 426506 264894
rect 426742 264658 444186 264894
rect 444422 264658 444506 264894
rect 444742 264658 462186 264894
rect 462422 264658 462506 264894
rect 462742 264658 480186 264894
rect 480422 264658 480506 264894
rect 480742 264658 498186 264894
rect 498422 264658 498506 264894
rect 498742 264658 516186 264894
rect 516422 264658 516506 264894
rect 516742 264658 534186 264894
rect 534422 264658 534506 264894
rect 534742 264658 546924 264894
rect 547160 264658 547244 264894
rect 547480 264658 548472 264894
rect -4476 264574 548472 264658
rect -4476 264338 -3484 264574
rect -3248 264338 -3164 264574
rect -2928 264338 12186 264574
rect 12422 264338 12506 264574
rect 12742 264338 30186 264574
rect 30422 264338 30506 264574
rect 30742 264338 48186 264574
rect 48422 264338 48506 264574
rect 48742 264338 66186 264574
rect 66422 264338 66506 264574
rect 66742 264338 84186 264574
rect 84422 264338 84506 264574
rect 84742 264338 102186 264574
rect 102422 264338 102506 264574
rect 102742 264338 120186 264574
rect 120422 264338 120506 264574
rect 120742 264338 138186 264574
rect 138422 264338 138506 264574
rect 138742 264338 156186 264574
rect 156422 264338 156506 264574
rect 156742 264338 174186 264574
rect 174422 264338 174506 264574
rect 174742 264338 192186 264574
rect 192422 264338 192506 264574
rect 192742 264338 210186 264574
rect 210422 264338 210506 264574
rect 210742 264338 228186 264574
rect 228422 264338 228506 264574
rect 228742 264338 246186 264574
rect 246422 264338 246506 264574
rect 246742 264338 264186 264574
rect 264422 264338 264506 264574
rect 264742 264338 282186 264574
rect 282422 264338 282506 264574
rect 282742 264338 300186 264574
rect 300422 264338 300506 264574
rect 300742 264338 318186 264574
rect 318422 264338 318506 264574
rect 318742 264338 336186 264574
rect 336422 264338 336506 264574
rect 336742 264338 354186 264574
rect 354422 264338 354506 264574
rect 354742 264338 372186 264574
rect 372422 264338 372506 264574
rect 372742 264338 390186 264574
rect 390422 264338 390506 264574
rect 390742 264338 408186 264574
rect 408422 264338 408506 264574
rect 408742 264338 426186 264574
rect 426422 264338 426506 264574
rect 426742 264338 444186 264574
rect 444422 264338 444506 264574
rect 444742 264338 462186 264574
rect 462422 264338 462506 264574
rect 462742 264338 480186 264574
rect 480422 264338 480506 264574
rect 480742 264338 498186 264574
rect 498422 264338 498506 264574
rect 498742 264338 516186 264574
rect 516422 264338 516506 264574
rect 516742 264338 534186 264574
rect 534422 264338 534506 264574
rect 534742 264338 546924 264574
rect 547160 264338 547244 264574
rect 547480 264338 548472 264574
rect -4476 264306 548472 264338
rect -4476 261174 548472 261206
rect -4476 260938 -2524 261174
rect -2288 260938 -2204 261174
rect -1968 260938 8466 261174
rect 8702 260938 8786 261174
rect 9022 260938 26466 261174
rect 26702 260938 26786 261174
rect 27022 260938 44466 261174
rect 44702 260938 44786 261174
rect 45022 260938 62466 261174
rect 62702 260938 62786 261174
rect 63022 260938 80466 261174
rect 80702 260938 80786 261174
rect 81022 260938 98466 261174
rect 98702 260938 98786 261174
rect 99022 260938 116466 261174
rect 116702 260938 116786 261174
rect 117022 260938 134466 261174
rect 134702 260938 134786 261174
rect 135022 260938 152466 261174
rect 152702 260938 152786 261174
rect 153022 260938 170466 261174
rect 170702 260938 170786 261174
rect 171022 260938 188466 261174
rect 188702 260938 188786 261174
rect 189022 260938 206466 261174
rect 206702 260938 206786 261174
rect 207022 260938 224466 261174
rect 224702 260938 224786 261174
rect 225022 260938 242466 261174
rect 242702 260938 242786 261174
rect 243022 260938 260466 261174
rect 260702 260938 260786 261174
rect 261022 260938 278466 261174
rect 278702 260938 278786 261174
rect 279022 260938 296466 261174
rect 296702 260938 296786 261174
rect 297022 260938 314466 261174
rect 314702 260938 314786 261174
rect 315022 260938 332466 261174
rect 332702 260938 332786 261174
rect 333022 260938 350466 261174
rect 350702 260938 350786 261174
rect 351022 260938 368466 261174
rect 368702 260938 368786 261174
rect 369022 260938 386466 261174
rect 386702 260938 386786 261174
rect 387022 260938 404466 261174
rect 404702 260938 404786 261174
rect 405022 260938 422466 261174
rect 422702 260938 422786 261174
rect 423022 260938 440466 261174
rect 440702 260938 440786 261174
rect 441022 260938 458466 261174
rect 458702 260938 458786 261174
rect 459022 260938 476466 261174
rect 476702 260938 476786 261174
rect 477022 260938 494466 261174
rect 494702 260938 494786 261174
rect 495022 260938 512466 261174
rect 512702 260938 512786 261174
rect 513022 260938 530466 261174
rect 530702 260938 530786 261174
rect 531022 260938 545964 261174
rect 546200 260938 546284 261174
rect 546520 260938 548472 261174
rect -4476 260854 548472 260938
rect -4476 260618 -2524 260854
rect -2288 260618 -2204 260854
rect -1968 260618 8466 260854
rect 8702 260618 8786 260854
rect 9022 260618 26466 260854
rect 26702 260618 26786 260854
rect 27022 260618 44466 260854
rect 44702 260618 44786 260854
rect 45022 260618 62466 260854
rect 62702 260618 62786 260854
rect 63022 260618 80466 260854
rect 80702 260618 80786 260854
rect 81022 260618 98466 260854
rect 98702 260618 98786 260854
rect 99022 260618 116466 260854
rect 116702 260618 116786 260854
rect 117022 260618 134466 260854
rect 134702 260618 134786 260854
rect 135022 260618 152466 260854
rect 152702 260618 152786 260854
rect 153022 260618 170466 260854
rect 170702 260618 170786 260854
rect 171022 260618 188466 260854
rect 188702 260618 188786 260854
rect 189022 260618 206466 260854
rect 206702 260618 206786 260854
rect 207022 260618 224466 260854
rect 224702 260618 224786 260854
rect 225022 260618 242466 260854
rect 242702 260618 242786 260854
rect 243022 260618 260466 260854
rect 260702 260618 260786 260854
rect 261022 260618 278466 260854
rect 278702 260618 278786 260854
rect 279022 260618 296466 260854
rect 296702 260618 296786 260854
rect 297022 260618 314466 260854
rect 314702 260618 314786 260854
rect 315022 260618 332466 260854
rect 332702 260618 332786 260854
rect 333022 260618 350466 260854
rect 350702 260618 350786 260854
rect 351022 260618 368466 260854
rect 368702 260618 368786 260854
rect 369022 260618 386466 260854
rect 386702 260618 386786 260854
rect 387022 260618 404466 260854
rect 404702 260618 404786 260854
rect 405022 260618 422466 260854
rect 422702 260618 422786 260854
rect 423022 260618 440466 260854
rect 440702 260618 440786 260854
rect 441022 260618 458466 260854
rect 458702 260618 458786 260854
rect 459022 260618 476466 260854
rect 476702 260618 476786 260854
rect 477022 260618 494466 260854
rect 494702 260618 494786 260854
rect 495022 260618 512466 260854
rect 512702 260618 512786 260854
rect 513022 260618 530466 260854
rect 530702 260618 530786 260854
rect 531022 260618 545964 260854
rect 546200 260618 546284 260854
rect 546520 260618 548472 260854
rect -4476 260586 548472 260618
rect -4476 257454 548472 257486
rect -4476 257218 -1564 257454
rect -1328 257218 -1244 257454
rect -1008 257218 4746 257454
rect 4982 257218 5066 257454
rect 5302 257218 22746 257454
rect 22982 257218 23066 257454
rect 23302 257218 40746 257454
rect 40982 257218 41066 257454
rect 41302 257218 58746 257454
rect 58982 257218 59066 257454
rect 59302 257218 76746 257454
rect 76982 257218 77066 257454
rect 77302 257218 94746 257454
rect 94982 257218 95066 257454
rect 95302 257218 112746 257454
rect 112982 257218 113066 257454
rect 113302 257218 130746 257454
rect 130982 257218 131066 257454
rect 131302 257218 148746 257454
rect 148982 257218 149066 257454
rect 149302 257218 166746 257454
rect 166982 257218 167066 257454
rect 167302 257218 184746 257454
rect 184982 257218 185066 257454
rect 185302 257218 202746 257454
rect 202982 257218 203066 257454
rect 203302 257218 220746 257454
rect 220982 257218 221066 257454
rect 221302 257218 238746 257454
rect 238982 257218 239066 257454
rect 239302 257218 256746 257454
rect 256982 257218 257066 257454
rect 257302 257218 274746 257454
rect 274982 257218 275066 257454
rect 275302 257218 292746 257454
rect 292982 257218 293066 257454
rect 293302 257218 310746 257454
rect 310982 257218 311066 257454
rect 311302 257218 328746 257454
rect 328982 257218 329066 257454
rect 329302 257218 346746 257454
rect 346982 257218 347066 257454
rect 347302 257218 364746 257454
rect 364982 257218 365066 257454
rect 365302 257218 382746 257454
rect 382982 257218 383066 257454
rect 383302 257218 400746 257454
rect 400982 257218 401066 257454
rect 401302 257218 418746 257454
rect 418982 257218 419066 257454
rect 419302 257218 436746 257454
rect 436982 257218 437066 257454
rect 437302 257218 454746 257454
rect 454982 257218 455066 257454
rect 455302 257218 472746 257454
rect 472982 257218 473066 257454
rect 473302 257218 490746 257454
rect 490982 257218 491066 257454
rect 491302 257218 508746 257454
rect 508982 257218 509066 257454
rect 509302 257218 526746 257454
rect 526982 257218 527066 257454
rect 527302 257218 545004 257454
rect 545240 257218 545324 257454
rect 545560 257218 548472 257454
rect -4476 257134 548472 257218
rect -4476 256898 -1564 257134
rect -1328 256898 -1244 257134
rect -1008 256898 4746 257134
rect 4982 256898 5066 257134
rect 5302 256898 22746 257134
rect 22982 256898 23066 257134
rect 23302 256898 40746 257134
rect 40982 256898 41066 257134
rect 41302 256898 58746 257134
rect 58982 256898 59066 257134
rect 59302 256898 76746 257134
rect 76982 256898 77066 257134
rect 77302 256898 94746 257134
rect 94982 256898 95066 257134
rect 95302 256898 112746 257134
rect 112982 256898 113066 257134
rect 113302 256898 130746 257134
rect 130982 256898 131066 257134
rect 131302 256898 148746 257134
rect 148982 256898 149066 257134
rect 149302 256898 166746 257134
rect 166982 256898 167066 257134
rect 167302 256898 184746 257134
rect 184982 256898 185066 257134
rect 185302 256898 202746 257134
rect 202982 256898 203066 257134
rect 203302 256898 220746 257134
rect 220982 256898 221066 257134
rect 221302 256898 238746 257134
rect 238982 256898 239066 257134
rect 239302 256898 256746 257134
rect 256982 256898 257066 257134
rect 257302 256898 274746 257134
rect 274982 256898 275066 257134
rect 275302 256898 292746 257134
rect 292982 256898 293066 257134
rect 293302 256898 310746 257134
rect 310982 256898 311066 257134
rect 311302 256898 328746 257134
rect 328982 256898 329066 257134
rect 329302 256898 346746 257134
rect 346982 256898 347066 257134
rect 347302 256898 364746 257134
rect 364982 256898 365066 257134
rect 365302 256898 382746 257134
rect 382982 256898 383066 257134
rect 383302 256898 400746 257134
rect 400982 256898 401066 257134
rect 401302 256898 418746 257134
rect 418982 256898 419066 257134
rect 419302 256898 436746 257134
rect 436982 256898 437066 257134
rect 437302 256898 454746 257134
rect 454982 256898 455066 257134
rect 455302 256898 472746 257134
rect 472982 256898 473066 257134
rect 473302 256898 490746 257134
rect 490982 256898 491066 257134
rect 491302 256898 508746 257134
rect 508982 256898 509066 257134
rect 509302 256898 526746 257134
rect 526982 256898 527066 257134
rect 527302 256898 545004 257134
rect 545240 256898 545324 257134
rect 545560 256898 548472 257134
rect -4476 256866 548472 256898
rect -4476 250614 548472 250646
rect -4476 250378 -4444 250614
rect -4208 250378 -4124 250614
rect -3888 250378 15906 250614
rect 16142 250378 16226 250614
rect 16462 250378 33906 250614
rect 34142 250378 34226 250614
rect 34462 250378 51906 250614
rect 52142 250378 52226 250614
rect 52462 250378 69906 250614
rect 70142 250378 70226 250614
rect 70462 250378 87906 250614
rect 88142 250378 88226 250614
rect 88462 250378 105906 250614
rect 106142 250378 106226 250614
rect 106462 250378 123906 250614
rect 124142 250378 124226 250614
rect 124462 250378 141906 250614
rect 142142 250378 142226 250614
rect 142462 250378 159906 250614
rect 160142 250378 160226 250614
rect 160462 250378 177906 250614
rect 178142 250378 178226 250614
rect 178462 250378 195906 250614
rect 196142 250378 196226 250614
rect 196462 250378 213906 250614
rect 214142 250378 214226 250614
rect 214462 250378 231906 250614
rect 232142 250378 232226 250614
rect 232462 250378 249906 250614
rect 250142 250378 250226 250614
rect 250462 250378 267906 250614
rect 268142 250378 268226 250614
rect 268462 250378 285906 250614
rect 286142 250378 286226 250614
rect 286462 250378 303906 250614
rect 304142 250378 304226 250614
rect 304462 250378 321906 250614
rect 322142 250378 322226 250614
rect 322462 250378 339906 250614
rect 340142 250378 340226 250614
rect 340462 250378 357906 250614
rect 358142 250378 358226 250614
rect 358462 250378 375906 250614
rect 376142 250378 376226 250614
rect 376462 250378 393906 250614
rect 394142 250378 394226 250614
rect 394462 250378 411906 250614
rect 412142 250378 412226 250614
rect 412462 250378 429906 250614
rect 430142 250378 430226 250614
rect 430462 250378 447906 250614
rect 448142 250378 448226 250614
rect 448462 250378 465906 250614
rect 466142 250378 466226 250614
rect 466462 250378 483906 250614
rect 484142 250378 484226 250614
rect 484462 250378 501906 250614
rect 502142 250378 502226 250614
rect 502462 250378 519906 250614
rect 520142 250378 520226 250614
rect 520462 250378 537906 250614
rect 538142 250378 538226 250614
rect 538462 250378 547884 250614
rect 548120 250378 548204 250614
rect 548440 250378 548472 250614
rect -4476 250294 548472 250378
rect -4476 250058 -4444 250294
rect -4208 250058 -4124 250294
rect -3888 250058 15906 250294
rect 16142 250058 16226 250294
rect 16462 250058 33906 250294
rect 34142 250058 34226 250294
rect 34462 250058 51906 250294
rect 52142 250058 52226 250294
rect 52462 250058 69906 250294
rect 70142 250058 70226 250294
rect 70462 250058 87906 250294
rect 88142 250058 88226 250294
rect 88462 250058 105906 250294
rect 106142 250058 106226 250294
rect 106462 250058 123906 250294
rect 124142 250058 124226 250294
rect 124462 250058 141906 250294
rect 142142 250058 142226 250294
rect 142462 250058 159906 250294
rect 160142 250058 160226 250294
rect 160462 250058 177906 250294
rect 178142 250058 178226 250294
rect 178462 250058 195906 250294
rect 196142 250058 196226 250294
rect 196462 250058 213906 250294
rect 214142 250058 214226 250294
rect 214462 250058 231906 250294
rect 232142 250058 232226 250294
rect 232462 250058 249906 250294
rect 250142 250058 250226 250294
rect 250462 250058 267906 250294
rect 268142 250058 268226 250294
rect 268462 250058 285906 250294
rect 286142 250058 286226 250294
rect 286462 250058 303906 250294
rect 304142 250058 304226 250294
rect 304462 250058 321906 250294
rect 322142 250058 322226 250294
rect 322462 250058 339906 250294
rect 340142 250058 340226 250294
rect 340462 250058 357906 250294
rect 358142 250058 358226 250294
rect 358462 250058 375906 250294
rect 376142 250058 376226 250294
rect 376462 250058 393906 250294
rect 394142 250058 394226 250294
rect 394462 250058 411906 250294
rect 412142 250058 412226 250294
rect 412462 250058 429906 250294
rect 430142 250058 430226 250294
rect 430462 250058 447906 250294
rect 448142 250058 448226 250294
rect 448462 250058 465906 250294
rect 466142 250058 466226 250294
rect 466462 250058 483906 250294
rect 484142 250058 484226 250294
rect 484462 250058 501906 250294
rect 502142 250058 502226 250294
rect 502462 250058 519906 250294
rect 520142 250058 520226 250294
rect 520462 250058 537906 250294
rect 538142 250058 538226 250294
rect 538462 250058 547884 250294
rect 548120 250058 548204 250294
rect 548440 250058 548472 250294
rect -4476 250026 548472 250058
rect -4476 246894 548472 246926
rect -4476 246658 -3484 246894
rect -3248 246658 -3164 246894
rect -2928 246658 12186 246894
rect 12422 246658 12506 246894
rect 12742 246658 30186 246894
rect 30422 246658 30506 246894
rect 30742 246658 48186 246894
rect 48422 246658 48506 246894
rect 48742 246658 66186 246894
rect 66422 246658 66506 246894
rect 66742 246658 84186 246894
rect 84422 246658 84506 246894
rect 84742 246658 102186 246894
rect 102422 246658 102506 246894
rect 102742 246658 120186 246894
rect 120422 246658 120506 246894
rect 120742 246658 138186 246894
rect 138422 246658 138506 246894
rect 138742 246658 156186 246894
rect 156422 246658 156506 246894
rect 156742 246658 174186 246894
rect 174422 246658 174506 246894
rect 174742 246658 192186 246894
rect 192422 246658 192506 246894
rect 192742 246658 210186 246894
rect 210422 246658 210506 246894
rect 210742 246658 228186 246894
rect 228422 246658 228506 246894
rect 228742 246658 246186 246894
rect 246422 246658 246506 246894
rect 246742 246658 264186 246894
rect 264422 246658 264506 246894
rect 264742 246658 282186 246894
rect 282422 246658 282506 246894
rect 282742 246658 300186 246894
rect 300422 246658 300506 246894
rect 300742 246658 318186 246894
rect 318422 246658 318506 246894
rect 318742 246658 336186 246894
rect 336422 246658 336506 246894
rect 336742 246658 354186 246894
rect 354422 246658 354506 246894
rect 354742 246658 372186 246894
rect 372422 246658 372506 246894
rect 372742 246658 390186 246894
rect 390422 246658 390506 246894
rect 390742 246658 408186 246894
rect 408422 246658 408506 246894
rect 408742 246658 426186 246894
rect 426422 246658 426506 246894
rect 426742 246658 444186 246894
rect 444422 246658 444506 246894
rect 444742 246658 462186 246894
rect 462422 246658 462506 246894
rect 462742 246658 480186 246894
rect 480422 246658 480506 246894
rect 480742 246658 498186 246894
rect 498422 246658 498506 246894
rect 498742 246658 516186 246894
rect 516422 246658 516506 246894
rect 516742 246658 534186 246894
rect 534422 246658 534506 246894
rect 534742 246658 546924 246894
rect 547160 246658 547244 246894
rect 547480 246658 548472 246894
rect -4476 246574 548472 246658
rect -4476 246338 -3484 246574
rect -3248 246338 -3164 246574
rect -2928 246338 12186 246574
rect 12422 246338 12506 246574
rect 12742 246338 30186 246574
rect 30422 246338 30506 246574
rect 30742 246338 48186 246574
rect 48422 246338 48506 246574
rect 48742 246338 66186 246574
rect 66422 246338 66506 246574
rect 66742 246338 84186 246574
rect 84422 246338 84506 246574
rect 84742 246338 102186 246574
rect 102422 246338 102506 246574
rect 102742 246338 120186 246574
rect 120422 246338 120506 246574
rect 120742 246338 138186 246574
rect 138422 246338 138506 246574
rect 138742 246338 156186 246574
rect 156422 246338 156506 246574
rect 156742 246338 174186 246574
rect 174422 246338 174506 246574
rect 174742 246338 192186 246574
rect 192422 246338 192506 246574
rect 192742 246338 210186 246574
rect 210422 246338 210506 246574
rect 210742 246338 228186 246574
rect 228422 246338 228506 246574
rect 228742 246338 246186 246574
rect 246422 246338 246506 246574
rect 246742 246338 264186 246574
rect 264422 246338 264506 246574
rect 264742 246338 282186 246574
rect 282422 246338 282506 246574
rect 282742 246338 300186 246574
rect 300422 246338 300506 246574
rect 300742 246338 318186 246574
rect 318422 246338 318506 246574
rect 318742 246338 336186 246574
rect 336422 246338 336506 246574
rect 336742 246338 354186 246574
rect 354422 246338 354506 246574
rect 354742 246338 372186 246574
rect 372422 246338 372506 246574
rect 372742 246338 390186 246574
rect 390422 246338 390506 246574
rect 390742 246338 408186 246574
rect 408422 246338 408506 246574
rect 408742 246338 426186 246574
rect 426422 246338 426506 246574
rect 426742 246338 444186 246574
rect 444422 246338 444506 246574
rect 444742 246338 462186 246574
rect 462422 246338 462506 246574
rect 462742 246338 480186 246574
rect 480422 246338 480506 246574
rect 480742 246338 498186 246574
rect 498422 246338 498506 246574
rect 498742 246338 516186 246574
rect 516422 246338 516506 246574
rect 516742 246338 534186 246574
rect 534422 246338 534506 246574
rect 534742 246338 546924 246574
rect 547160 246338 547244 246574
rect 547480 246338 548472 246574
rect -4476 246306 548472 246338
rect -4476 243174 548472 243206
rect -4476 242938 -2524 243174
rect -2288 242938 -2204 243174
rect -1968 242938 8466 243174
rect 8702 242938 8786 243174
rect 9022 242938 26466 243174
rect 26702 242938 26786 243174
rect 27022 242938 44466 243174
rect 44702 242938 44786 243174
rect 45022 242938 62466 243174
rect 62702 242938 62786 243174
rect 63022 242938 80466 243174
rect 80702 242938 80786 243174
rect 81022 242938 98466 243174
rect 98702 242938 98786 243174
rect 99022 242938 116466 243174
rect 116702 242938 116786 243174
rect 117022 242938 134466 243174
rect 134702 242938 134786 243174
rect 135022 242938 152466 243174
rect 152702 242938 152786 243174
rect 153022 242938 170466 243174
rect 170702 242938 170786 243174
rect 171022 242938 188466 243174
rect 188702 242938 188786 243174
rect 189022 242938 206466 243174
rect 206702 242938 206786 243174
rect 207022 242938 224466 243174
rect 224702 242938 224786 243174
rect 225022 242938 242466 243174
rect 242702 242938 242786 243174
rect 243022 242938 260466 243174
rect 260702 242938 260786 243174
rect 261022 242938 278466 243174
rect 278702 242938 278786 243174
rect 279022 242938 296466 243174
rect 296702 242938 296786 243174
rect 297022 242938 314466 243174
rect 314702 242938 314786 243174
rect 315022 242938 332466 243174
rect 332702 242938 332786 243174
rect 333022 242938 350466 243174
rect 350702 242938 350786 243174
rect 351022 242938 368466 243174
rect 368702 242938 368786 243174
rect 369022 242938 386466 243174
rect 386702 242938 386786 243174
rect 387022 242938 404466 243174
rect 404702 242938 404786 243174
rect 405022 242938 422466 243174
rect 422702 242938 422786 243174
rect 423022 242938 440466 243174
rect 440702 242938 440786 243174
rect 441022 242938 458466 243174
rect 458702 242938 458786 243174
rect 459022 242938 476466 243174
rect 476702 242938 476786 243174
rect 477022 242938 494466 243174
rect 494702 242938 494786 243174
rect 495022 242938 512466 243174
rect 512702 242938 512786 243174
rect 513022 242938 530466 243174
rect 530702 242938 530786 243174
rect 531022 242938 545964 243174
rect 546200 242938 546284 243174
rect 546520 242938 548472 243174
rect -4476 242854 548472 242938
rect -4476 242618 -2524 242854
rect -2288 242618 -2204 242854
rect -1968 242618 8466 242854
rect 8702 242618 8786 242854
rect 9022 242618 26466 242854
rect 26702 242618 26786 242854
rect 27022 242618 44466 242854
rect 44702 242618 44786 242854
rect 45022 242618 62466 242854
rect 62702 242618 62786 242854
rect 63022 242618 80466 242854
rect 80702 242618 80786 242854
rect 81022 242618 98466 242854
rect 98702 242618 98786 242854
rect 99022 242618 116466 242854
rect 116702 242618 116786 242854
rect 117022 242618 134466 242854
rect 134702 242618 134786 242854
rect 135022 242618 152466 242854
rect 152702 242618 152786 242854
rect 153022 242618 170466 242854
rect 170702 242618 170786 242854
rect 171022 242618 188466 242854
rect 188702 242618 188786 242854
rect 189022 242618 206466 242854
rect 206702 242618 206786 242854
rect 207022 242618 224466 242854
rect 224702 242618 224786 242854
rect 225022 242618 242466 242854
rect 242702 242618 242786 242854
rect 243022 242618 260466 242854
rect 260702 242618 260786 242854
rect 261022 242618 278466 242854
rect 278702 242618 278786 242854
rect 279022 242618 296466 242854
rect 296702 242618 296786 242854
rect 297022 242618 314466 242854
rect 314702 242618 314786 242854
rect 315022 242618 332466 242854
rect 332702 242618 332786 242854
rect 333022 242618 350466 242854
rect 350702 242618 350786 242854
rect 351022 242618 368466 242854
rect 368702 242618 368786 242854
rect 369022 242618 386466 242854
rect 386702 242618 386786 242854
rect 387022 242618 404466 242854
rect 404702 242618 404786 242854
rect 405022 242618 422466 242854
rect 422702 242618 422786 242854
rect 423022 242618 440466 242854
rect 440702 242618 440786 242854
rect 441022 242618 458466 242854
rect 458702 242618 458786 242854
rect 459022 242618 476466 242854
rect 476702 242618 476786 242854
rect 477022 242618 494466 242854
rect 494702 242618 494786 242854
rect 495022 242618 512466 242854
rect 512702 242618 512786 242854
rect 513022 242618 530466 242854
rect 530702 242618 530786 242854
rect 531022 242618 545964 242854
rect 546200 242618 546284 242854
rect 546520 242618 548472 242854
rect -4476 242586 548472 242618
rect -4476 239454 548472 239486
rect -4476 239218 -1564 239454
rect -1328 239218 -1244 239454
rect -1008 239218 4746 239454
rect 4982 239218 5066 239454
rect 5302 239218 22746 239454
rect 22982 239218 23066 239454
rect 23302 239218 40746 239454
rect 40982 239218 41066 239454
rect 41302 239218 58746 239454
rect 58982 239218 59066 239454
rect 59302 239218 76746 239454
rect 76982 239218 77066 239454
rect 77302 239218 94746 239454
rect 94982 239218 95066 239454
rect 95302 239218 112746 239454
rect 112982 239218 113066 239454
rect 113302 239218 130746 239454
rect 130982 239218 131066 239454
rect 131302 239218 148746 239454
rect 148982 239218 149066 239454
rect 149302 239218 166746 239454
rect 166982 239218 167066 239454
rect 167302 239218 184746 239454
rect 184982 239218 185066 239454
rect 185302 239218 202746 239454
rect 202982 239218 203066 239454
rect 203302 239218 220746 239454
rect 220982 239218 221066 239454
rect 221302 239218 238746 239454
rect 238982 239218 239066 239454
rect 239302 239218 256746 239454
rect 256982 239218 257066 239454
rect 257302 239218 274746 239454
rect 274982 239218 275066 239454
rect 275302 239218 292746 239454
rect 292982 239218 293066 239454
rect 293302 239218 310746 239454
rect 310982 239218 311066 239454
rect 311302 239218 328746 239454
rect 328982 239218 329066 239454
rect 329302 239218 346746 239454
rect 346982 239218 347066 239454
rect 347302 239218 364746 239454
rect 364982 239218 365066 239454
rect 365302 239218 382746 239454
rect 382982 239218 383066 239454
rect 383302 239218 400746 239454
rect 400982 239218 401066 239454
rect 401302 239218 418746 239454
rect 418982 239218 419066 239454
rect 419302 239218 436746 239454
rect 436982 239218 437066 239454
rect 437302 239218 454746 239454
rect 454982 239218 455066 239454
rect 455302 239218 472746 239454
rect 472982 239218 473066 239454
rect 473302 239218 490746 239454
rect 490982 239218 491066 239454
rect 491302 239218 508746 239454
rect 508982 239218 509066 239454
rect 509302 239218 526746 239454
rect 526982 239218 527066 239454
rect 527302 239218 545004 239454
rect 545240 239218 545324 239454
rect 545560 239218 548472 239454
rect -4476 239134 548472 239218
rect -4476 238898 -1564 239134
rect -1328 238898 -1244 239134
rect -1008 238898 4746 239134
rect 4982 238898 5066 239134
rect 5302 238898 22746 239134
rect 22982 238898 23066 239134
rect 23302 238898 40746 239134
rect 40982 238898 41066 239134
rect 41302 238898 58746 239134
rect 58982 238898 59066 239134
rect 59302 238898 76746 239134
rect 76982 238898 77066 239134
rect 77302 238898 94746 239134
rect 94982 238898 95066 239134
rect 95302 238898 112746 239134
rect 112982 238898 113066 239134
rect 113302 238898 130746 239134
rect 130982 238898 131066 239134
rect 131302 238898 148746 239134
rect 148982 238898 149066 239134
rect 149302 238898 166746 239134
rect 166982 238898 167066 239134
rect 167302 238898 184746 239134
rect 184982 238898 185066 239134
rect 185302 238898 202746 239134
rect 202982 238898 203066 239134
rect 203302 238898 220746 239134
rect 220982 238898 221066 239134
rect 221302 238898 238746 239134
rect 238982 238898 239066 239134
rect 239302 238898 256746 239134
rect 256982 238898 257066 239134
rect 257302 238898 274746 239134
rect 274982 238898 275066 239134
rect 275302 238898 292746 239134
rect 292982 238898 293066 239134
rect 293302 238898 310746 239134
rect 310982 238898 311066 239134
rect 311302 238898 328746 239134
rect 328982 238898 329066 239134
rect 329302 238898 346746 239134
rect 346982 238898 347066 239134
rect 347302 238898 364746 239134
rect 364982 238898 365066 239134
rect 365302 238898 382746 239134
rect 382982 238898 383066 239134
rect 383302 238898 400746 239134
rect 400982 238898 401066 239134
rect 401302 238898 418746 239134
rect 418982 238898 419066 239134
rect 419302 238898 436746 239134
rect 436982 238898 437066 239134
rect 437302 238898 454746 239134
rect 454982 238898 455066 239134
rect 455302 238898 472746 239134
rect 472982 238898 473066 239134
rect 473302 238898 490746 239134
rect 490982 238898 491066 239134
rect 491302 238898 508746 239134
rect 508982 238898 509066 239134
rect 509302 238898 526746 239134
rect 526982 238898 527066 239134
rect 527302 238898 545004 239134
rect 545240 238898 545324 239134
rect 545560 238898 548472 239134
rect -4476 238866 548472 238898
rect -4476 232614 548472 232646
rect -4476 232378 -4444 232614
rect -4208 232378 -4124 232614
rect -3888 232378 15906 232614
rect 16142 232378 16226 232614
rect 16462 232378 33906 232614
rect 34142 232378 34226 232614
rect 34462 232378 51906 232614
rect 52142 232378 52226 232614
rect 52462 232378 69906 232614
rect 70142 232378 70226 232614
rect 70462 232378 87906 232614
rect 88142 232378 88226 232614
rect 88462 232378 105906 232614
rect 106142 232378 106226 232614
rect 106462 232378 123906 232614
rect 124142 232378 124226 232614
rect 124462 232378 141906 232614
rect 142142 232378 142226 232614
rect 142462 232378 159906 232614
rect 160142 232378 160226 232614
rect 160462 232378 177906 232614
rect 178142 232378 178226 232614
rect 178462 232378 195906 232614
rect 196142 232378 196226 232614
rect 196462 232378 213906 232614
rect 214142 232378 214226 232614
rect 214462 232378 231906 232614
rect 232142 232378 232226 232614
rect 232462 232378 249906 232614
rect 250142 232378 250226 232614
rect 250462 232378 267906 232614
rect 268142 232378 268226 232614
rect 268462 232378 285906 232614
rect 286142 232378 286226 232614
rect 286462 232378 303906 232614
rect 304142 232378 304226 232614
rect 304462 232378 321906 232614
rect 322142 232378 322226 232614
rect 322462 232378 339906 232614
rect 340142 232378 340226 232614
rect 340462 232378 357906 232614
rect 358142 232378 358226 232614
rect 358462 232378 375906 232614
rect 376142 232378 376226 232614
rect 376462 232378 393906 232614
rect 394142 232378 394226 232614
rect 394462 232378 411906 232614
rect 412142 232378 412226 232614
rect 412462 232378 429906 232614
rect 430142 232378 430226 232614
rect 430462 232378 447906 232614
rect 448142 232378 448226 232614
rect 448462 232378 465906 232614
rect 466142 232378 466226 232614
rect 466462 232378 483906 232614
rect 484142 232378 484226 232614
rect 484462 232378 501906 232614
rect 502142 232378 502226 232614
rect 502462 232378 519906 232614
rect 520142 232378 520226 232614
rect 520462 232378 537906 232614
rect 538142 232378 538226 232614
rect 538462 232378 547884 232614
rect 548120 232378 548204 232614
rect 548440 232378 548472 232614
rect -4476 232294 548472 232378
rect -4476 232058 -4444 232294
rect -4208 232058 -4124 232294
rect -3888 232058 15906 232294
rect 16142 232058 16226 232294
rect 16462 232058 33906 232294
rect 34142 232058 34226 232294
rect 34462 232058 51906 232294
rect 52142 232058 52226 232294
rect 52462 232058 69906 232294
rect 70142 232058 70226 232294
rect 70462 232058 87906 232294
rect 88142 232058 88226 232294
rect 88462 232058 105906 232294
rect 106142 232058 106226 232294
rect 106462 232058 123906 232294
rect 124142 232058 124226 232294
rect 124462 232058 141906 232294
rect 142142 232058 142226 232294
rect 142462 232058 159906 232294
rect 160142 232058 160226 232294
rect 160462 232058 177906 232294
rect 178142 232058 178226 232294
rect 178462 232058 195906 232294
rect 196142 232058 196226 232294
rect 196462 232058 213906 232294
rect 214142 232058 214226 232294
rect 214462 232058 231906 232294
rect 232142 232058 232226 232294
rect 232462 232058 249906 232294
rect 250142 232058 250226 232294
rect 250462 232058 267906 232294
rect 268142 232058 268226 232294
rect 268462 232058 285906 232294
rect 286142 232058 286226 232294
rect 286462 232058 303906 232294
rect 304142 232058 304226 232294
rect 304462 232058 321906 232294
rect 322142 232058 322226 232294
rect 322462 232058 339906 232294
rect 340142 232058 340226 232294
rect 340462 232058 357906 232294
rect 358142 232058 358226 232294
rect 358462 232058 375906 232294
rect 376142 232058 376226 232294
rect 376462 232058 393906 232294
rect 394142 232058 394226 232294
rect 394462 232058 411906 232294
rect 412142 232058 412226 232294
rect 412462 232058 429906 232294
rect 430142 232058 430226 232294
rect 430462 232058 447906 232294
rect 448142 232058 448226 232294
rect 448462 232058 465906 232294
rect 466142 232058 466226 232294
rect 466462 232058 483906 232294
rect 484142 232058 484226 232294
rect 484462 232058 501906 232294
rect 502142 232058 502226 232294
rect 502462 232058 519906 232294
rect 520142 232058 520226 232294
rect 520462 232058 537906 232294
rect 538142 232058 538226 232294
rect 538462 232058 547884 232294
rect 548120 232058 548204 232294
rect 548440 232058 548472 232294
rect -4476 232026 548472 232058
rect -4476 228894 548472 228926
rect -4476 228658 -3484 228894
rect -3248 228658 -3164 228894
rect -2928 228658 12186 228894
rect 12422 228658 12506 228894
rect 12742 228658 30186 228894
rect 30422 228658 30506 228894
rect 30742 228658 48186 228894
rect 48422 228658 48506 228894
rect 48742 228658 66186 228894
rect 66422 228658 66506 228894
rect 66742 228658 84186 228894
rect 84422 228658 84506 228894
rect 84742 228658 102186 228894
rect 102422 228658 102506 228894
rect 102742 228658 120186 228894
rect 120422 228658 120506 228894
rect 120742 228658 138186 228894
rect 138422 228658 138506 228894
rect 138742 228658 156186 228894
rect 156422 228658 156506 228894
rect 156742 228658 174186 228894
rect 174422 228658 174506 228894
rect 174742 228658 192186 228894
rect 192422 228658 192506 228894
rect 192742 228658 210186 228894
rect 210422 228658 210506 228894
rect 210742 228658 228186 228894
rect 228422 228658 228506 228894
rect 228742 228658 246186 228894
rect 246422 228658 246506 228894
rect 246742 228658 264186 228894
rect 264422 228658 264506 228894
rect 264742 228658 282186 228894
rect 282422 228658 282506 228894
rect 282742 228658 300186 228894
rect 300422 228658 300506 228894
rect 300742 228658 318186 228894
rect 318422 228658 318506 228894
rect 318742 228658 336186 228894
rect 336422 228658 336506 228894
rect 336742 228658 354186 228894
rect 354422 228658 354506 228894
rect 354742 228658 372186 228894
rect 372422 228658 372506 228894
rect 372742 228658 390186 228894
rect 390422 228658 390506 228894
rect 390742 228658 408186 228894
rect 408422 228658 408506 228894
rect 408742 228658 426186 228894
rect 426422 228658 426506 228894
rect 426742 228658 444186 228894
rect 444422 228658 444506 228894
rect 444742 228658 462186 228894
rect 462422 228658 462506 228894
rect 462742 228658 480186 228894
rect 480422 228658 480506 228894
rect 480742 228658 498186 228894
rect 498422 228658 498506 228894
rect 498742 228658 516186 228894
rect 516422 228658 516506 228894
rect 516742 228658 534186 228894
rect 534422 228658 534506 228894
rect 534742 228658 546924 228894
rect 547160 228658 547244 228894
rect 547480 228658 548472 228894
rect -4476 228574 548472 228658
rect -4476 228338 -3484 228574
rect -3248 228338 -3164 228574
rect -2928 228338 12186 228574
rect 12422 228338 12506 228574
rect 12742 228338 30186 228574
rect 30422 228338 30506 228574
rect 30742 228338 48186 228574
rect 48422 228338 48506 228574
rect 48742 228338 66186 228574
rect 66422 228338 66506 228574
rect 66742 228338 84186 228574
rect 84422 228338 84506 228574
rect 84742 228338 102186 228574
rect 102422 228338 102506 228574
rect 102742 228338 120186 228574
rect 120422 228338 120506 228574
rect 120742 228338 138186 228574
rect 138422 228338 138506 228574
rect 138742 228338 156186 228574
rect 156422 228338 156506 228574
rect 156742 228338 174186 228574
rect 174422 228338 174506 228574
rect 174742 228338 192186 228574
rect 192422 228338 192506 228574
rect 192742 228338 210186 228574
rect 210422 228338 210506 228574
rect 210742 228338 228186 228574
rect 228422 228338 228506 228574
rect 228742 228338 246186 228574
rect 246422 228338 246506 228574
rect 246742 228338 264186 228574
rect 264422 228338 264506 228574
rect 264742 228338 282186 228574
rect 282422 228338 282506 228574
rect 282742 228338 300186 228574
rect 300422 228338 300506 228574
rect 300742 228338 318186 228574
rect 318422 228338 318506 228574
rect 318742 228338 336186 228574
rect 336422 228338 336506 228574
rect 336742 228338 354186 228574
rect 354422 228338 354506 228574
rect 354742 228338 372186 228574
rect 372422 228338 372506 228574
rect 372742 228338 390186 228574
rect 390422 228338 390506 228574
rect 390742 228338 408186 228574
rect 408422 228338 408506 228574
rect 408742 228338 426186 228574
rect 426422 228338 426506 228574
rect 426742 228338 444186 228574
rect 444422 228338 444506 228574
rect 444742 228338 462186 228574
rect 462422 228338 462506 228574
rect 462742 228338 480186 228574
rect 480422 228338 480506 228574
rect 480742 228338 498186 228574
rect 498422 228338 498506 228574
rect 498742 228338 516186 228574
rect 516422 228338 516506 228574
rect 516742 228338 534186 228574
rect 534422 228338 534506 228574
rect 534742 228338 546924 228574
rect 547160 228338 547244 228574
rect 547480 228338 548472 228574
rect -4476 228306 548472 228338
rect -4476 225174 548472 225206
rect -4476 224938 -2524 225174
rect -2288 224938 -2204 225174
rect -1968 224938 8466 225174
rect 8702 224938 8786 225174
rect 9022 224938 26466 225174
rect 26702 224938 26786 225174
rect 27022 224938 44466 225174
rect 44702 224938 44786 225174
rect 45022 224938 62466 225174
rect 62702 224938 62786 225174
rect 63022 224938 80466 225174
rect 80702 224938 80786 225174
rect 81022 224938 98466 225174
rect 98702 224938 98786 225174
rect 99022 224938 116466 225174
rect 116702 224938 116786 225174
rect 117022 224938 134466 225174
rect 134702 224938 134786 225174
rect 135022 224938 152466 225174
rect 152702 224938 152786 225174
rect 153022 224938 170466 225174
rect 170702 224938 170786 225174
rect 171022 224938 188466 225174
rect 188702 224938 188786 225174
rect 189022 224938 206466 225174
rect 206702 224938 206786 225174
rect 207022 224938 224466 225174
rect 224702 224938 224786 225174
rect 225022 224938 242466 225174
rect 242702 224938 242786 225174
rect 243022 224938 260466 225174
rect 260702 224938 260786 225174
rect 261022 224938 278466 225174
rect 278702 224938 278786 225174
rect 279022 224938 296466 225174
rect 296702 224938 296786 225174
rect 297022 224938 314466 225174
rect 314702 224938 314786 225174
rect 315022 224938 332466 225174
rect 332702 224938 332786 225174
rect 333022 224938 350466 225174
rect 350702 224938 350786 225174
rect 351022 224938 368466 225174
rect 368702 224938 368786 225174
rect 369022 224938 386466 225174
rect 386702 224938 386786 225174
rect 387022 224938 404466 225174
rect 404702 224938 404786 225174
rect 405022 224938 422466 225174
rect 422702 224938 422786 225174
rect 423022 224938 440466 225174
rect 440702 224938 440786 225174
rect 441022 224938 458466 225174
rect 458702 224938 458786 225174
rect 459022 224938 476466 225174
rect 476702 224938 476786 225174
rect 477022 224938 494466 225174
rect 494702 224938 494786 225174
rect 495022 224938 512466 225174
rect 512702 224938 512786 225174
rect 513022 224938 530466 225174
rect 530702 224938 530786 225174
rect 531022 224938 545964 225174
rect 546200 224938 546284 225174
rect 546520 224938 548472 225174
rect -4476 224854 548472 224938
rect -4476 224618 -2524 224854
rect -2288 224618 -2204 224854
rect -1968 224618 8466 224854
rect 8702 224618 8786 224854
rect 9022 224618 26466 224854
rect 26702 224618 26786 224854
rect 27022 224618 44466 224854
rect 44702 224618 44786 224854
rect 45022 224618 62466 224854
rect 62702 224618 62786 224854
rect 63022 224618 80466 224854
rect 80702 224618 80786 224854
rect 81022 224618 98466 224854
rect 98702 224618 98786 224854
rect 99022 224618 116466 224854
rect 116702 224618 116786 224854
rect 117022 224618 134466 224854
rect 134702 224618 134786 224854
rect 135022 224618 152466 224854
rect 152702 224618 152786 224854
rect 153022 224618 170466 224854
rect 170702 224618 170786 224854
rect 171022 224618 188466 224854
rect 188702 224618 188786 224854
rect 189022 224618 206466 224854
rect 206702 224618 206786 224854
rect 207022 224618 224466 224854
rect 224702 224618 224786 224854
rect 225022 224618 242466 224854
rect 242702 224618 242786 224854
rect 243022 224618 260466 224854
rect 260702 224618 260786 224854
rect 261022 224618 278466 224854
rect 278702 224618 278786 224854
rect 279022 224618 296466 224854
rect 296702 224618 296786 224854
rect 297022 224618 314466 224854
rect 314702 224618 314786 224854
rect 315022 224618 332466 224854
rect 332702 224618 332786 224854
rect 333022 224618 350466 224854
rect 350702 224618 350786 224854
rect 351022 224618 368466 224854
rect 368702 224618 368786 224854
rect 369022 224618 386466 224854
rect 386702 224618 386786 224854
rect 387022 224618 404466 224854
rect 404702 224618 404786 224854
rect 405022 224618 422466 224854
rect 422702 224618 422786 224854
rect 423022 224618 440466 224854
rect 440702 224618 440786 224854
rect 441022 224618 458466 224854
rect 458702 224618 458786 224854
rect 459022 224618 476466 224854
rect 476702 224618 476786 224854
rect 477022 224618 494466 224854
rect 494702 224618 494786 224854
rect 495022 224618 512466 224854
rect 512702 224618 512786 224854
rect 513022 224618 530466 224854
rect 530702 224618 530786 224854
rect 531022 224618 545964 224854
rect 546200 224618 546284 224854
rect 546520 224618 548472 224854
rect -4476 224586 548472 224618
rect -4476 221454 548472 221486
rect -4476 221218 -1564 221454
rect -1328 221218 -1244 221454
rect -1008 221218 4746 221454
rect 4982 221218 5066 221454
rect 5302 221218 22746 221454
rect 22982 221218 23066 221454
rect 23302 221218 40746 221454
rect 40982 221218 41066 221454
rect 41302 221218 58746 221454
rect 58982 221218 59066 221454
rect 59302 221218 76746 221454
rect 76982 221218 77066 221454
rect 77302 221218 94746 221454
rect 94982 221218 95066 221454
rect 95302 221218 112746 221454
rect 112982 221218 113066 221454
rect 113302 221218 130746 221454
rect 130982 221218 131066 221454
rect 131302 221218 148746 221454
rect 148982 221218 149066 221454
rect 149302 221218 166746 221454
rect 166982 221218 167066 221454
rect 167302 221218 184746 221454
rect 184982 221218 185066 221454
rect 185302 221218 202746 221454
rect 202982 221218 203066 221454
rect 203302 221218 220746 221454
rect 220982 221218 221066 221454
rect 221302 221218 238746 221454
rect 238982 221218 239066 221454
rect 239302 221218 256746 221454
rect 256982 221218 257066 221454
rect 257302 221218 274746 221454
rect 274982 221218 275066 221454
rect 275302 221218 292746 221454
rect 292982 221218 293066 221454
rect 293302 221218 310746 221454
rect 310982 221218 311066 221454
rect 311302 221218 328746 221454
rect 328982 221218 329066 221454
rect 329302 221218 346746 221454
rect 346982 221218 347066 221454
rect 347302 221218 364746 221454
rect 364982 221218 365066 221454
rect 365302 221218 382746 221454
rect 382982 221218 383066 221454
rect 383302 221218 400746 221454
rect 400982 221218 401066 221454
rect 401302 221218 418746 221454
rect 418982 221218 419066 221454
rect 419302 221218 436746 221454
rect 436982 221218 437066 221454
rect 437302 221218 454746 221454
rect 454982 221218 455066 221454
rect 455302 221218 472746 221454
rect 472982 221218 473066 221454
rect 473302 221218 490746 221454
rect 490982 221218 491066 221454
rect 491302 221218 508746 221454
rect 508982 221218 509066 221454
rect 509302 221218 526746 221454
rect 526982 221218 527066 221454
rect 527302 221218 545004 221454
rect 545240 221218 545324 221454
rect 545560 221218 548472 221454
rect -4476 221134 548472 221218
rect -4476 220898 -1564 221134
rect -1328 220898 -1244 221134
rect -1008 220898 4746 221134
rect 4982 220898 5066 221134
rect 5302 220898 22746 221134
rect 22982 220898 23066 221134
rect 23302 220898 40746 221134
rect 40982 220898 41066 221134
rect 41302 220898 58746 221134
rect 58982 220898 59066 221134
rect 59302 220898 76746 221134
rect 76982 220898 77066 221134
rect 77302 220898 94746 221134
rect 94982 220898 95066 221134
rect 95302 220898 112746 221134
rect 112982 220898 113066 221134
rect 113302 220898 130746 221134
rect 130982 220898 131066 221134
rect 131302 220898 148746 221134
rect 148982 220898 149066 221134
rect 149302 220898 166746 221134
rect 166982 220898 167066 221134
rect 167302 220898 184746 221134
rect 184982 220898 185066 221134
rect 185302 220898 202746 221134
rect 202982 220898 203066 221134
rect 203302 220898 220746 221134
rect 220982 220898 221066 221134
rect 221302 220898 238746 221134
rect 238982 220898 239066 221134
rect 239302 220898 256746 221134
rect 256982 220898 257066 221134
rect 257302 220898 274746 221134
rect 274982 220898 275066 221134
rect 275302 220898 292746 221134
rect 292982 220898 293066 221134
rect 293302 220898 310746 221134
rect 310982 220898 311066 221134
rect 311302 220898 328746 221134
rect 328982 220898 329066 221134
rect 329302 220898 346746 221134
rect 346982 220898 347066 221134
rect 347302 220898 364746 221134
rect 364982 220898 365066 221134
rect 365302 220898 382746 221134
rect 382982 220898 383066 221134
rect 383302 220898 400746 221134
rect 400982 220898 401066 221134
rect 401302 220898 418746 221134
rect 418982 220898 419066 221134
rect 419302 220898 436746 221134
rect 436982 220898 437066 221134
rect 437302 220898 454746 221134
rect 454982 220898 455066 221134
rect 455302 220898 472746 221134
rect 472982 220898 473066 221134
rect 473302 220898 490746 221134
rect 490982 220898 491066 221134
rect 491302 220898 508746 221134
rect 508982 220898 509066 221134
rect 509302 220898 526746 221134
rect 526982 220898 527066 221134
rect 527302 220898 545004 221134
rect 545240 220898 545324 221134
rect 545560 220898 548472 221134
rect -4476 220866 548472 220898
rect -4476 214614 548472 214646
rect -4476 214378 -4444 214614
rect -4208 214378 -4124 214614
rect -3888 214378 15906 214614
rect 16142 214378 16226 214614
rect 16462 214378 33906 214614
rect 34142 214378 34226 214614
rect 34462 214378 51906 214614
rect 52142 214378 52226 214614
rect 52462 214378 69906 214614
rect 70142 214378 70226 214614
rect 70462 214378 87906 214614
rect 88142 214378 88226 214614
rect 88462 214378 105906 214614
rect 106142 214378 106226 214614
rect 106462 214378 123906 214614
rect 124142 214378 124226 214614
rect 124462 214378 141906 214614
rect 142142 214378 142226 214614
rect 142462 214378 159906 214614
rect 160142 214378 160226 214614
rect 160462 214378 177906 214614
rect 178142 214378 178226 214614
rect 178462 214378 195906 214614
rect 196142 214378 196226 214614
rect 196462 214378 213906 214614
rect 214142 214378 214226 214614
rect 214462 214378 231906 214614
rect 232142 214378 232226 214614
rect 232462 214378 249906 214614
rect 250142 214378 250226 214614
rect 250462 214378 267906 214614
rect 268142 214378 268226 214614
rect 268462 214378 285906 214614
rect 286142 214378 286226 214614
rect 286462 214378 303906 214614
rect 304142 214378 304226 214614
rect 304462 214378 321906 214614
rect 322142 214378 322226 214614
rect 322462 214378 339906 214614
rect 340142 214378 340226 214614
rect 340462 214378 357906 214614
rect 358142 214378 358226 214614
rect 358462 214378 375906 214614
rect 376142 214378 376226 214614
rect 376462 214378 393906 214614
rect 394142 214378 394226 214614
rect 394462 214378 411906 214614
rect 412142 214378 412226 214614
rect 412462 214378 429906 214614
rect 430142 214378 430226 214614
rect 430462 214378 447906 214614
rect 448142 214378 448226 214614
rect 448462 214378 465906 214614
rect 466142 214378 466226 214614
rect 466462 214378 483906 214614
rect 484142 214378 484226 214614
rect 484462 214378 501906 214614
rect 502142 214378 502226 214614
rect 502462 214378 519906 214614
rect 520142 214378 520226 214614
rect 520462 214378 537906 214614
rect 538142 214378 538226 214614
rect 538462 214378 547884 214614
rect 548120 214378 548204 214614
rect 548440 214378 548472 214614
rect -4476 214294 548472 214378
rect -4476 214058 -4444 214294
rect -4208 214058 -4124 214294
rect -3888 214058 15906 214294
rect 16142 214058 16226 214294
rect 16462 214058 33906 214294
rect 34142 214058 34226 214294
rect 34462 214058 51906 214294
rect 52142 214058 52226 214294
rect 52462 214058 69906 214294
rect 70142 214058 70226 214294
rect 70462 214058 87906 214294
rect 88142 214058 88226 214294
rect 88462 214058 105906 214294
rect 106142 214058 106226 214294
rect 106462 214058 123906 214294
rect 124142 214058 124226 214294
rect 124462 214058 141906 214294
rect 142142 214058 142226 214294
rect 142462 214058 159906 214294
rect 160142 214058 160226 214294
rect 160462 214058 177906 214294
rect 178142 214058 178226 214294
rect 178462 214058 195906 214294
rect 196142 214058 196226 214294
rect 196462 214058 213906 214294
rect 214142 214058 214226 214294
rect 214462 214058 231906 214294
rect 232142 214058 232226 214294
rect 232462 214058 249906 214294
rect 250142 214058 250226 214294
rect 250462 214058 267906 214294
rect 268142 214058 268226 214294
rect 268462 214058 285906 214294
rect 286142 214058 286226 214294
rect 286462 214058 303906 214294
rect 304142 214058 304226 214294
rect 304462 214058 321906 214294
rect 322142 214058 322226 214294
rect 322462 214058 339906 214294
rect 340142 214058 340226 214294
rect 340462 214058 357906 214294
rect 358142 214058 358226 214294
rect 358462 214058 375906 214294
rect 376142 214058 376226 214294
rect 376462 214058 393906 214294
rect 394142 214058 394226 214294
rect 394462 214058 411906 214294
rect 412142 214058 412226 214294
rect 412462 214058 429906 214294
rect 430142 214058 430226 214294
rect 430462 214058 447906 214294
rect 448142 214058 448226 214294
rect 448462 214058 465906 214294
rect 466142 214058 466226 214294
rect 466462 214058 483906 214294
rect 484142 214058 484226 214294
rect 484462 214058 501906 214294
rect 502142 214058 502226 214294
rect 502462 214058 519906 214294
rect 520142 214058 520226 214294
rect 520462 214058 537906 214294
rect 538142 214058 538226 214294
rect 538462 214058 547884 214294
rect 548120 214058 548204 214294
rect 548440 214058 548472 214294
rect -4476 214026 548472 214058
rect -4476 210894 548472 210926
rect -4476 210658 -3484 210894
rect -3248 210658 -3164 210894
rect -2928 210658 12186 210894
rect 12422 210658 12506 210894
rect 12742 210658 30186 210894
rect 30422 210658 30506 210894
rect 30742 210658 48186 210894
rect 48422 210658 48506 210894
rect 48742 210658 66186 210894
rect 66422 210658 66506 210894
rect 66742 210658 84186 210894
rect 84422 210658 84506 210894
rect 84742 210658 102186 210894
rect 102422 210658 102506 210894
rect 102742 210658 120186 210894
rect 120422 210658 120506 210894
rect 120742 210658 138186 210894
rect 138422 210658 138506 210894
rect 138742 210658 156186 210894
rect 156422 210658 156506 210894
rect 156742 210658 174186 210894
rect 174422 210658 174506 210894
rect 174742 210658 192186 210894
rect 192422 210658 192506 210894
rect 192742 210658 210186 210894
rect 210422 210658 210506 210894
rect 210742 210658 228186 210894
rect 228422 210658 228506 210894
rect 228742 210658 246186 210894
rect 246422 210658 246506 210894
rect 246742 210658 264186 210894
rect 264422 210658 264506 210894
rect 264742 210658 282186 210894
rect 282422 210658 282506 210894
rect 282742 210658 300186 210894
rect 300422 210658 300506 210894
rect 300742 210658 318186 210894
rect 318422 210658 318506 210894
rect 318742 210658 336186 210894
rect 336422 210658 336506 210894
rect 336742 210658 354186 210894
rect 354422 210658 354506 210894
rect 354742 210658 372186 210894
rect 372422 210658 372506 210894
rect 372742 210658 390186 210894
rect 390422 210658 390506 210894
rect 390742 210658 408186 210894
rect 408422 210658 408506 210894
rect 408742 210658 426186 210894
rect 426422 210658 426506 210894
rect 426742 210658 444186 210894
rect 444422 210658 444506 210894
rect 444742 210658 462186 210894
rect 462422 210658 462506 210894
rect 462742 210658 480186 210894
rect 480422 210658 480506 210894
rect 480742 210658 498186 210894
rect 498422 210658 498506 210894
rect 498742 210658 516186 210894
rect 516422 210658 516506 210894
rect 516742 210658 534186 210894
rect 534422 210658 534506 210894
rect 534742 210658 546924 210894
rect 547160 210658 547244 210894
rect 547480 210658 548472 210894
rect -4476 210574 548472 210658
rect -4476 210338 -3484 210574
rect -3248 210338 -3164 210574
rect -2928 210338 12186 210574
rect 12422 210338 12506 210574
rect 12742 210338 30186 210574
rect 30422 210338 30506 210574
rect 30742 210338 48186 210574
rect 48422 210338 48506 210574
rect 48742 210338 66186 210574
rect 66422 210338 66506 210574
rect 66742 210338 84186 210574
rect 84422 210338 84506 210574
rect 84742 210338 102186 210574
rect 102422 210338 102506 210574
rect 102742 210338 120186 210574
rect 120422 210338 120506 210574
rect 120742 210338 138186 210574
rect 138422 210338 138506 210574
rect 138742 210338 156186 210574
rect 156422 210338 156506 210574
rect 156742 210338 174186 210574
rect 174422 210338 174506 210574
rect 174742 210338 192186 210574
rect 192422 210338 192506 210574
rect 192742 210338 210186 210574
rect 210422 210338 210506 210574
rect 210742 210338 228186 210574
rect 228422 210338 228506 210574
rect 228742 210338 246186 210574
rect 246422 210338 246506 210574
rect 246742 210338 264186 210574
rect 264422 210338 264506 210574
rect 264742 210338 282186 210574
rect 282422 210338 282506 210574
rect 282742 210338 300186 210574
rect 300422 210338 300506 210574
rect 300742 210338 318186 210574
rect 318422 210338 318506 210574
rect 318742 210338 336186 210574
rect 336422 210338 336506 210574
rect 336742 210338 354186 210574
rect 354422 210338 354506 210574
rect 354742 210338 372186 210574
rect 372422 210338 372506 210574
rect 372742 210338 390186 210574
rect 390422 210338 390506 210574
rect 390742 210338 408186 210574
rect 408422 210338 408506 210574
rect 408742 210338 426186 210574
rect 426422 210338 426506 210574
rect 426742 210338 444186 210574
rect 444422 210338 444506 210574
rect 444742 210338 462186 210574
rect 462422 210338 462506 210574
rect 462742 210338 480186 210574
rect 480422 210338 480506 210574
rect 480742 210338 498186 210574
rect 498422 210338 498506 210574
rect 498742 210338 516186 210574
rect 516422 210338 516506 210574
rect 516742 210338 534186 210574
rect 534422 210338 534506 210574
rect 534742 210338 546924 210574
rect 547160 210338 547244 210574
rect 547480 210338 548472 210574
rect -4476 210306 548472 210338
rect -4476 207174 548472 207206
rect -4476 206938 -2524 207174
rect -2288 206938 -2204 207174
rect -1968 206938 8466 207174
rect 8702 206938 8786 207174
rect 9022 206938 26466 207174
rect 26702 206938 26786 207174
rect 27022 206938 44466 207174
rect 44702 206938 44786 207174
rect 45022 206938 62466 207174
rect 62702 206938 62786 207174
rect 63022 206938 80466 207174
rect 80702 206938 80786 207174
rect 81022 206938 98466 207174
rect 98702 206938 98786 207174
rect 99022 206938 116466 207174
rect 116702 206938 116786 207174
rect 117022 206938 134466 207174
rect 134702 206938 134786 207174
rect 135022 206938 152466 207174
rect 152702 206938 152786 207174
rect 153022 206938 170466 207174
rect 170702 206938 170786 207174
rect 171022 206938 188466 207174
rect 188702 206938 188786 207174
rect 189022 206938 206466 207174
rect 206702 206938 206786 207174
rect 207022 206938 224466 207174
rect 224702 206938 224786 207174
rect 225022 206938 242466 207174
rect 242702 206938 242786 207174
rect 243022 206938 260466 207174
rect 260702 206938 260786 207174
rect 261022 206938 278466 207174
rect 278702 206938 278786 207174
rect 279022 206938 296466 207174
rect 296702 206938 296786 207174
rect 297022 206938 314466 207174
rect 314702 206938 314786 207174
rect 315022 206938 332466 207174
rect 332702 206938 332786 207174
rect 333022 206938 350466 207174
rect 350702 206938 350786 207174
rect 351022 206938 368466 207174
rect 368702 206938 368786 207174
rect 369022 206938 386466 207174
rect 386702 206938 386786 207174
rect 387022 206938 404466 207174
rect 404702 206938 404786 207174
rect 405022 206938 422466 207174
rect 422702 206938 422786 207174
rect 423022 206938 440466 207174
rect 440702 206938 440786 207174
rect 441022 206938 458466 207174
rect 458702 206938 458786 207174
rect 459022 206938 476466 207174
rect 476702 206938 476786 207174
rect 477022 206938 494466 207174
rect 494702 206938 494786 207174
rect 495022 206938 512466 207174
rect 512702 206938 512786 207174
rect 513022 206938 530466 207174
rect 530702 206938 530786 207174
rect 531022 206938 545964 207174
rect 546200 206938 546284 207174
rect 546520 206938 548472 207174
rect -4476 206854 548472 206938
rect -4476 206618 -2524 206854
rect -2288 206618 -2204 206854
rect -1968 206618 8466 206854
rect 8702 206618 8786 206854
rect 9022 206618 26466 206854
rect 26702 206618 26786 206854
rect 27022 206618 44466 206854
rect 44702 206618 44786 206854
rect 45022 206618 62466 206854
rect 62702 206618 62786 206854
rect 63022 206618 80466 206854
rect 80702 206618 80786 206854
rect 81022 206618 98466 206854
rect 98702 206618 98786 206854
rect 99022 206618 116466 206854
rect 116702 206618 116786 206854
rect 117022 206618 134466 206854
rect 134702 206618 134786 206854
rect 135022 206618 152466 206854
rect 152702 206618 152786 206854
rect 153022 206618 170466 206854
rect 170702 206618 170786 206854
rect 171022 206618 188466 206854
rect 188702 206618 188786 206854
rect 189022 206618 206466 206854
rect 206702 206618 206786 206854
rect 207022 206618 224466 206854
rect 224702 206618 224786 206854
rect 225022 206618 242466 206854
rect 242702 206618 242786 206854
rect 243022 206618 260466 206854
rect 260702 206618 260786 206854
rect 261022 206618 278466 206854
rect 278702 206618 278786 206854
rect 279022 206618 296466 206854
rect 296702 206618 296786 206854
rect 297022 206618 314466 206854
rect 314702 206618 314786 206854
rect 315022 206618 332466 206854
rect 332702 206618 332786 206854
rect 333022 206618 350466 206854
rect 350702 206618 350786 206854
rect 351022 206618 368466 206854
rect 368702 206618 368786 206854
rect 369022 206618 386466 206854
rect 386702 206618 386786 206854
rect 387022 206618 404466 206854
rect 404702 206618 404786 206854
rect 405022 206618 422466 206854
rect 422702 206618 422786 206854
rect 423022 206618 440466 206854
rect 440702 206618 440786 206854
rect 441022 206618 458466 206854
rect 458702 206618 458786 206854
rect 459022 206618 476466 206854
rect 476702 206618 476786 206854
rect 477022 206618 494466 206854
rect 494702 206618 494786 206854
rect 495022 206618 512466 206854
rect 512702 206618 512786 206854
rect 513022 206618 530466 206854
rect 530702 206618 530786 206854
rect 531022 206618 545964 206854
rect 546200 206618 546284 206854
rect 546520 206618 548472 206854
rect -4476 206586 548472 206618
rect -4476 203454 548472 203486
rect -4476 203218 -1564 203454
rect -1328 203218 -1244 203454
rect -1008 203218 4746 203454
rect 4982 203218 5066 203454
rect 5302 203218 22746 203454
rect 22982 203218 23066 203454
rect 23302 203218 40746 203454
rect 40982 203218 41066 203454
rect 41302 203218 58746 203454
rect 58982 203218 59066 203454
rect 59302 203218 76746 203454
rect 76982 203218 77066 203454
rect 77302 203218 94746 203454
rect 94982 203218 95066 203454
rect 95302 203218 112746 203454
rect 112982 203218 113066 203454
rect 113302 203218 130746 203454
rect 130982 203218 131066 203454
rect 131302 203218 148746 203454
rect 148982 203218 149066 203454
rect 149302 203218 166746 203454
rect 166982 203218 167066 203454
rect 167302 203218 184746 203454
rect 184982 203218 185066 203454
rect 185302 203218 202746 203454
rect 202982 203218 203066 203454
rect 203302 203218 220746 203454
rect 220982 203218 221066 203454
rect 221302 203218 238746 203454
rect 238982 203218 239066 203454
rect 239302 203218 256746 203454
rect 256982 203218 257066 203454
rect 257302 203218 274746 203454
rect 274982 203218 275066 203454
rect 275302 203218 292746 203454
rect 292982 203218 293066 203454
rect 293302 203218 310746 203454
rect 310982 203218 311066 203454
rect 311302 203218 328746 203454
rect 328982 203218 329066 203454
rect 329302 203218 346746 203454
rect 346982 203218 347066 203454
rect 347302 203218 364746 203454
rect 364982 203218 365066 203454
rect 365302 203218 382746 203454
rect 382982 203218 383066 203454
rect 383302 203218 400746 203454
rect 400982 203218 401066 203454
rect 401302 203218 418746 203454
rect 418982 203218 419066 203454
rect 419302 203218 436746 203454
rect 436982 203218 437066 203454
rect 437302 203218 454746 203454
rect 454982 203218 455066 203454
rect 455302 203218 472746 203454
rect 472982 203218 473066 203454
rect 473302 203218 490746 203454
rect 490982 203218 491066 203454
rect 491302 203218 508746 203454
rect 508982 203218 509066 203454
rect 509302 203218 526746 203454
rect 526982 203218 527066 203454
rect 527302 203218 545004 203454
rect 545240 203218 545324 203454
rect 545560 203218 548472 203454
rect -4476 203134 548472 203218
rect -4476 202898 -1564 203134
rect -1328 202898 -1244 203134
rect -1008 202898 4746 203134
rect 4982 202898 5066 203134
rect 5302 202898 22746 203134
rect 22982 202898 23066 203134
rect 23302 202898 40746 203134
rect 40982 202898 41066 203134
rect 41302 202898 58746 203134
rect 58982 202898 59066 203134
rect 59302 202898 76746 203134
rect 76982 202898 77066 203134
rect 77302 202898 94746 203134
rect 94982 202898 95066 203134
rect 95302 202898 112746 203134
rect 112982 202898 113066 203134
rect 113302 202898 130746 203134
rect 130982 202898 131066 203134
rect 131302 202898 148746 203134
rect 148982 202898 149066 203134
rect 149302 202898 166746 203134
rect 166982 202898 167066 203134
rect 167302 202898 184746 203134
rect 184982 202898 185066 203134
rect 185302 202898 202746 203134
rect 202982 202898 203066 203134
rect 203302 202898 220746 203134
rect 220982 202898 221066 203134
rect 221302 202898 238746 203134
rect 238982 202898 239066 203134
rect 239302 202898 256746 203134
rect 256982 202898 257066 203134
rect 257302 202898 274746 203134
rect 274982 202898 275066 203134
rect 275302 202898 292746 203134
rect 292982 202898 293066 203134
rect 293302 202898 310746 203134
rect 310982 202898 311066 203134
rect 311302 202898 328746 203134
rect 328982 202898 329066 203134
rect 329302 202898 346746 203134
rect 346982 202898 347066 203134
rect 347302 202898 364746 203134
rect 364982 202898 365066 203134
rect 365302 202898 382746 203134
rect 382982 202898 383066 203134
rect 383302 202898 400746 203134
rect 400982 202898 401066 203134
rect 401302 202898 418746 203134
rect 418982 202898 419066 203134
rect 419302 202898 436746 203134
rect 436982 202898 437066 203134
rect 437302 202898 454746 203134
rect 454982 202898 455066 203134
rect 455302 202898 472746 203134
rect 472982 202898 473066 203134
rect 473302 202898 490746 203134
rect 490982 202898 491066 203134
rect 491302 202898 508746 203134
rect 508982 202898 509066 203134
rect 509302 202898 526746 203134
rect 526982 202898 527066 203134
rect 527302 202898 545004 203134
rect 545240 202898 545324 203134
rect 545560 202898 548472 203134
rect -4476 202866 548472 202898
rect -4476 196614 548472 196646
rect -4476 196378 -4444 196614
rect -4208 196378 -4124 196614
rect -3888 196378 15906 196614
rect 16142 196378 16226 196614
rect 16462 196378 33906 196614
rect 34142 196378 34226 196614
rect 34462 196378 51906 196614
rect 52142 196378 52226 196614
rect 52462 196378 69906 196614
rect 70142 196378 70226 196614
rect 70462 196378 87906 196614
rect 88142 196378 88226 196614
rect 88462 196378 105906 196614
rect 106142 196378 106226 196614
rect 106462 196378 123906 196614
rect 124142 196378 124226 196614
rect 124462 196378 141906 196614
rect 142142 196378 142226 196614
rect 142462 196378 159906 196614
rect 160142 196378 160226 196614
rect 160462 196378 177906 196614
rect 178142 196378 178226 196614
rect 178462 196378 195906 196614
rect 196142 196378 196226 196614
rect 196462 196378 213906 196614
rect 214142 196378 214226 196614
rect 214462 196378 231906 196614
rect 232142 196378 232226 196614
rect 232462 196378 249906 196614
rect 250142 196378 250226 196614
rect 250462 196378 267906 196614
rect 268142 196378 268226 196614
rect 268462 196378 285906 196614
rect 286142 196378 286226 196614
rect 286462 196378 303906 196614
rect 304142 196378 304226 196614
rect 304462 196378 321906 196614
rect 322142 196378 322226 196614
rect 322462 196378 339906 196614
rect 340142 196378 340226 196614
rect 340462 196378 357906 196614
rect 358142 196378 358226 196614
rect 358462 196378 375906 196614
rect 376142 196378 376226 196614
rect 376462 196378 393906 196614
rect 394142 196378 394226 196614
rect 394462 196378 411906 196614
rect 412142 196378 412226 196614
rect 412462 196378 429906 196614
rect 430142 196378 430226 196614
rect 430462 196378 447906 196614
rect 448142 196378 448226 196614
rect 448462 196378 465906 196614
rect 466142 196378 466226 196614
rect 466462 196378 483906 196614
rect 484142 196378 484226 196614
rect 484462 196378 501906 196614
rect 502142 196378 502226 196614
rect 502462 196378 519906 196614
rect 520142 196378 520226 196614
rect 520462 196378 537906 196614
rect 538142 196378 538226 196614
rect 538462 196378 547884 196614
rect 548120 196378 548204 196614
rect 548440 196378 548472 196614
rect -4476 196294 548472 196378
rect -4476 196058 -4444 196294
rect -4208 196058 -4124 196294
rect -3888 196058 15906 196294
rect 16142 196058 16226 196294
rect 16462 196058 33906 196294
rect 34142 196058 34226 196294
rect 34462 196058 51906 196294
rect 52142 196058 52226 196294
rect 52462 196058 69906 196294
rect 70142 196058 70226 196294
rect 70462 196058 87906 196294
rect 88142 196058 88226 196294
rect 88462 196058 105906 196294
rect 106142 196058 106226 196294
rect 106462 196058 123906 196294
rect 124142 196058 124226 196294
rect 124462 196058 141906 196294
rect 142142 196058 142226 196294
rect 142462 196058 159906 196294
rect 160142 196058 160226 196294
rect 160462 196058 177906 196294
rect 178142 196058 178226 196294
rect 178462 196058 195906 196294
rect 196142 196058 196226 196294
rect 196462 196058 213906 196294
rect 214142 196058 214226 196294
rect 214462 196058 231906 196294
rect 232142 196058 232226 196294
rect 232462 196058 249906 196294
rect 250142 196058 250226 196294
rect 250462 196058 267906 196294
rect 268142 196058 268226 196294
rect 268462 196058 285906 196294
rect 286142 196058 286226 196294
rect 286462 196058 303906 196294
rect 304142 196058 304226 196294
rect 304462 196058 321906 196294
rect 322142 196058 322226 196294
rect 322462 196058 339906 196294
rect 340142 196058 340226 196294
rect 340462 196058 357906 196294
rect 358142 196058 358226 196294
rect 358462 196058 375906 196294
rect 376142 196058 376226 196294
rect 376462 196058 393906 196294
rect 394142 196058 394226 196294
rect 394462 196058 411906 196294
rect 412142 196058 412226 196294
rect 412462 196058 429906 196294
rect 430142 196058 430226 196294
rect 430462 196058 447906 196294
rect 448142 196058 448226 196294
rect 448462 196058 465906 196294
rect 466142 196058 466226 196294
rect 466462 196058 483906 196294
rect 484142 196058 484226 196294
rect 484462 196058 501906 196294
rect 502142 196058 502226 196294
rect 502462 196058 519906 196294
rect 520142 196058 520226 196294
rect 520462 196058 537906 196294
rect 538142 196058 538226 196294
rect 538462 196058 547884 196294
rect 548120 196058 548204 196294
rect 548440 196058 548472 196294
rect -4476 196026 548472 196058
rect -4476 192894 548472 192926
rect -4476 192658 -3484 192894
rect -3248 192658 -3164 192894
rect -2928 192658 12186 192894
rect 12422 192658 12506 192894
rect 12742 192658 30186 192894
rect 30422 192658 30506 192894
rect 30742 192658 48186 192894
rect 48422 192658 48506 192894
rect 48742 192658 66186 192894
rect 66422 192658 66506 192894
rect 66742 192658 84186 192894
rect 84422 192658 84506 192894
rect 84742 192658 102186 192894
rect 102422 192658 102506 192894
rect 102742 192658 120186 192894
rect 120422 192658 120506 192894
rect 120742 192658 138186 192894
rect 138422 192658 138506 192894
rect 138742 192658 156186 192894
rect 156422 192658 156506 192894
rect 156742 192658 174186 192894
rect 174422 192658 174506 192894
rect 174742 192658 192186 192894
rect 192422 192658 192506 192894
rect 192742 192658 210186 192894
rect 210422 192658 210506 192894
rect 210742 192658 228186 192894
rect 228422 192658 228506 192894
rect 228742 192658 246186 192894
rect 246422 192658 246506 192894
rect 246742 192658 264186 192894
rect 264422 192658 264506 192894
rect 264742 192658 282186 192894
rect 282422 192658 282506 192894
rect 282742 192658 300186 192894
rect 300422 192658 300506 192894
rect 300742 192658 318186 192894
rect 318422 192658 318506 192894
rect 318742 192658 336186 192894
rect 336422 192658 336506 192894
rect 336742 192658 354186 192894
rect 354422 192658 354506 192894
rect 354742 192658 372186 192894
rect 372422 192658 372506 192894
rect 372742 192658 390186 192894
rect 390422 192658 390506 192894
rect 390742 192658 408186 192894
rect 408422 192658 408506 192894
rect 408742 192658 426186 192894
rect 426422 192658 426506 192894
rect 426742 192658 444186 192894
rect 444422 192658 444506 192894
rect 444742 192658 462186 192894
rect 462422 192658 462506 192894
rect 462742 192658 480186 192894
rect 480422 192658 480506 192894
rect 480742 192658 498186 192894
rect 498422 192658 498506 192894
rect 498742 192658 516186 192894
rect 516422 192658 516506 192894
rect 516742 192658 534186 192894
rect 534422 192658 534506 192894
rect 534742 192658 546924 192894
rect 547160 192658 547244 192894
rect 547480 192658 548472 192894
rect -4476 192574 548472 192658
rect -4476 192338 -3484 192574
rect -3248 192338 -3164 192574
rect -2928 192338 12186 192574
rect 12422 192338 12506 192574
rect 12742 192338 30186 192574
rect 30422 192338 30506 192574
rect 30742 192338 48186 192574
rect 48422 192338 48506 192574
rect 48742 192338 66186 192574
rect 66422 192338 66506 192574
rect 66742 192338 84186 192574
rect 84422 192338 84506 192574
rect 84742 192338 102186 192574
rect 102422 192338 102506 192574
rect 102742 192338 120186 192574
rect 120422 192338 120506 192574
rect 120742 192338 138186 192574
rect 138422 192338 138506 192574
rect 138742 192338 156186 192574
rect 156422 192338 156506 192574
rect 156742 192338 174186 192574
rect 174422 192338 174506 192574
rect 174742 192338 192186 192574
rect 192422 192338 192506 192574
rect 192742 192338 210186 192574
rect 210422 192338 210506 192574
rect 210742 192338 228186 192574
rect 228422 192338 228506 192574
rect 228742 192338 246186 192574
rect 246422 192338 246506 192574
rect 246742 192338 264186 192574
rect 264422 192338 264506 192574
rect 264742 192338 282186 192574
rect 282422 192338 282506 192574
rect 282742 192338 300186 192574
rect 300422 192338 300506 192574
rect 300742 192338 318186 192574
rect 318422 192338 318506 192574
rect 318742 192338 336186 192574
rect 336422 192338 336506 192574
rect 336742 192338 354186 192574
rect 354422 192338 354506 192574
rect 354742 192338 372186 192574
rect 372422 192338 372506 192574
rect 372742 192338 390186 192574
rect 390422 192338 390506 192574
rect 390742 192338 408186 192574
rect 408422 192338 408506 192574
rect 408742 192338 426186 192574
rect 426422 192338 426506 192574
rect 426742 192338 444186 192574
rect 444422 192338 444506 192574
rect 444742 192338 462186 192574
rect 462422 192338 462506 192574
rect 462742 192338 480186 192574
rect 480422 192338 480506 192574
rect 480742 192338 498186 192574
rect 498422 192338 498506 192574
rect 498742 192338 516186 192574
rect 516422 192338 516506 192574
rect 516742 192338 534186 192574
rect 534422 192338 534506 192574
rect 534742 192338 546924 192574
rect 547160 192338 547244 192574
rect 547480 192338 548472 192574
rect -4476 192306 548472 192338
rect -4476 189174 548472 189206
rect -4476 188938 -2524 189174
rect -2288 188938 -2204 189174
rect -1968 188938 8466 189174
rect 8702 188938 8786 189174
rect 9022 188938 26466 189174
rect 26702 188938 26786 189174
rect 27022 188938 44466 189174
rect 44702 188938 44786 189174
rect 45022 188938 62466 189174
rect 62702 188938 62786 189174
rect 63022 188938 80466 189174
rect 80702 188938 80786 189174
rect 81022 188938 98466 189174
rect 98702 188938 98786 189174
rect 99022 188938 116466 189174
rect 116702 188938 116786 189174
rect 117022 188938 134466 189174
rect 134702 188938 134786 189174
rect 135022 188938 152466 189174
rect 152702 188938 152786 189174
rect 153022 188938 170466 189174
rect 170702 188938 170786 189174
rect 171022 188938 188466 189174
rect 188702 188938 188786 189174
rect 189022 188938 206466 189174
rect 206702 188938 206786 189174
rect 207022 188938 224466 189174
rect 224702 188938 224786 189174
rect 225022 188938 242466 189174
rect 242702 188938 242786 189174
rect 243022 188938 260466 189174
rect 260702 188938 260786 189174
rect 261022 188938 278466 189174
rect 278702 188938 278786 189174
rect 279022 188938 296466 189174
rect 296702 188938 296786 189174
rect 297022 188938 314466 189174
rect 314702 188938 314786 189174
rect 315022 188938 332466 189174
rect 332702 188938 332786 189174
rect 333022 188938 350466 189174
rect 350702 188938 350786 189174
rect 351022 188938 368466 189174
rect 368702 188938 368786 189174
rect 369022 188938 386466 189174
rect 386702 188938 386786 189174
rect 387022 188938 404466 189174
rect 404702 188938 404786 189174
rect 405022 188938 422466 189174
rect 422702 188938 422786 189174
rect 423022 188938 440466 189174
rect 440702 188938 440786 189174
rect 441022 188938 458466 189174
rect 458702 188938 458786 189174
rect 459022 188938 476466 189174
rect 476702 188938 476786 189174
rect 477022 188938 494466 189174
rect 494702 188938 494786 189174
rect 495022 188938 512466 189174
rect 512702 188938 512786 189174
rect 513022 188938 530466 189174
rect 530702 188938 530786 189174
rect 531022 188938 545964 189174
rect 546200 188938 546284 189174
rect 546520 188938 548472 189174
rect -4476 188854 548472 188938
rect -4476 188618 -2524 188854
rect -2288 188618 -2204 188854
rect -1968 188618 8466 188854
rect 8702 188618 8786 188854
rect 9022 188618 26466 188854
rect 26702 188618 26786 188854
rect 27022 188618 44466 188854
rect 44702 188618 44786 188854
rect 45022 188618 62466 188854
rect 62702 188618 62786 188854
rect 63022 188618 80466 188854
rect 80702 188618 80786 188854
rect 81022 188618 98466 188854
rect 98702 188618 98786 188854
rect 99022 188618 116466 188854
rect 116702 188618 116786 188854
rect 117022 188618 134466 188854
rect 134702 188618 134786 188854
rect 135022 188618 152466 188854
rect 152702 188618 152786 188854
rect 153022 188618 170466 188854
rect 170702 188618 170786 188854
rect 171022 188618 188466 188854
rect 188702 188618 188786 188854
rect 189022 188618 206466 188854
rect 206702 188618 206786 188854
rect 207022 188618 224466 188854
rect 224702 188618 224786 188854
rect 225022 188618 242466 188854
rect 242702 188618 242786 188854
rect 243022 188618 260466 188854
rect 260702 188618 260786 188854
rect 261022 188618 278466 188854
rect 278702 188618 278786 188854
rect 279022 188618 296466 188854
rect 296702 188618 296786 188854
rect 297022 188618 314466 188854
rect 314702 188618 314786 188854
rect 315022 188618 332466 188854
rect 332702 188618 332786 188854
rect 333022 188618 350466 188854
rect 350702 188618 350786 188854
rect 351022 188618 368466 188854
rect 368702 188618 368786 188854
rect 369022 188618 386466 188854
rect 386702 188618 386786 188854
rect 387022 188618 404466 188854
rect 404702 188618 404786 188854
rect 405022 188618 422466 188854
rect 422702 188618 422786 188854
rect 423022 188618 440466 188854
rect 440702 188618 440786 188854
rect 441022 188618 458466 188854
rect 458702 188618 458786 188854
rect 459022 188618 476466 188854
rect 476702 188618 476786 188854
rect 477022 188618 494466 188854
rect 494702 188618 494786 188854
rect 495022 188618 512466 188854
rect 512702 188618 512786 188854
rect 513022 188618 530466 188854
rect 530702 188618 530786 188854
rect 531022 188618 545964 188854
rect 546200 188618 546284 188854
rect 546520 188618 548472 188854
rect -4476 188586 548472 188618
rect -4476 185454 548472 185486
rect -4476 185218 -1564 185454
rect -1328 185218 -1244 185454
rect -1008 185218 4746 185454
rect 4982 185218 5066 185454
rect 5302 185218 22746 185454
rect 22982 185218 23066 185454
rect 23302 185218 40746 185454
rect 40982 185218 41066 185454
rect 41302 185218 58746 185454
rect 58982 185218 59066 185454
rect 59302 185218 76746 185454
rect 76982 185218 77066 185454
rect 77302 185218 94746 185454
rect 94982 185218 95066 185454
rect 95302 185218 112746 185454
rect 112982 185218 113066 185454
rect 113302 185218 130746 185454
rect 130982 185218 131066 185454
rect 131302 185218 148746 185454
rect 148982 185218 149066 185454
rect 149302 185218 166746 185454
rect 166982 185218 167066 185454
rect 167302 185218 184746 185454
rect 184982 185218 185066 185454
rect 185302 185218 202746 185454
rect 202982 185218 203066 185454
rect 203302 185218 220746 185454
rect 220982 185218 221066 185454
rect 221302 185218 238746 185454
rect 238982 185218 239066 185454
rect 239302 185218 256746 185454
rect 256982 185218 257066 185454
rect 257302 185218 274746 185454
rect 274982 185218 275066 185454
rect 275302 185218 292746 185454
rect 292982 185218 293066 185454
rect 293302 185218 310746 185454
rect 310982 185218 311066 185454
rect 311302 185218 328746 185454
rect 328982 185218 329066 185454
rect 329302 185218 346746 185454
rect 346982 185218 347066 185454
rect 347302 185218 364746 185454
rect 364982 185218 365066 185454
rect 365302 185218 382746 185454
rect 382982 185218 383066 185454
rect 383302 185218 400746 185454
rect 400982 185218 401066 185454
rect 401302 185218 418746 185454
rect 418982 185218 419066 185454
rect 419302 185218 436746 185454
rect 436982 185218 437066 185454
rect 437302 185218 454746 185454
rect 454982 185218 455066 185454
rect 455302 185218 472746 185454
rect 472982 185218 473066 185454
rect 473302 185218 490746 185454
rect 490982 185218 491066 185454
rect 491302 185218 508746 185454
rect 508982 185218 509066 185454
rect 509302 185218 526746 185454
rect 526982 185218 527066 185454
rect 527302 185218 545004 185454
rect 545240 185218 545324 185454
rect 545560 185218 548472 185454
rect -4476 185134 548472 185218
rect -4476 184898 -1564 185134
rect -1328 184898 -1244 185134
rect -1008 184898 4746 185134
rect 4982 184898 5066 185134
rect 5302 184898 22746 185134
rect 22982 184898 23066 185134
rect 23302 184898 40746 185134
rect 40982 184898 41066 185134
rect 41302 184898 58746 185134
rect 58982 184898 59066 185134
rect 59302 184898 76746 185134
rect 76982 184898 77066 185134
rect 77302 184898 94746 185134
rect 94982 184898 95066 185134
rect 95302 184898 112746 185134
rect 112982 184898 113066 185134
rect 113302 184898 130746 185134
rect 130982 184898 131066 185134
rect 131302 184898 148746 185134
rect 148982 184898 149066 185134
rect 149302 184898 166746 185134
rect 166982 184898 167066 185134
rect 167302 184898 184746 185134
rect 184982 184898 185066 185134
rect 185302 184898 202746 185134
rect 202982 184898 203066 185134
rect 203302 184898 220746 185134
rect 220982 184898 221066 185134
rect 221302 184898 238746 185134
rect 238982 184898 239066 185134
rect 239302 184898 256746 185134
rect 256982 184898 257066 185134
rect 257302 184898 274746 185134
rect 274982 184898 275066 185134
rect 275302 184898 292746 185134
rect 292982 184898 293066 185134
rect 293302 184898 310746 185134
rect 310982 184898 311066 185134
rect 311302 184898 328746 185134
rect 328982 184898 329066 185134
rect 329302 184898 346746 185134
rect 346982 184898 347066 185134
rect 347302 184898 364746 185134
rect 364982 184898 365066 185134
rect 365302 184898 382746 185134
rect 382982 184898 383066 185134
rect 383302 184898 400746 185134
rect 400982 184898 401066 185134
rect 401302 184898 418746 185134
rect 418982 184898 419066 185134
rect 419302 184898 436746 185134
rect 436982 184898 437066 185134
rect 437302 184898 454746 185134
rect 454982 184898 455066 185134
rect 455302 184898 472746 185134
rect 472982 184898 473066 185134
rect 473302 184898 490746 185134
rect 490982 184898 491066 185134
rect 491302 184898 508746 185134
rect 508982 184898 509066 185134
rect 509302 184898 526746 185134
rect 526982 184898 527066 185134
rect 527302 184898 545004 185134
rect 545240 184898 545324 185134
rect 545560 184898 548472 185134
rect -4476 184866 548472 184898
rect -4476 178614 548472 178646
rect -4476 178378 -4444 178614
rect -4208 178378 -4124 178614
rect -3888 178378 15906 178614
rect 16142 178378 16226 178614
rect 16462 178378 33906 178614
rect 34142 178378 34226 178614
rect 34462 178378 51906 178614
rect 52142 178378 52226 178614
rect 52462 178378 69906 178614
rect 70142 178378 70226 178614
rect 70462 178378 87906 178614
rect 88142 178378 88226 178614
rect 88462 178378 105906 178614
rect 106142 178378 106226 178614
rect 106462 178378 123906 178614
rect 124142 178378 124226 178614
rect 124462 178378 141906 178614
rect 142142 178378 142226 178614
rect 142462 178378 159906 178614
rect 160142 178378 160226 178614
rect 160462 178378 177906 178614
rect 178142 178378 178226 178614
rect 178462 178378 195906 178614
rect 196142 178378 196226 178614
rect 196462 178378 213906 178614
rect 214142 178378 214226 178614
rect 214462 178378 231906 178614
rect 232142 178378 232226 178614
rect 232462 178378 249906 178614
rect 250142 178378 250226 178614
rect 250462 178378 267906 178614
rect 268142 178378 268226 178614
rect 268462 178378 285906 178614
rect 286142 178378 286226 178614
rect 286462 178378 303906 178614
rect 304142 178378 304226 178614
rect 304462 178378 321906 178614
rect 322142 178378 322226 178614
rect 322462 178378 339906 178614
rect 340142 178378 340226 178614
rect 340462 178378 357906 178614
rect 358142 178378 358226 178614
rect 358462 178378 375906 178614
rect 376142 178378 376226 178614
rect 376462 178378 393906 178614
rect 394142 178378 394226 178614
rect 394462 178378 411906 178614
rect 412142 178378 412226 178614
rect 412462 178378 429906 178614
rect 430142 178378 430226 178614
rect 430462 178378 447906 178614
rect 448142 178378 448226 178614
rect 448462 178378 465906 178614
rect 466142 178378 466226 178614
rect 466462 178378 483906 178614
rect 484142 178378 484226 178614
rect 484462 178378 501906 178614
rect 502142 178378 502226 178614
rect 502462 178378 519906 178614
rect 520142 178378 520226 178614
rect 520462 178378 537906 178614
rect 538142 178378 538226 178614
rect 538462 178378 547884 178614
rect 548120 178378 548204 178614
rect 548440 178378 548472 178614
rect -4476 178294 548472 178378
rect -4476 178058 -4444 178294
rect -4208 178058 -4124 178294
rect -3888 178058 15906 178294
rect 16142 178058 16226 178294
rect 16462 178058 33906 178294
rect 34142 178058 34226 178294
rect 34462 178058 51906 178294
rect 52142 178058 52226 178294
rect 52462 178058 69906 178294
rect 70142 178058 70226 178294
rect 70462 178058 87906 178294
rect 88142 178058 88226 178294
rect 88462 178058 105906 178294
rect 106142 178058 106226 178294
rect 106462 178058 123906 178294
rect 124142 178058 124226 178294
rect 124462 178058 141906 178294
rect 142142 178058 142226 178294
rect 142462 178058 159906 178294
rect 160142 178058 160226 178294
rect 160462 178058 177906 178294
rect 178142 178058 178226 178294
rect 178462 178058 195906 178294
rect 196142 178058 196226 178294
rect 196462 178058 213906 178294
rect 214142 178058 214226 178294
rect 214462 178058 231906 178294
rect 232142 178058 232226 178294
rect 232462 178058 249906 178294
rect 250142 178058 250226 178294
rect 250462 178058 267906 178294
rect 268142 178058 268226 178294
rect 268462 178058 285906 178294
rect 286142 178058 286226 178294
rect 286462 178058 303906 178294
rect 304142 178058 304226 178294
rect 304462 178058 321906 178294
rect 322142 178058 322226 178294
rect 322462 178058 339906 178294
rect 340142 178058 340226 178294
rect 340462 178058 357906 178294
rect 358142 178058 358226 178294
rect 358462 178058 375906 178294
rect 376142 178058 376226 178294
rect 376462 178058 393906 178294
rect 394142 178058 394226 178294
rect 394462 178058 411906 178294
rect 412142 178058 412226 178294
rect 412462 178058 429906 178294
rect 430142 178058 430226 178294
rect 430462 178058 447906 178294
rect 448142 178058 448226 178294
rect 448462 178058 465906 178294
rect 466142 178058 466226 178294
rect 466462 178058 483906 178294
rect 484142 178058 484226 178294
rect 484462 178058 501906 178294
rect 502142 178058 502226 178294
rect 502462 178058 519906 178294
rect 520142 178058 520226 178294
rect 520462 178058 537906 178294
rect 538142 178058 538226 178294
rect 538462 178058 547884 178294
rect 548120 178058 548204 178294
rect 548440 178058 548472 178294
rect -4476 178026 548472 178058
rect -4476 174894 548472 174926
rect -4476 174658 -3484 174894
rect -3248 174658 -3164 174894
rect -2928 174658 12186 174894
rect 12422 174658 12506 174894
rect 12742 174658 30186 174894
rect 30422 174658 30506 174894
rect 30742 174658 48186 174894
rect 48422 174658 48506 174894
rect 48742 174658 66186 174894
rect 66422 174658 66506 174894
rect 66742 174658 84186 174894
rect 84422 174658 84506 174894
rect 84742 174658 102186 174894
rect 102422 174658 102506 174894
rect 102742 174658 120186 174894
rect 120422 174658 120506 174894
rect 120742 174658 138186 174894
rect 138422 174658 138506 174894
rect 138742 174658 156186 174894
rect 156422 174658 156506 174894
rect 156742 174658 174186 174894
rect 174422 174658 174506 174894
rect 174742 174658 192186 174894
rect 192422 174658 192506 174894
rect 192742 174658 210186 174894
rect 210422 174658 210506 174894
rect 210742 174658 228186 174894
rect 228422 174658 228506 174894
rect 228742 174658 246186 174894
rect 246422 174658 246506 174894
rect 246742 174658 264186 174894
rect 264422 174658 264506 174894
rect 264742 174658 282186 174894
rect 282422 174658 282506 174894
rect 282742 174658 300186 174894
rect 300422 174658 300506 174894
rect 300742 174658 318186 174894
rect 318422 174658 318506 174894
rect 318742 174658 336186 174894
rect 336422 174658 336506 174894
rect 336742 174658 354186 174894
rect 354422 174658 354506 174894
rect 354742 174658 372186 174894
rect 372422 174658 372506 174894
rect 372742 174658 390186 174894
rect 390422 174658 390506 174894
rect 390742 174658 408186 174894
rect 408422 174658 408506 174894
rect 408742 174658 426186 174894
rect 426422 174658 426506 174894
rect 426742 174658 444186 174894
rect 444422 174658 444506 174894
rect 444742 174658 462186 174894
rect 462422 174658 462506 174894
rect 462742 174658 480186 174894
rect 480422 174658 480506 174894
rect 480742 174658 498186 174894
rect 498422 174658 498506 174894
rect 498742 174658 516186 174894
rect 516422 174658 516506 174894
rect 516742 174658 534186 174894
rect 534422 174658 534506 174894
rect 534742 174658 546924 174894
rect 547160 174658 547244 174894
rect 547480 174658 548472 174894
rect -4476 174574 548472 174658
rect -4476 174338 -3484 174574
rect -3248 174338 -3164 174574
rect -2928 174338 12186 174574
rect 12422 174338 12506 174574
rect 12742 174338 30186 174574
rect 30422 174338 30506 174574
rect 30742 174338 48186 174574
rect 48422 174338 48506 174574
rect 48742 174338 66186 174574
rect 66422 174338 66506 174574
rect 66742 174338 84186 174574
rect 84422 174338 84506 174574
rect 84742 174338 102186 174574
rect 102422 174338 102506 174574
rect 102742 174338 120186 174574
rect 120422 174338 120506 174574
rect 120742 174338 138186 174574
rect 138422 174338 138506 174574
rect 138742 174338 156186 174574
rect 156422 174338 156506 174574
rect 156742 174338 174186 174574
rect 174422 174338 174506 174574
rect 174742 174338 192186 174574
rect 192422 174338 192506 174574
rect 192742 174338 210186 174574
rect 210422 174338 210506 174574
rect 210742 174338 228186 174574
rect 228422 174338 228506 174574
rect 228742 174338 246186 174574
rect 246422 174338 246506 174574
rect 246742 174338 264186 174574
rect 264422 174338 264506 174574
rect 264742 174338 282186 174574
rect 282422 174338 282506 174574
rect 282742 174338 300186 174574
rect 300422 174338 300506 174574
rect 300742 174338 318186 174574
rect 318422 174338 318506 174574
rect 318742 174338 336186 174574
rect 336422 174338 336506 174574
rect 336742 174338 354186 174574
rect 354422 174338 354506 174574
rect 354742 174338 372186 174574
rect 372422 174338 372506 174574
rect 372742 174338 390186 174574
rect 390422 174338 390506 174574
rect 390742 174338 408186 174574
rect 408422 174338 408506 174574
rect 408742 174338 426186 174574
rect 426422 174338 426506 174574
rect 426742 174338 444186 174574
rect 444422 174338 444506 174574
rect 444742 174338 462186 174574
rect 462422 174338 462506 174574
rect 462742 174338 480186 174574
rect 480422 174338 480506 174574
rect 480742 174338 498186 174574
rect 498422 174338 498506 174574
rect 498742 174338 516186 174574
rect 516422 174338 516506 174574
rect 516742 174338 534186 174574
rect 534422 174338 534506 174574
rect 534742 174338 546924 174574
rect 547160 174338 547244 174574
rect 547480 174338 548472 174574
rect -4476 174306 548472 174338
rect -4476 171174 548472 171206
rect -4476 170938 -2524 171174
rect -2288 170938 -2204 171174
rect -1968 170938 8466 171174
rect 8702 170938 8786 171174
rect 9022 170938 26466 171174
rect 26702 170938 26786 171174
rect 27022 170938 44466 171174
rect 44702 170938 44786 171174
rect 45022 170938 62466 171174
rect 62702 170938 62786 171174
rect 63022 170938 80466 171174
rect 80702 170938 80786 171174
rect 81022 170938 98466 171174
rect 98702 170938 98786 171174
rect 99022 170938 116466 171174
rect 116702 170938 116786 171174
rect 117022 170938 134466 171174
rect 134702 170938 134786 171174
rect 135022 170938 152466 171174
rect 152702 170938 152786 171174
rect 153022 170938 170466 171174
rect 170702 170938 170786 171174
rect 171022 170938 188466 171174
rect 188702 170938 188786 171174
rect 189022 170938 206466 171174
rect 206702 170938 206786 171174
rect 207022 170938 224466 171174
rect 224702 170938 224786 171174
rect 225022 170938 242466 171174
rect 242702 170938 242786 171174
rect 243022 170938 260466 171174
rect 260702 170938 260786 171174
rect 261022 170938 278466 171174
rect 278702 170938 278786 171174
rect 279022 170938 296466 171174
rect 296702 170938 296786 171174
rect 297022 170938 314466 171174
rect 314702 170938 314786 171174
rect 315022 170938 332466 171174
rect 332702 170938 332786 171174
rect 333022 170938 350466 171174
rect 350702 170938 350786 171174
rect 351022 170938 368466 171174
rect 368702 170938 368786 171174
rect 369022 170938 386466 171174
rect 386702 170938 386786 171174
rect 387022 170938 404466 171174
rect 404702 170938 404786 171174
rect 405022 170938 422466 171174
rect 422702 170938 422786 171174
rect 423022 170938 440466 171174
rect 440702 170938 440786 171174
rect 441022 170938 458466 171174
rect 458702 170938 458786 171174
rect 459022 170938 476466 171174
rect 476702 170938 476786 171174
rect 477022 170938 494466 171174
rect 494702 170938 494786 171174
rect 495022 170938 512466 171174
rect 512702 170938 512786 171174
rect 513022 170938 530466 171174
rect 530702 170938 530786 171174
rect 531022 170938 545964 171174
rect 546200 170938 546284 171174
rect 546520 170938 548472 171174
rect -4476 170854 548472 170938
rect -4476 170618 -2524 170854
rect -2288 170618 -2204 170854
rect -1968 170618 8466 170854
rect 8702 170618 8786 170854
rect 9022 170618 26466 170854
rect 26702 170618 26786 170854
rect 27022 170618 44466 170854
rect 44702 170618 44786 170854
rect 45022 170618 62466 170854
rect 62702 170618 62786 170854
rect 63022 170618 80466 170854
rect 80702 170618 80786 170854
rect 81022 170618 98466 170854
rect 98702 170618 98786 170854
rect 99022 170618 116466 170854
rect 116702 170618 116786 170854
rect 117022 170618 134466 170854
rect 134702 170618 134786 170854
rect 135022 170618 152466 170854
rect 152702 170618 152786 170854
rect 153022 170618 170466 170854
rect 170702 170618 170786 170854
rect 171022 170618 188466 170854
rect 188702 170618 188786 170854
rect 189022 170618 206466 170854
rect 206702 170618 206786 170854
rect 207022 170618 224466 170854
rect 224702 170618 224786 170854
rect 225022 170618 242466 170854
rect 242702 170618 242786 170854
rect 243022 170618 260466 170854
rect 260702 170618 260786 170854
rect 261022 170618 278466 170854
rect 278702 170618 278786 170854
rect 279022 170618 296466 170854
rect 296702 170618 296786 170854
rect 297022 170618 314466 170854
rect 314702 170618 314786 170854
rect 315022 170618 332466 170854
rect 332702 170618 332786 170854
rect 333022 170618 350466 170854
rect 350702 170618 350786 170854
rect 351022 170618 368466 170854
rect 368702 170618 368786 170854
rect 369022 170618 386466 170854
rect 386702 170618 386786 170854
rect 387022 170618 404466 170854
rect 404702 170618 404786 170854
rect 405022 170618 422466 170854
rect 422702 170618 422786 170854
rect 423022 170618 440466 170854
rect 440702 170618 440786 170854
rect 441022 170618 458466 170854
rect 458702 170618 458786 170854
rect 459022 170618 476466 170854
rect 476702 170618 476786 170854
rect 477022 170618 494466 170854
rect 494702 170618 494786 170854
rect 495022 170618 512466 170854
rect 512702 170618 512786 170854
rect 513022 170618 530466 170854
rect 530702 170618 530786 170854
rect 531022 170618 545964 170854
rect 546200 170618 546284 170854
rect 546520 170618 548472 170854
rect -4476 170586 548472 170618
rect -4476 167454 548472 167486
rect -4476 167218 -1564 167454
rect -1328 167218 -1244 167454
rect -1008 167218 4746 167454
rect 4982 167218 5066 167454
rect 5302 167218 22746 167454
rect 22982 167218 23066 167454
rect 23302 167218 40746 167454
rect 40982 167218 41066 167454
rect 41302 167218 58746 167454
rect 58982 167218 59066 167454
rect 59302 167218 76746 167454
rect 76982 167218 77066 167454
rect 77302 167218 94746 167454
rect 94982 167218 95066 167454
rect 95302 167218 112746 167454
rect 112982 167218 113066 167454
rect 113302 167218 130746 167454
rect 130982 167218 131066 167454
rect 131302 167218 148746 167454
rect 148982 167218 149066 167454
rect 149302 167218 166746 167454
rect 166982 167218 167066 167454
rect 167302 167218 184746 167454
rect 184982 167218 185066 167454
rect 185302 167218 202746 167454
rect 202982 167218 203066 167454
rect 203302 167218 220746 167454
rect 220982 167218 221066 167454
rect 221302 167218 238746 167454
rect 238982 167218 239066 167454
rect 239302 167218 256746 167454
rect 256982 167218 257066 167454
rect 257302 167218 274746 167454
rect 274982 167218 275066 167454
rect 275302 167218 292746 167454
rect 292982 167218 293066 167454
rect 293302 167218 310746 167454
rect 310982 167218 311066 167454
rect 311302 167218 328746 167454
rect 328982 167218 329066 167454
rect 329302 167218 346746 167454
rect 346982 167218 347066 167454
rect 347302 167218 364746 167454
rect 364982 167218 365066 167454
rect 365302 167218 382746 167454
rect 382982 167218 383066 167454
rect 383302 167218 400746 167454
rect 400982 167218 401066 167454
rect 401302 167218 418746 167454
rect 418982 167218 419066 167454
rect 419302 167218 436746 167454
rect 436982 167218 437066 167454
rect 437302 167218 454746 167454
rect 454982 167218 455066 167454
rect 455302 167218 472746 167454
rect 472982 167218 473066 167454
rect 473302 167218 490746 167454
rect 490982 167218 491066 167454
rect 491302 167218 508746 167454
rect 508982 167218 509066 167454
rect 509302 167218 526746 167454
rect 526982 167218 527066 167454
rect 527302 167218 545004 167454
rect 545240 167218 545324 167454
rect 545560 167218 548472 167454
rect -4476 167134 548472 167218
rect -4476 166898 -1564 167134
rect -1328 166898 -1244 167134
rect -1008 166898 4746 167134
rect 4982 166898 5066 167134
rect 5302 166898 22746 167134
rect 22982 166898 23066 167134
rect 23302 166898 40746 167134
rect 40982 166898 41066 167134
rect 41302 166898 58746 167134
rect 58982 166898 59066 167134
rect 59302 166898 76746 167134
rect 76982 166898 77066 167134
rect 77302 166898 94746 167134
rect 94982 166898 95066 167134
rect 95302 166898 112746 167134
rect 112982 166898 113066 167134
rect 113302 166898 130746 167134
rect 130982 166898 131066 167134
rect 131302 166898 148746 167134
rect 148982 166898 149066 167134
rect 149302 166898 166746 167134
rect 166982 166898 167066 167134
rect 167302 166898 184746 167134
rect 184982 166898 185066 167134
rect 185302 166898 202746 167134
rect 202982 166898 203066 167134
rect 203302 166898 220746 167134
rect 220982 166898 221066 167134
rect 221302 166898 238746 167134
rect 238982 166898 239066 167134
rect 239302 166898 256746 167134
rect 256982 166898 257066 167134
rect 257302 166898 274746 167134
rect 274982 166898 275066 167134
rect 275302 166898 292746 167134
rect 292982 166898 293066 167134
rect 293302 166898 310746 167134
rect 310982 166898 311066 167134
rect 311302 166898 328746 167134
rect 328982 166898 329066 167134
rect 329302 166898 346746 167134
rect 346982 166898 347066 167134
rect 347302 166898 364746 167134
rect 364982 166898 365066 167134
rect 365302 166898 382746 167134
rect 382982 166898 383066 167134
rect 383302 166898 400746 167134
rect 400982 166898 401066 167134
rect 401302 166898 418746 167134
rect 418982 166898 419066 167134
rect 419302 166898 436746 167134
rect 436982 166898 437066 167134
rect 437302 166898 454746 167134
rect 454982 166898 455066 167134
rect 455302 166898 472746 167134
rect 472982 166898 473066 167134
rect 473302 166898 490746 167134
rect 490982 166898 491066 167134
rect 491302 166898 508746 167134
rect 508982 166898 509066 167134
rect 509302 166898 526746 167134
rect 526982 166898 527066 167134
rect 527302 166898 545004 167134
rect 545240 166898 545324 167134
rect 545560 166898 548472 167134
rect -4476 166866 548472 166898
rect -4476 160614 548472 160646
rect -4476 160378 -4444 160614
rect -4208 160378 -4124 160614
rect -3888 160378 15906 160614
rect 16142 160378 16226 160614
rect 16462 160378 33906 160614
rect 34142 160378 34226 160614
rect 34462 160378 51906 160614
rect 52142 160378 52226 160614
rect 52462 160378 69906 160614
rect 70142 160378 70226 160614
rect 70462 160378 87906 160614
rect 88142 160378 88226 160614
rect 88462 160378 105906 160614
rect 106142 160378 106226 160614
rect 106462 160378 123906 160614
rect 124142 160378 124226 160614
rect 124462 160378 141906 160614
rect 142142 160378 142226 160614
rect 142462 160378 159906 160614
rect 160142 160378 160226 160614
rect 160462 160378 177906 160614
rect 178142 160378 178226 160614
rect 178462 160378 195906 160614
rect 196142 160378 196226 160614
rect 196462 160378 213906 160614
rect 214142 160378 214226 160614
rect 214462 160378 231906 160614
rect 232142 160378 232226 160614
rect 232462 160378 249906 160614
rect 250142 160378 250226 160614
rect 250462 160378 267906 160614
rect 268142 160378 268226 160614
rect 268462 160378 285906 160614
rect 286142 160378 286226 160614
rect 286462 160378 303906 160614
rect 304142 160378 304226 160614
rect 304462 160378 321906 160614
rect 322142 160378 322226 160614
rect 322462 160378 339906 160614
rect 340142 160378 340226 160614
rect 340462 160378 357906 160614
rect 358142 160378 358226 160614
rect 358462 160378 375906 160614
rect 376142 160378 376226 160614
rect 376462 160378 393906 160614
rect 394142 160378 394226 160614
rect 394462 160378 411906 160614
rect 412142 160378 412226 160614
rect 412462 160378 429906 160614
rect 430142 160378 430226 160614
rect 430462 160378 447906 160614
rect 448142 160378 448226 160614
rect 448462 160378 465906 160614
rect 466142 160378 466226 160614
rect 466462 160378 483906 160614
rect 484142 160378 484226 160614
rect 484462 160378 501906 160614
rect 502142 160378 502226 160614
rect 502462 160378 519906 160614
rect 520142 160378 520226 160614
rect 520462 160378 537906 160614
rect 538142 160378 538226 160614
rect 538462 160378 547884 160614
rect 548120 160378 548204 160614
rect 548440 160378 548472 160614
rect -4476 160294 548472 160378
rect -4476 160058 -4444 160294
rect -4208 160058 -4124 160294
rect -3888 160058 15906 160294
rect 16142 160058 16226 160294
rect 16462 160058 33906 160294
rect 34142 160058 34226 160294
rect 34462 160058 51906 160294
rect 52142 160058 52226 160294
rect 52462 160058 69906 160294
rect 70142 160058 70226 160294
rect 70462 160058 87906 160294
rect 88142 160058 88226 160294
rect 88462 160058 105906 160294
rect 106142 160058 106226 160294
rect 106462 160058 123906 160294
rect 124142 160058 124226 160294
rect 124462 160058 141906 160294
rect 142142 160058 142226 160294
rect 142462 160058 159906 160294
rect 160142 160058 160226 160294
rect 160462 160058 177906 160294
rect 178142 160058 178226 160294
rect 178462 160058 195906 160294
rect 196142 160058 196226 160294
rect 196462 160058 213906 160294
rect 214142 160058 214226 160294
rect 214462 160058 231906 160294
rect 232142 160058 232226 160294
rect 232462 160058 249906 160294
rect 250142 160058 250226 160294
rect 250462 160058 267906 160294
rect 268142 160058 268226 160294
rect 268462 160058 285906 160294
rect 286142 160058 286226 160294
rect 286462 160058 303906 160294
rect 304142 160058 304226 160294
rect 304462 160058 321906 160294
rect 322142 160058 322226 160294
rect 322462 160058 339906 160294
rect 340142 160058 340226 160294
rect 340462 160058 357906 160294
rect 358142 160058 358226 160294
rect 358462 160058 375906 160294
rect 376142 160058 376226 160294
rect 376462 160058 393906 160294
rect 394142 160058 394226 160294
rect 394462 160058 411906 160294
rect 412142 160058 412226 160294
rect 412462 160058 429906 160294
rect 430142 160058 430226 160294
rect 430462 160058 447906 160294
rect 448142 160058 448226 160294
rect 448462 160058 465906 160294
rect 466142 160058 466226 160294
rect 466462 160058 483906 160294
rect 484142 160058 484226 160294
rect 484462 160058 501906 160294
rect 502142 160058 502226 160294
rect 502462 160058 519906 160294
rect 520142 160058 520226 160294
rect 520462 160058 537906 160294
rect 538142 160058 538226 160294
rect 538462 160058 547884 160294
rect 548120 160058 548204 160294
rect 548440 160058 548472 160294
rect -4476 160026 548472 160058
rect -4476 156894 548472 156926
rect -4476 156658 -3484 156894
rect -3248 156658 -3164 156894
rect -2928 156658 12186 156894
rect 12422 156658 12506 156894
rect 12742 156658 30186 156894
rect 30422 156658 30506 156894
rect 30742 156658 48186 156894
rect 48422 156658 48506 156894
rect 48742 156658 66186 156894
rect 66422 156658 66506 156894
rect 66742 156658 84186 156894
rect 84422 156658 84506 156894
rect 84742 156658 102186 156894
rect 102422 156658 102506 156894
rect 102742 156658 120186 156894
rect 120422 156658 120506 156894
rect 120742 156658 138186 156894
rect 138422 156658 138506 156894
rect 138742 156658 156186 156894
rect 156422 156658 156506 156894
rect 156742 156658 174186 156894
rect 174422 156658 174506 156894
rect 174742 156658 192186 156894
rect 192422 156658 192506 156894
rect 192742 156658 210186 156894
rect 210422 156658 210506 156894
rect 210742 156658 228186 156894
rect 228422 156658 228506 156894
rect 228742 156658 246186 156894
rect 246422 156658 246506 156894
rect 246742 156658 264186 156894
rect 264422 156658 264506 156894
rect 264742 156658 282186 156894
rect 282422 156658 282506 156894
rect 282742 156658 300186 156894
rect 300422 156658 300506 156894
rect 300742 156658 318186 156894
rect 318422 156658 318506 156894
rect 318742 156658 336186 156894
rect 336422 156658 336506 156894
rect 336742 156658 354186 156894
rect 354422 156658 354506 156894
rect 354742 156658 372186 156894
rect 372422 156658 372506 156894
rect 372742 156658 390186 156894
rect 390422 156658 390506 156894
rect 390742 156658 408186 156894
rect 408422 156658 408506 156894
rect 408742 156658 426186 156894
rect 426422 156658 426506 156894
rect 426742 156658 444186 156894
rect 444422 156658 444506 156894
rect 444742 156658 462186 156894
rect 462422 156658 462506 156894
rect 462742 156658 480186 156894
rect 480422 156658 480506 156894
rect 480742 156658 498186 156894
rect 498422 156658 498506 156894
rect 498742 156658 516186 156894
rect 516422 156658 516506 156894
rect 516742 156658 534186 156894
rect 534422 156658 534506 156894
rect 534742 156658 546924 156894
rect 547160 156658 547244 156894
rect 547480 156658 548472 156894
rect -4476 156574 548472 156658
rect -4476 156338 -3484 156574
rect -3248 156338 -3164 156574
rect -2928 156338 12186 156574
rect 12422 156338 12506 156574
rect 12742 156338 30186 156574
rect 30422 156338 30506 156574
rect 30742 156338 48186 156574
rect 48422 156338 48506 156574
rect 48742 156338 66186 156574
rect 66422 156338 66506 156574
rect 66742 156338 84186 156574
rect 84422 156338 84506 156574
rect 84742 156338 102186 156574
rect 102422 156338 102506 156574
rect 102742 156338 120186 156574
rect 120422 156338 120506 156574
rect 120742 156338 138186 156574
rect 138422 156338 138506 156574
rect 138742 156338 156186 156574
rect 156422 156338 156506 156574
rect 156742 156338 174186 156574
rect 174422 156338 174506 156574
rect 174742 156338 192186 156574
rect 192422 156338 192506 156574
rect 192742 156338 210186 156574
rect 210422 156338 210506 156574
rect 210742 156338 228186 156574
rect 228422 156338 228506 156574
rect 228742 156338 246186 156574
rect 246422 156338 246506 156574
rect 246742 156338 264186 156574
rect 264422 156338 264506 156574
rect 264742 156338 282186 156574
rect 282422 156338 282506 156574
rect 282742 156338 300186 156574
rect 300422 156338 300506 156574
rect 300742 156338 318186 156574
rect 318422 156338 318506 156574
rect 318742 156338 336186 156574
rect 336422 156338 336506 156574
rect 336742 156338 354186 156574
rect 354422 156338 354506 156574
rect 354742 156338 372186 156574
rect 372422 156338 372506 156574
rect 372742 156338 390186 156574
rect 390422 156338 390506 156574
rect 390742 156338 408186 156574
rect 408422 156338 408506 156574
rect 408742 156338 426186 156574
rect 426422 156338 426506 156574
rect 426742 156338 444186 156574
rect 444422 156338 444506 156574
rect 444742 156338 462186 156574
rect 462422 156338 462506 156574
rect 462742 156338 480186 156574
rect 480422 156338 480506 156574
rect 480742 156338 498186 156574
rect 498422 156338 498506 156574
rect 498742 156338 516186 156574
rect 516422 156338 516506 156574
rect 516742 156338 534186 156574
rect 534422 156338 534506 156574
rect 534742 156338 546924 156574
rect 547160 156338 547244 156574
rect 547480 156338 548472 156574
rect -4476 156306 548472 156338
rect -4476 153174 548472 153206
rect -4476 152938 -2524 153174
rect -2288 152938 -2204 153174
rect -1968 152938 8466 153174
rect 8702 152938 8786 153174
rect 9022 152938 26466 153174
rect 26702 152938 26786 153174
rect 27022 152938 44466 153174
rect 44702 152938 44786 153174
rect 45022 152938 62466 153174
rect 62702 152938 62786 153174
rect 63022 152938 80466 153174
rect 80702 152938 80786 153174
rect 81022 152938 98466 153174
rect 98702 152938 98786 153174
rect 99022 152938 116466 153174
rect 116702 152938 116786 153174
rect 117022 152938 134466 153174
rect 134702 152938 134786 153174
rect 135022 152938 152466 153174
rect 152702 152938 152786 153174
rect 153022 152938 170466 153174
rect 170702 152938 170786 153174
rect 171022 152938 188466 153174
rect 188702 152938 188786 153174
rect 189022 152938 206466 153174
rect 206702 152938 206786 153174
rect 207022 152938 224466 153174
rect 224702 152938 224786 153174
rect 225022 152938 242466 153174
rect 242702 152938 242786 153174
rect 243022 152938 260466 153174
rect 260702 152938 260786 153174
rect 261022 152938 278466 153174
rect 278702 152938 278786 153174
rect 279022 152938 296466 153174
rect 296702 152938 296786 153174
rect 297022 152938 314466 153174
rect 314702 152938 314786 153174
rect 315022 152938 332466 153174
rect 332702 152938 332786 153174
rect 333022 152938 350466 153174
rect 350702 152938 350786 153174
rect 351022 152938 368466 153174
rect 368702 152938 368786 153174
rect 369022 152938 386466 153174
rect 386702 152938 386786 153174
rect 387022 152938 404466 153174
rect 404702 152938 404786 153174
rect 405022 152938 422466 153174
rect 422702 152938 422786 153174
rect 423022 152938 440466 153174
rect 440702 152938 440786 153174
rect 441022 152938 458466 153174
rect 458702 152938 458786 153174
rect 459022 152938 476466 153174
rect 476702 152938 476786 153174
rect 477022 152938 494466 153174
rect 494702 152938 494786 153174
rect 495022 152938 512466 153174
rect 512702 152938 512786 153174
rect 513022 152938 530466 153174
rect 530702 152938 530786 153174
rect 531022 152938 545964 153174
rect 546200 152938 546284 153174
rect 546520 152938 548472 153174
rect -4476 152854 548472 152938
rect -4476 152618 -2524 152854
rect -2288 152618 -2204 152854
rect -1968 152618 8466 152854
rect 8702 152618 8786 152854
rect 9022 152618 26466 152854
rect 26702 152618 26786 152854
rect 27022 152618 44466 152854
rect 44702 152618 44786 152854
rect 45022 152618 62466 152854
rect 62702 152618 62786 152854
rect 63022 152618 80466 152854
rect 80702 152618 80786 152854
rect 81022 152618 98466 152854
rect 98702 152618 98786 152854
rect 99022 152618 116466 152854
rect 116702 152618 116786 152854
rect 117022 152618 134466 152854
rect 134702 152618 134786 152854
rect 135022 152618 152466 152854
rect 152702 152618 152786 152854
rect 153022 152618 170466 152854
rect 170702 152618 170786 152854
rect 171022 152618 188466 152854
rect 188702 152618 188786 152854
rect 189022 152618 206466 152854
rect 206702 152618 206786 152854
rect 207022 152618 224466 152854
rect 224702 152618 224786 152854
rect 225022 152618 242466 152854
rect 242702 152618 242786 152854
rect 243022 152618 260466 152854
rect 260702 152618 260786 152854
rect 261022 152618 278466 152854
rect 278702 152618 278786 152854
rect 279022 152618 296466 152854
rect 296702 152618 296786 152854
rect 297022 152618 314466 152854
rect 314702 152618 314786 152854
rect 315022 152618 332466 152854
rect 332702 152618 332786 152854
rect 333022 152618 350466 152854
rect 350702 152618 350786 152854
rect 351022 152618 368466 152854
rect 368702 152618 368786 152854
rect 369022 152618 386466 152854
rect 386702 152618 386786 152854
rect 387022 152618 404466 152854
rect 404702 152618 404786 152854
rect 405022 152618 422466 152854
rect 422702 152618 422786 152854
rect 423022 152618 440466 152854
rect 440702 152618 440786 152854
rect 441022 152618 458466 152854
rect 458702 152618 458786 152854
rect 459022 152618 476466 152854
rect 476702 152618 476786 152854
rect 477022 152618 494466 152854
rect 494702 152618 494786 152854
rect 495022 152618 512466 152854
rect 512702 152618 512786 152854
rect 513022 152618 530466 152854
rect 530702 152618 530786 152854
rect 531022 152618 545964 152854
rect 546200 152618 546284 152854
rect 546520 152618 548472 152854
rect -4476 152586 548472 152618
rect -4476 149454 548472 149486
rect -4476 149218 -1564 149454
rect -1328 149218 -1244 149454
rect -1008 149218 4746 149454
rect 4982 149218 5066 149454
rect 5302 149218 22746 149454
rect 22982 149218 23066 149454
rect 23302 149218 40746 149454
rect 40982 149218 41066 149454
rect 41302 149218 58746 149454
rect 58982 149218 59066 149454
rect 59302 149218 76746 149454
rect 76982 149218 77066 149454
rect 77302 149218 94746 149454
rect 94982 149218 95066 149454
rect 95302 149218 112746 149454
rect 112982 149218 113066 149454
rect 113302 149218 130746 149454
rect 130982 149218 131066 149454
rect 131302 149218 148746 149454
rect 148982 149218 149066 149454
rect 149302 149218 166746 149454
rect 166982 149218 167066 149454
rect 167302 149218 184746 149454
rect 184982 149218 185066 149454
rect 185302 149218 202746 149454
rect 202982 149218 203066 149454
rect 203302 149218 220746 149454
rect 220982 149218 221066 149454
rect 221302 149218 238746 149454
rect 238982 149218 239066 149454
rect 239302 149218 256746 149454
rect 256982 149218 257066 149454
rect 257302 149218 274746 149454
rect 274982 149218 275066 149454
rect 275302 149218 292746 149454
rect 292982 149218 293066 149454
rect 293302 149218 310746 149454
rect 310982 149218 311066 149454
rect 311302 149218 328746 149454
rect 328982 149218 329066 149454
rect 329302 149218 346746 149454
rect 346982 149218 347066 149454
rect 347302 149218 364746 149454
rect 364982 149218 365066 149454
rect 365302 149218 382746 149454
rect 382982 149218 383066 149454
rect 383302 149218 400746 149454
rect 400982 149218 401066 149454
rect 401302 149218 418746 149454
rect 418982 149218 419066 149454
rect 419302 149218 436746 149454
rect 436982 149218 437066 149454
rect 437302 149218 454746 149454
rect 454982 149218 455066 149454
rect 455302 149218 472746 149454
rect 472982 149218 473066 149454
rect 473302 149218 490746 149454
rect 490982 149218 491066 149454
rect 491302 149218 508746 149454
rect 508982 149218 509066 149454
rect 509302 149218 526746 149454
rect 526982 149218 527066 149454
rect 527302 149218 545004 149454
rect 545240 149218 545324 149454
rect 545560 149218 548472 149454
rect -4476 149134 548472 149218
rect -4476 148898 -1564 149134
rect -1328 148898 -1244 149134
rect -1008 148898 4746 149134
rect 4982 148898 5066 149134
rect 5302 148898 22746 149134
rect 22982 148898 23066 149134
rect 23302 148898 40746 149134
rect 40982 148898 41066 149134
rect 41302 148898 58746 149134
rect 58982 148898 59066 149134
rect 59302 148898 76746 149134
rect 76982 148898 77066 149134
rect 77302 148898 94746 149134
rect 94982 148898 95066 149134
rect 95302 148898 112746 149134
rect 112982 148898 113066 149134
rect 113302 148898 130746 149134
rect 130982 148898 131066 149134
rect 131302 148898 148746 149134
rect 148982 148898 149066 149134
rect 149302 148898 166746 149134
rect 166982 148898 167066 149134
rect 167302 148898 184746 149134
rect 184982 148898 185066 149134
rect 185302 148898 202746 149134
rect 202982 148898 203066 149134
rect 203302 148898 220746 149134
rect 220982 148898 221066 149134
rect 221302 148898 238746 149134
rect 238982 148898 239066 149134
rect 239302 148898 256746 149134
rect 256982 148898 257066 149134
rect 257302 148898 274746 149134
rect 274982 148898 275066 149134
rect 275302 148898 292746 149134
rect 292982 148898 293066 149134
rect 293302 148898 310746 149134
rect 310982 148898 311066 149134
rect 311302 148898 328746 149134
rect 328982 148898 329066 149134
rect 329302 148898 346746 149134
rect 346982 148898 347066 149134
rect 347302 148898 364746 149134
rect 364982 148898 365066 149134
rect 365302 148898 382746 149134
rect 382982 148898 383066 149134
rect 383302 148898 400746 149134
rect 400982 148898 401066 149134
rect 401302 148898 418746 149134
rect 418982 148898 419066 149134
rect 419302 148898 436746 149134
rect 436982 148898 437066 149134
rect 437302 148898 454746 149134
rect 454982 148898 455066 149134
rect 455302 148898 472746 149134
rect 472982 148898 473066 149134
rect 473302 148898 490746 149134
rect 490982 148898 491066 149134
rect 491302 148898 508746 149134
rect 508982 148898 509066 149134
rect 509302 148898 526746 149134
rect 526982 148898 527066 149134
rect 527302 148898 545004 149134
rect 545240 148898 545324 149134
rect 545560 148898 548472 149134
rect -4476 148866 548472 148898
rect -4476 142614 548472 142646
rect -4476 142378 -4444 142614
rect -4208 142378 -4124 142614
rect -3888 142378 15906 142614
rect 16142 142378 16226 142614
rect 16462 142378 33906 142614
rect 34142 142378 34226 142614
rect 34462 142378 51906 142614
rect 52142 142378 52226 142614
rect 52462 142378 69906 142614
rect 70142 142378 70226 142614
rect 70462 142378 87906 142614
rect 88142 142378 88226 142614
rect 88462 142378 105906 142614
rect 106142 142378 106226 142614
rect 106462 142378 123906 142614
rect 124142 142378 124226 142614
rect 124462 142378 141906 142614
rect 142142 142378 142226 142614
rect 142462 142378 159906 142614
rect 160142 142378 160226 142614
rect 160462 142378 177906 142614
rect 178142 142378 178226 142614
rect 178462 142378 195906 142614
rect 196142 142378 196226 142614
rect 196462 142378 213906 142614
rect 214142 142378 214226 142614
rect 214462 142378 231906 142614
rect 232142 142378 232226 142614
rect 232462 142378 249906 142614
rect 250142 142378 250226 142614
rect 250462 142378 267906 142614
rect 268142 142378 268226 142614
rect 268462 142378 285906 142614
rect 286142 142378 286226 142614
rect 286462 142378 303906 142614
rect 304142 142378 304226 142614
rect 304462 142378 321906 142614
rect 322142 142378 322226 142614
rect 322462 142378 339906 142614
rect 340142 142378 340226 142614
rect 340462 142378 357906 142614
rect 358142 142378 358226 142614
rect 358462 142378 375906 142614
rect 376142 142378 376226 142614
rect 376462 142378 393906 142614
rect 394142 142378 394226 142614
rect 394462 142378 411906 142614
rect 412142 142378 412226 142614
rect 412462 142378 429906 142614
rect 430142 142378 430226 142614
rect 430462 142378 447906 142614
rect 448142 142378 448226 142614
rect 448462 142378 465906 142614
rect 466142 142378 466226 142614
rect 466462 142378 483906 142614
rect 484142 142378 484226 142614
rect 484462 142378 501906 142614
rect 502142 142378 502226 142614
rect 502462 142378 519906 142614
rect 520142 142378 520226 142614
rect 520462 142378 537906 142614
rect 538142 142378 538226 142614
rect 538462 142378 547884 142614
rect 548120 142378 548204 142614
rect 548440 142378 548472 142614
rect -4476 142294 548472 142378
rect -4476 142058 -4444 142294
rect -4208 142058 -4124 142294
rect -3888 142058 15906 142294
rect 16142 142058 16226 142294
rect 16462 142058 33906 142294
rect 34142 142058 34226 142294
rect 34462 142058 51906 142294
rect 52142 142058 52226 142294
rect 52462 142058 69906 142294
rect 70142 142058 70226 142294
rect 70462 142058 87906 142294
rect 88142 142058 88226 142294
rect 88462 142058 105906 142294
rect 106142 142058 106226 142294
rect 106462 142058 123906 142294
rect 124142 142058 124226 142294
rect 124462 142058 141906 142294
rect 142142 142058 142226 142294
rect 142462 142058 159906 142294
rect 160142 142058 160226 142294
rect 160462 142058 177906 142294
rect 178142 142058 178226 142294
rect 178462 142058 195906 142294
rect 196142 142058 196226 142294
rect 196462 142058 213906 142294
rect 214142 142058 214226 142294
rect 214462 142058 231906 142294
rect 232142 142058 232226 142294
rect 232462 142058 249906 142294
rect 250142 142058 250226 142294
rect 250462 142058 267906 142294
rect 268142 142058 268226 142294
rect 268462 142058 285906 142294
rect 286142 142058 286226 142294
rect 286462 142058 303906 142294
rect 304142 142058 304226 142294
rect 304462 142058 321906 142294
rect 322142 142058 322226 142294
rect 322462 142058 339906 142294
rect 340142 142058 340226 142294
rect 340462 142058 357906 142294
rect 358142 142058 358226 142294
rect 358462 142058 375906 142294
rect 376142 142058 376226 142294
rect 376462 142058 393906 142294
rect 394142 142058 394226 142294
rect 394462 142058 411906 142294
rect 412142 142058 412226 142294
rect 412462 142058 429906 142294
rect 430142 142058 430226 142294
rect 430462 142058 447906 142294
rect 448142 142058 448226 142294
rect 448462 142058 465906 142294
rect 466142 142058 466226 142294
rect 466462 142058 483906 142294
rect 484142 142058 484226 142294
rect 484462 142058 501906 142294
rect 502142 142058 502226 142294
rect 502462 142058 519906 142294
rect 520142 142058 520226 142294
rect 520462 142058 537906 142294
rect 538142 142058 538226 142294
rect 538462 142058 547884 142294
rect 548120 142058 548204 142294
rect 548440 142058 548472 142294
rect -4476 142026 548472 142058
rect -4476 138894 548472 138926
rect -4476 138658 -3484 138894
rect -3248 138658 -3164 138894
rect -2928 138658 12186 138894
rect 12422 138658 12506 138894
rect 12742 138658 30186 138894
rect 30422 138658 30506 138894
rect 30742 138658 48186 138894
rect 48422 138658 48506 138894
rect 48742 138658 66186 138894
rect 66422 138658 66506 138894
rect 66742 138658 84186 138894
rect 84422 138658 84506 138894
rect 84742 138658 102186 138894
rect 102422 138658 102506 138894
rect 102742 138658 120186 138894
rect 120422 138658 120506 138894
rect 120742 138658 138186 138894
rect 138422 138658 138506 138894
rect 138742 138658 156186 138894
rect 156422 138658 156506 138894
rect 156742 138658 174186 138894
rect 174422 138658 174506 138894
rect 174742 138658 192186 138894
rect 192422 138658 192506 138894
rect 192742 138658 210186 138894
rect 210422 138658 210506 138894
rect 210742 138658 228186 138894
rect 228422 138658 228506 138894
rect 228742 138658 246186 138894
rect 246422 138658 246506 138894
rect 246742 138658 264186 138894
rect 264422 138658 264506 138894
rect 264742 138658 282186 138894
rect 282422 138658 282506 138894
rect 282742 138658 300186 138894
rect 300422 138658 300506 138894
rect 300742 138658 318186 138894
rect 318422 138658 318506 138894
rect 318742 138658 336186 138894
rect 336422 138658 336506 138894
rect 336742 138658 354186 138894
rect 354422 138658 354506 138894
rect 354742 138658 372186 138894
rect 372422 138658 372506 138894
rect 372742 138658 390186 138894
rect 390422 138658 390506 138894
rect 390742 138658 408186 138894
rect 408422 138658 408506 138894
rect 408742 138658 426186 138894
rect 426422 138658 426506 138894
rect 426742 138658 444186 138894
rect 444422 138658 444506 138894
rect 444742 138658 462186 138894
rect 462422 138658 462506 138894
rect 462742 138658 480186 138894
rect 480422 138658 480506 138894
rect 480742 138658 498186 138894
rect 498422 138658 498506 138894
rect 498742 138658 516186 138894
rect 516422 138658 516506 138894
rect 516742 138658 534186 138894
rect 534422 138658 534506 138894
rect 534742 138658 546924 138894
rect 547160 138658 547244 138894
rect 547480 138658 548472 138894
rect -4476 138574 548472 138658
rect -4476 138338 -3484 138574
rect -3248 138338 -3164 138574
rect -2928 138338 12186 138574
rect 12422 138338 12506 138574
rect 12742 138338 30186 138574
rect 30422 138338 30506 138574
rect 30742 138338 48186 138574
rect 48422 138338 48506 138574
rect 48742 138338 66186 138574
rect 66422 138338 66506 138574
rect 66742 138338 84186 138574
rect 84422 138338 84506 138574
rect 84742 138338 102186 138574
rect 102422 138338 102506 138574
rect 102742 138338 120186 138574
rect 120422 138338 120506 138574
rect 120742 138338 138186 138574
rect 138422 138338 138506 138574
rect 138742 138338 156186 138574
rect 156422 138338 156506 138574
rect 156742 138338 174186 138574
rect 174422 138338 174506 138574
rect 174742 138338 192186 138574
rect 192422 138338 192506 138574
rect 192742 138338 210186 138574
rect 210422 138338 210506 138574
rect 210742 138338 228186 138574
rect 228422 138338 228506 138574
rect 228742 138338 246186 138574
rect 246422 138338 246506 138574
rect 246742 138338 264186 138574
rect 264422 138338 264506 138574
rect 264742 138338 282186 138574
rect 282422 138338 282506 138574
rect 282742 138338 300186 138574
rect 300422 138338 300506 138574
rect 300742 138338 318186 138574
rect 318422 138338 318506 138574
rect 318742 138338 336186 138574
rect 336422 138338 336506 138574
rect 336742 138338 354186 138574
rect 354422 138338 354506 138574
rect 354742 138338 372186 138574
rect 372422 138338 372506 138574
rect 372742 138338 390186 138574
rect 390422 138338 390506 138574
rect 390742 138338 408186 138574
rect 408422 138338 408506 138574
rect 408742 138338 426186 138574
rect 426422 138338 426506 138574
rect 426742 138338 444186 138574
rect 444422 138338 444506 138574
rect 444742 138338 462186 138574
rect 462422 138338 462506 138574
rect 462742 138338 480186 138574
rect 480422 138338 480506 138574
rect 480742 138338 498186 138574
rect 498422 138338 498506 138574
rect 498742 138338 516186 138574
rect 516422 138338 516506 138574
rect 516742 138338 534186 138574
rect 534422 138338 534506 138574
rect 534742 138338 546924 138574
rect 547160 138338 547244 138574
rect 547480 138338 548472 138574
rect -4476 138306 548472 138338
rect -4476 135174 548472 135206
rect -4476 134938 -2524 135174
rect -2288 134938 -2204 135174
rect -1968 134938 8466 135174
rect 8702 134938 8786 135174
rect 9022 134938 26466 135174
rect 26702 134938 26786 135174
rect 27022 134938 44466 135174
rect 44702 134938 44786 135174
rect 45022 134938 62466 135174
rect 62702 134938 62786 135174
rect 63022 134938 80466 135174
rect 80702 134938 80786 135174
rect 81022 134938 98466 135174
rect 98702 134938 98786 135174
rect 99022 134938 116466 135174
rect 116702 134938 116786 135174
rect 117022 134938 134466 135174
rect 134702 134938 134786 135174
rect 135022 134938 152466 135174
rect 152702 134938 152786 135174
rect 153022 134938 170466 135174
rect 170702 134938 170786 135174
rect 171022 134938 188466 135174
rect 188702 134938 188786 135174
rect 189022 134938 206466 135174
rect 206702 134938 206786 135174
rect 207022 134938 224466 135174
rect 224702 134938 224786 135174
rect 225022 134938 242466 135174
rect 242702 134938 242786 135174
rect 243022 134938 260466 135174
rect 260702 134938 260786 135174
rect 261022 134938 278466 135174
rect 278702 134938 278786 135174
rect 279022 134938 296466 135174
rect 296702 134938 296786 135174
rect 297022 134938 314466 135174
rect 314702 134938 314786 135174
rect 315022 134938 332466 135174
rect 332702 134938 332786 135174
rect 333022 134938 350466 135174
rect 350702 134938 350786 135174
rect 351022 134938 368466 135174
rect 368702 134938 368786 135174
rect 369022 134938 386466 135174
rect 386702 134938 386786 135174
rect 387022 134938 404466 135174
rect 404702 134938 404786 135174
rect 405022 134938 422466 135174
rect 422702 134938 422786 135174
rect 423022 134938 440466 135174
rect 440702 134938 440786 135174
rect 441022 134938 458466 135174
rect 458702 134938 458786 135174
rect 459022 134938 476466 135174
rect 476702 134938 476786 135174
rect 477022 134938 494466 135174
rect 494702 134938 494786 135174
rect 495022 134938 512466 135174
rect 512702 134938 512786 135174
rect 513022 134938 530466 135174
rect 530702 134938 530786 135174
rect 531022 134938 545964 135174
rect 546200 134938 546284 135174
rect 546520 134938 548472 135174
rect -4476 134854 548472 134938
rect -4476 134618 -2524 134854
rect -2288 134618 -2204 134854
rect -1968 134618 8466 134854
rect 8702 134618 8786 134854
rect 9022 134618 26466 134854
rect 26702 134618 26786 134854
rect 27022 134618 44466 134854
rect 44702 134618 44786 134854
rect 45022 134618 62466 134854
rect 62702 134618 62786 134854
rect 63022 134618 80466 134854
rect 80702 134618 80786 134854
rect 81022 134618 98466 134854
rect 98702 134618 98786 134854
rect 99022 134618 116466 134854
rect 116702 134618 116786 134854
rect 117022 134618 134466 134854
rect 134702 134618 134786 134854
rect 135022 134618 152466 134854
rect 152702 134618 152786 134854
rect 153022 134618 170466 134854
rect 170702 134618 170786 134854
rect 171022 134618 188466 134854
rect 188702 134618 188786 134854
rect 189022 134618 206466 134854
rect 206702 134618 206786 134854
rect 207022 134618 224466 134854
rect 224702 134618 224786 134854
rect 225022 134618 242466 134854
rect 242702 134618 242786 134854
rect 243022 134618 260466 134854
rect 260702 134618 260786 134854
rect 261022 134618 278466 134854
rect 278702 134618 278786 134854
rect 279022 134618 296466 134854
rect 296702 134618 296786 134854
rect 297022 134618 314466 134854
rect 314702 134618 314786 134854
rect 315022 134618 332466 134854
rect 332702 134618 332786 134854
rect 333022 134618 350466 134854
rect 350702 134618 350786 134854
rect 351022 134618 368466 134854
rect 368702 134618 368786 134854
rect 369022 134618 386466 134854
rect 386702 134618 386786 134854
rect 387022 134618 404466 134854
rect 404702 134618 404786 134854
rect 405022 134618 422466 134854
rect 422702 134618 422786 134854
rect 423022 134618 440466 134854
rect 440702 134618 440786 134854
rect 441022 134618 458466 134854
rect 458702 134618 458786 134854
rect 459022 134618 476466 134854
rect 476702 134618 476786 134854
rect 477022 134618 494466 134854
rect 494702 134618 494786 134854
rect 495022 134618 512466 134854
rect 512702 134618 512786 134854
rect 513022 134618 530466 134854
rect 530702 134618 530786 134854
rect 531022 134618 545964 134854
rect 546200 134618 546284 134854
rect 546520 134618 548472 134854
rect -4476 134586 548472 134618
rect -4476 131454 548472 131486
rect -4476 131218 -1564 131454
rect -1328 131218 -1244 131454
rect -1008 131218 4746 131454
rect 4982 131218 5066 131454
rect 5302 131218 22746 131454
rect 22982 131218 23066 131454
rect 23302 131218 40746 131454
rect 40982 131218 41066 131454
rect 41302 131218 58746 131454
rect 58982 131218 59066 131454
rect 59302 131218 76746 131454
rect 76982 131218 77066 131454
rect 77302 131218 94746 131454
rect 94982 131218 95066 131454
rect 95302 131218 112746 131454
rect 112982 131218 113066 131454
rect 113302 131218 130746 131454
rect 130982 131218 131066 131454
rect 131302 131218 148746 131454
rect 148982 131218 149066 131454
rect 149302 131218 166746 131454
rect 166982 131218 167066 131454
rect 167302 131218 184746 131454
rect 184982 131218 185066 131454
rect 185302 131218 202746 131454
rect 202982 131218 203066 131454
rect 203302 131218 220746 131454
rect 220982 131218 221066 131454
rect 221302 131218 238746 131454
rect 238982 131218 239066 131454
rect 239302 131218 256746 131454
rect 256982 131218 257066 131454
rect 257302 131218 274746 131454
rect 274982 131218 275066 131454
rect 275302 131218 292746 131454
rect 292982 131218 293066 131454
rect 293302 131218 310746 131454
rect 310982 131218 311066 131454
rect 311302 131218 328746 131454
rect 328982 131218 329066 131454
rect 329302 131218 346746 131454
rect 346982 131218 347066 131454
rect 347302 131218 364746 131454
rect 364982 131218 365066 131454
rect 365302 131218 382746 131454
rect 382982 131218 383066 131454
rect 383302 131218 400746 131454
rect 400982 131218 401066 131454
rect 401302 131218 418746 131454
rect 418982 131218 419066 131454
rect 419302 131218 436746 131454
rect 436982 131218 437066 131454
rect 437302 131218 454746 131454
rect 454982 131218 455066 131454
rect 455302 131218 472746 131454
rect 472982 131218 473066 131454
rect 473302 131218 490746 131454
rect 490982 131218 491066 131454
rect 491302 131218 508746 131454
rect 508982 131218 509066 131454
rect 509302 131218 526746 131454
rect 526982 131218 527066 131454
rect 527302 131218 545004 131454
rect 545240 131218 545324 131454
rect 545560 131218 548472 131454
rect -4476 131134 548472 131218
rect -4476 130898 -1564 131134
rect -1328 130898 -1244 131134
rect -1008 130898 4746 131134
rect 4982 130898 5066 131134
rect 5302 130898 22746 131134
rect 22982 130898 23066 131134
rect 23302 130898 40746 131134
rect 40982 130898 41066 131134
rect 41302 130898 58746 131134
rect 58982 130898 59066 131134
rect 59302 130898 76746 131134
rect 76982 130898 77066 131134
rect 77302 130898 94746 131134
rect 94982 130898 95066 131134
rect 95302 130898 112746 131134
rect 112982 130898 113066 131134
rect 113302 130898 130746 131134
rect 130982 130898 131066 131134
rect 131302 130898 148746 131134
rect 148982 130898 149066 131134
rect 149302 130898 166746 131134
rect 166982 130898 167066 131134
rect 167302 130898 184746 131134
rect 184982 130898 185066 131134
rect 185302 130898 202746 131134
rect 202982 130898 203066 131134
rect 203302 130898 220746 131134
rect 220982 130898 221066 131134
rect 221302 130898 238746 131134
rect 238982 130898 239066 131134
rect 239302 130898 256746 131134
rect 256982 130898 257066 131134
rect 257302 130898 274746 131134
rect 274982 130898 275066 131134
rect 275302 130898 292746 131134
rect 292982 130898 293066 131134
rect 293302 130898 310746 131134
rect 310982 130898 311066 131134
rect 311302 130898 328746 131134
rect 328982 130898 329066 131134
rect 329302 130898 346746 131134
rect 346982 130898 347066 131134
rect 347302 130898 364746 131134
rect 364982 130898 365066 131134
rect 365302 130898 382746 131134
rect 382982 130898 383066 131134
rect 383302 130898 400746 131134
rect 400982 130898 401066 131134
rect 401302 130898 418746 131134
rect 418982 130898 419066 131134
rect 419302 130898 436746 131134
rect 436982 130898 437066 131134
rect 437302 130898 454746 131134
rect 454982 130898 455066 131134
rect 455302 130898 472746 131134
rect 472982 130898 473066 131134
rect 473302 130898 490746 131134
rect 490982 130898 491066 131134
rect 491302 130898 508746 131134
rect 508982 130898 509066 131134
rect 509302 130898 526746 131134
rect 526982 130898 527066 131134
rect 527302 130898 545004 131134
rect 545240 130898 545324 131134
rect 545560 130898 548472 131134
rect -4476 130866 548472 130898
rect -4476 124614 548472 124646
rect -4476 124378 -4444 124614
rect -4208 124378 -4124 124614
rect -3888 124378 15906 124614
rect 16142 124378 16226 124614
rect 16462 124378 33906 124614
rect 34142 124378 34226 124614
rect 34462 124378 51906 124614
rect 52142 124378 52226 124614
rect 52462 124378 69906 124614
rect 70142 124378 70226 124614
rect 70462 124378 87906 124614
rect 88142 124378 88226 124614
rect 88462 124378 105906 124614
rect 106142 124378 106226 124614
rect 106462 124378 123906 124614
rect 124142 124378 124226 124614
rect 124462 124378 141906 124614
rect 142142 124378 142226 124614
rect 142462 124378 159906 124614
rect 160142 124378 160226 124614
rect 160462 124378 177906 124614
rect 178142 124378 178226 124614
rect 178462 124378 195906 124614
rect 196142 124378 196226 124614
rect 196462 124378 213906 124614
rect 214142 124378 214226 124614
rect 214462 124378 231906 124614
rect 232142 124378 232226 124614
rect 232462 124378 249906 124614
rect 250142 124378 250226 124614
rect 250462 124378 267906 124614
rect 268142 124378 268226 124614
rect 268462 124378 285906 124614
rect 286142 124378 286226 124614
rect 286462 124378 303906 124614
rect 304142 124378 304226 124614
rect 304462 124378 321906 124614
rect 322142 124378 322226 124614
rect 322462 124378 339906 124614
rect 340142 124378 340226 124614
rect 340462 124378 357906 124614
rect 358142 124378 358226 124614
rect 358462 124378 375906 124614
rect 376142 124378 376226 124614
rect 376462 124378 393906 124614
rect 394142 124378 394226 124614
rect 394462 124378 411906 124614
rect 412142 124378 412226 124614
rect 412462 124378 429906 124614
rect 430142 124378 430226 124614
rect 430462 124378 447906 124614
rect 448142 124378 448226 124614
rect 448462 124378 465906 124614
rect 466142 124378 466226 124614
rect 466462 124378 483906 124614
rect 484142 124378 484226 124614
rect 484462 124378 501906 124614
rect 502142 124378 502226 124614
rect 502462 124378 519906 124614
rect 520142 124378 520226 124614
rect 520462 124378 537906 124614
rect 538142 124378 538226 124614
rect 538462 124378 547884 124614
rect 548120 124378 548204 124614
rect 548440 124378 548472 124614
rect -4476 124294 548472 124378
rect -4476 124058 -4444 124294
rect -4208 124058 -4124 124294
rect -3888 124058 15906 124294
rect 16142 124058 16226 124294
rect 16462 124058 33906 124294
rect 34142 124058 34226 124294
rect 34462 124058 51906 124294
rect 52142 124058 52226 124294
rect 52462 124058 69906 124294
rect 70142 124058 70226 124294
rect 70462 124058 87906 124294
rect 88142 124058 88226 124294
rect 88462 124058 105906 124294
rect 106142 124058 106226 124294
rect 106462 124058 123906 124294
rect 124142 124058 124226 124294
rect 124462 124058 141906 124294
rect 142142 124058 142226 124294
rect 142462 124058 159906 124294
rect 160142 124058 160226 124294
rect 160462 124058 177906 124294
rect 178142 124058 178226 124294
rect 178462 124058 195906 124294
rect 196142 124058 196226 124294
rect 196462 124058 213906 124294
rect 214142 124058 214226 124294
rect 214462 124058 231906 124294
rect 232142 124058 232226 124294
rect 232462 124058 249906 124294
rect 250142 124058 250226 124294
rect 250462 124058 267906 124294
rect 268142 124058 268226 124294
rect 268462 124058 285906 124294
rect 286142 124058 286226 124294
rect 286462 124058 303906 124294
rect 304142 124058 304226 124294
rect 304462 124058 321906 124294
rect 322142 124058 322226 124294
rect 322462 124058 339906 124294
rect 340142 124058 340226 124294
rect 340462 124058 357906 124294
rect 358142 124058 358226 124294
rect 358462 124058 375906 124294
rect 376142 124058 376226 124294
rect 376462 124058 393906 124294
rect 394142 124058 394226 124294
rect 394462 124058 411906 124294
rect 412142 124058 412226 124294
rect 412462 124058 429906 124294
rect 430142 124058 430226 124294
rect 430462 124058 447906 124294
rect 448142 124058 448226 124294
rect 448462 124058 465906 124294
rect 466142 124058 466226 124294
rect 466462 124058 483906 124294
rect 484142 124058 484226 124294
rect 484462 124058 501906 124294
rect 502142 124058 502226 124294
rect 502462 124058 519906 124294
rect 520142 124058 520226 124294
rect 520462 124058 537906 124294
rect 538142 124058 538226 124294
rect 538462 124058 547884 124294
rect 548120 124058 548204 124294
rect 548440 124058 548472 124294
rect -4476 124026 548472 124058
rect -4476 120894 548472 120926
rect -4476 120658 -3484 120894
rect -3248 120658 -3164 120894
rect -2928 120658 12186 120894
rect 12422 120658 12506 120894
rect 12742 120658 30186 120894
rect 30422 120658 30506 120894
rect 30742 120658 48186 120894
rect 48422 120658 48506 120894
rect 48742 120658 66186 120894
rect 66422 120658 66506 120894
rect 66742 120658 84186 120894
rect 84422 120658 84506 120894
rect 84742 120658 102186 120894
rect 102422 120658 102506 120894
rect 102742 120658 120186 120894
rect 120422 120658 120506 120894
rect 120742 120658 138186 120894
rect 138422 120658 138506 120894
rect 138742 120658 156186 120894
rect 156422 120658 156506 120894
rect 156742 120658 174186 120894
rect 174422 120658 174506 120894
rect 174742 120658 192186 120894
rect 192422 120658 192506 120894
rect 192742 120658 210186 120894
rect 210422 120658 210506 120894
rect 210742 120658 228186 120894
rect 228422 120658 228506 120894
rect 228742 120658 246186 120894
rect 246422 120658 246506 120894
rect 246742 120658 264186 120894
rect 264422 120658 264506 120894
rect 264742 120658 282186 120894
rect 282422 120658 282506 120894
rect 282742 120658 300186 120894
rect 300422 120658 300506 120894
rect 300742 120658 318186 120894
rect 318422 120658 318506 120894
rect 318742 120658 336186 120894
rect 336422 120658 336506 120894
rect 336742 120658 354186 120894
rect 354422 120658 354506 120894
rect 354742 120658 372186 120894
rect 372422 120658 372506 120894
rect 372742 120658 390186 120894
rect 390422 120658 390506 120894
rect 390742 120658 408186 120894
rect 408422 120658 408506 120894
rect 408742 120658 426186 120894
rect 426422 120658 426506 120894
rect 426742 120658 444186 120894
rect 444422 120658 444506 120894
rect 444742 120658 462186 120894
rect 462422 120658 462506 120894
rect 462742 120658 480186 120894
rect 480422 120658 480506 120894
rect 480742 120658 498186 120894
rect 498422 120658 498506 120894
rect 498742 120658 516186 120894
rect 516422 120658 516506 120894
rect 516742 120658 534186 120894
rect 534422 120658 534506 120894
rect 534742 120658 546924 120894
rect 547160 120658 547244 120894
rect 547480 120658 548472 120894
rect -4476 120574 548472 120658
rect -4476 120338 -3484 120574
rect -3248 120338 -3164 120574
rect -2928 120338 12186 120574
rect 12422 120338 12506 120574
rect 12742 120338 30186 120574
rect 30422 120338 30506 120574
rect 30742 120338 48186 120574
rect 48422 120338 48506 120574
rect 48742 120338 66186 120574
rect 66422 120338 66506 120574
rect 66742 120338 84186 120574
rect 84422 120338 84506 120574
rect 84742 120338 102186 120574
rect 102422 120338 102506 120574
rect 102742 120338 120186 120574
rect 120422 120338 120506 120574
rect 120742 120338 138186 120574
rect 138422 120338 138506 120574
rect 138742 120338 156186 120574
rect 156422 120338 156506 120574
rect 156742 120338 174186 120574
rect 174422 120338 174506 120574
rect 174742 120338 192186 120574
rect 192422 120338 192506 120574
rect 192742 120338 210186 120574
rect 210422 120338 210506 120574
rect 210742 120338 228186 120574
rect 228422 120338 228506 120574
rect 228742 120338 246186 120574
rect 246422 120338 246506 120574
rect 246742 120338 264186 120574
rect 264422 120338 264506 120574
rect 264742 120338 282186 120574
rect 282422 120338 282506 120574
rect 282742 120338 300186 120574
rect 300422 120338 300506 120574
rect 300742 120338 318186 120574
rect 318422 120338 318506 120574
rect 318742 120338 336186 120574
rect 336422 120338 336506 120574
rect 336742 120338 354186 120574
rect 354422 120338 354506 120574
rect 354742 120338 372186 120574
rect 372422 120338 372506 120574
rect 372742 120338 390186 120574
rect 390422 120338 390506 120574
rect 390742 120338 408186 120574
rect 408422 120338 408506 120574
rect 408742 120338 426186 120574
rect 426422 120338 426506 120574
rect 426742 120338 444186 120574
rect 444422 120338 444506 120574
rect 444742 120338 462186 120574
rect 462422 120338 462506 120574
rect 462742 120338 480186 120574
rect 480422 120338 480506 120574
rect 480742 120338 498186 120574
rect 498422 120338 498506 120574
rect 498742 120338 516186 120574
rect 516422 120338 516506 120574
rect 516742 120338 534186 120574
rect 534422 120338 534506 120574
rect 534742 120338 546924 120574
rect 547160 120338 547244 120574
rect 547480 120338 548472 120574
rect -4476 120306 548472 120338
rect -4476 117174 548472 117206
rect -4476 116938 -2524 117174
rect -2288 116938 -2204 117174
rect -1968 116938 8466 117174
rect 8702 116938 8786 117174
rect 9022 116938 26466 117174
rect 26702 116938 26786 117174
rect 27022 116938 44466 117174
rect 44702 116938 44786 117174
rect 45022 116938 62466 117174
rect 62702 116938 62786 117174
rect 63022 116938 80466 117174
rect 80702 116938 80786 117174
rect 81022 116938 98466 117174
rect 98702 116938 98786 117174
rect 99022 116938 116466 117174
rect 116702 116938 116786 117174
rect 117022 116938 134466 117174
rect 134702 116938 134786 117174
rect 135022 116938 152466 117174
rect 152702 116938 152786 117174
rect 153022 116938 170466 117174
rect 170702 116938 170786 117174
rect 171022 116938 188466 117174
rect 188702 116938 188786 117174
rect 189022 116938 206466 117174
rect 206702 116938 206786 117174
rect 207022 116938 224466 117174
rect 224702 116938 224786 117174
rect 225022 116938 242466 117174
rect 242702 116938 242786 117174
rect 243022 116938 260466 117174
rect 260702 116938 260786 117174
rect 261022 116938 278466 117174
rect 278702 116938 278786 117174
rect 279022 116938 296466 117174
rect 296702 116938 296786 117174
rect 297022 116938 314466 117174
rect 314702 116938 314786 117174
rect 315022 116938 332466 117174
rect 332702 116938 332786 117174
rect 333022 116938 350466 117174
rect 350702 116938 350786 117174
rect 351022 116938 368466 117174
rect 368702 116938 368786 117174
rect 369022 116938 386466 117174
rect 386702 116938 386786 117174
rect 387022 116938 404466 117174
rect 404702 116938 404786 117174
rect 405022 116938 422466 117174
rect 422702 116938 422786 117174
rect 423022 116938 440466 117174
rect 440702 116938 440786 117174
rect 441022 116938 458466 117174
rect 458702 116938 458786 117174
rect 459022 116938 476466 117174
rect 476702 116938 476786 117174
rect 477022 116938 494466 117174
rect 494702 116938 494786 117174
rect 495022 116938 512466 117174
rect 512702 116938 512786 117174
rect 513022 116938 530466 117174
rect 530702 116938 530786 117174
rect 531022 116938 545964 117174
rect 546200 116938 546284 117174
rect 546520 116938 548472 117174
rect -4476 116854 548472 116938
rect -4476 116618 -2524 116854
rect -2288 116618 -2204 116854
rect -1968 116618 8466 116854
rect 8702 116618 8786 116854
rect 9022 116618 26466 116854
rect 26702 116618 26786 116854
rect 27022 116618 44466 116854
rect 44702 116618 44786 116854
rect 45022 116618 62466 116854
rect 62702 116618 62786 116854
rect 63022 116618 80466 116854
rect 80702 116618 80786 116854
rect 81022 116618 98466 116854
rect 98702 116618 98786 116854
rect 99022 116618 116466 116854
rect 116702 116618 116786 116854
rect 117022 116618 134466 116854
rect 134702 116618 134786 116854
rect 135022 116618 152466 116854
rect 152702 116618 152786 116854
rect 153022 116618 170466 116854
rect 170702 116618 170786 116854
rect 171022 116618 188466 116854
rect 188702 116618 188786 116854
rect 189022 116618 206466 116854
rect 206702 116618 206786 116854
rect 207022 116618 224466 116854
rect 224702 116618 224786 116854
rect 225022 116618 242466 116854
rect 242702 116618 242786 116854
rect 243022 116618 260466 116854
rect 260702 116618 260786 116854
rect 261022 116618 278466 116854
rect 278702 116618 278786 116854
rect 279022 116618 296466 116854
rect 296702 116618 296786 116854
rect 297022 116618 314466 116854
rect 314702 116618 314786 116854
rect 315022 116618 332466 116854
rect 332702 116618 332786 116854
rect 333022 116618 350466 116854
rect 350702 116618 350786 116854
rect 351022 116618 368466 116854
rect 368702 116618 368786 116854
rect 369022 116618 386466 116854
rect 386702 116618 386786 116854
rect 387022 116618 404466 116854
rect 404702 116618 404786 116854
rect 405022 116618 422466 116854
rect 422702 116618 422786 116854
rect 423022 116618 440466 116854
rect 440702 116618 440786 116854
rect 441022 116618 458466 116854
rect 458702 116618 458786 116854
rect 459022 116618 476466 116854
rect 476702 116618 476786 116854
rect 477022 116618 494466 116854
rect 494702 116618 494786 116854
rect 495022 116618 512466 116854
rect 512702 116618 512786 116854
rect 513022 116618 530466 116854
rect 530702 116618 530786 116854
rect 531022 116618 545964 116854
rect 546200 116618 546284 116854
rect 546520 116618 548472 116854
rect -4476 116586 548472 116618
rect -4476 113454 548472 113486
rect -4476 113218 -1564 113454
rect -1328 113218 -1244 113454
rect -1008 113218 4746 113454
rect 4982 113218 5066 113454
rect 5302 113218 22746 113454
rect 22982 113218 23066 113454
rect 23302 113218 40746 113454
rect 40982 113218 41066 113454
rect 41302 113218 58746 113454
rect 58982 113218 59066 113454
rect 59302 113218 76746 113454
rect 76982 113218 77066 113454
rect 77302 113218 94746 113454
rect 94982 113218 95066 113454
rect 95302 113218 112746 113454
rect 112982 113218 113066 113454
rect 113302 113218 130746 113454
rect 130982 113218 131066 113454
rect 131302 113218 148746 113454
rect 148982 113218 149066 113454
rect 149302 113218 166746 113454
rect 166982 113218 167066 113454
rect 167302 113218 184746 113454
rect 184982 113218 185066 113454
rect 185302 113218 202746 113454
rect 202982 113218 203066 113454
rect 203302 113218 220746 113454
rect 220982 113218 221066 113454
rect 221302 113218 238746 113454
rect 238982 113218 239066 113454
rect 239302 113218 256746 113454
rect 256982 113218 257066 113454
rect 257302 113218 274746 113454
rect 274982 113218 275066 113454
rect 275302 113218 292746 113454
rect 292982 113218 293066 113454
rect 293302 113218 310746 113454
rect 310982 113218 311066 113454
rect 311302 113218 328746 113454
rect 328982 113218 329066 113454
rect 329302 113218 346746 113454
rect 346982 113218 347066 113454
rect 347302 113218 364746 113454
rect 364982 113218 365066 113454
rect 365302 113218 382746 113454
rect 382982 113218 383066 113454
rect 383302 113218 400746 113454
rect 400982 113218 401066 113454
rect 401302 113218 418746 113454
rect 418982 113218 419066 113454
rect 419302 113218 436746 113454
rect 436982 113218 437066 113454
rect 437302 113218 454746 113454
rect 454982 113218 455066 113454
rect 455302 113218 472746 113454
rect 472982 113218 473066 113454
rect 473302 113218 490746 113454
rect 490982 113218 491066 113454
rect 491302 113218 508746 113454
rect 508982 113218 509066 113454
rect 509302 113218 526746 113454
rect 526982 113218 527066 113454
rect 527302 113218 545004 113454
rect 545240 113218 545324 113454
rect 545560 113218 548472 113454
rect -4476 113134 548472 113218
rect -4476 112898 -1564 113134
rect -1328 112898 -1244 113134
rect -1008 112898 4746 113134
rect 4982 112898 5066 113134
rect 5302 112898 22746 113134
rect 22982 112898 23066 113134
rect 23302 112898 40746 113134
rect 40982 112898 41066 113134
rect 41302 112898 58746 113134
rect 58982 112898 59066 113134
rect 59302 112898 76746 113134
rect 76982 112898 77066 113134
rect 77302 112898 94746 113134
rect 94982 112898 95066 113134
rect 95302 112898 112746 113134
rect 112982 112898 113066 113134
rect 113302 112898 130746 113134
rect 130982 112898 131066 113134
rect 131302 112898 148746 113134
rect 148982 112898 149066 113134
rect 149302 112898 166746 113134
rect 166982 112898 167066 113134
rect 167302 112898 184746 113134
rect 184982 112898 185066 113134
rect 185302 112898 202746 113134
rect 202982 112898 203066 113134
rect 203302 112898 220746 113134
rect 220982 112898 221066 113134
rect 221302 112898 238746 113134
rect 238982 112898 239066 113134
rect 239302 112898 256746 113134
rect 256982 112898 257066 113134
rect 257302 112898 274746 113134
rect 274982 112898 275066 113134
rect 275302 112898 292746 113134
rect 292982 112898 293066 113134
rect 293302 112898 310746 113134
rect 310982 112898 311066 113134
rect 311302 112898 328746 113134
rect 328982 112898 329066 113134
rect 329302 112898 346746 113134
rect 346982 112898 347066 113134
rect 347302 112898 364746 113134
rect 364982 112898 365066 113134
rect 365302 112898 382746 113134
rect 382982 112898 383066 113134
rect 383302 112898 400746 113134
rect 400982 112898 401066 113134
rect 401302 112898 418746 113134
rect 418982 112898 419066 113134
rect 419302 112898 436746 113134
rect 436982 112898 437066 113134
rect 437302 112898 454746 113134
rect 454982 112898 455066 113134
rect 455302 112898 472746 113134
rect 472982 112898 473066 113134
rect 473302 112898 490746 113134
rect 490982 112898 491066 113134
rect 491302 112898 508746 113134
rect 508982 112898 509066 113134
rect 509302 112898 526746 113134
rect 526982 112898 527066 113134
rect 527302 112898 545004 113134
rect 545240 112898 545324 113134
rect 545560 112898 548472 113134
rect -4476 112866 548472 112898
rect -4476 106614 548472 106646
rect -4476 106378 -4444 106614
rect -4208 106378 -4124 106614
rect -3888 106378 15906 106614
rect 16142 106378 16226 106614
rect 16462 106378 33906 106614
rect 34142 106378 34226 106614
rect 34462 106378 51906 106614
rect 52142 106378 52226 106614
rect 52462 106378 69906 106614
rect 70142 106378 70226 106614
rect 70462 106378 87906 106614
rect 88142 106378 88226 106614
rect 88462 106378 105906 106614
rect 106142 106378 106226 106614
rect 106462 106378 123906 106614
rect 124142 106378 124226 106614
rect 124462 106378 141906 106614
rect 142142 106378 142226 106614
rect 142462 106378 159906 106614
rect 160142 106378 160226 106614
rect 160462 106378 177906 106614
rect 178142 106378 178226 106614
rect 178462 106378 195906 106614
rect 196142 106378 196226 106614
rect 196462 106378 213906 106614
rect 214142 106378 214226 106614
rect 214462 106378 231906 106614
rect 232142 106378 232226 106614
rect 232462 106378 249906 106614
rect 250142 106378 250226 106614
rect 250462 106378 267906 106614
rect 268142 106378 268226 106614
rect 268462 106378 285906 106614
rect 286142 106378 286226 106614
rect 286462 106378 303906 106614
rect 304142 106378 304226 106614
rect 304462 106378 321906 106614
rect 322142 106378 322226 106614
rect 322462 106378 339906 106614
rect 340142 106378 340226 106614
rect 340462 106378 357906 106614
rect 358142 106378 358226 106614
rect 358462 106378 375906 106614
rect 376142 106378 376226 106614
rect 376462 106378 393906 106614
rect 394142 106378 394226 106614
rect 394462 106378 411906 106614
rect 412142 106378 412226 106614
rect 412462 106378 429906 106614
rect 430142 106378 430226 106614
rect 430462 106378 447906 106614
rect 448142 106378 448226 106614
rect 448462 106378 465906 106614
rect 466142 106378 466226 106614
rect 466462 106378 483906 106614
rect 484142 106378 484226 106614
rect 484462 106378 501906 106614
rect 502142 106378 502226 106614
rect 502462 106378 519906 106614
rect 520142 106378 520226 106614
rect 520462 106378 537906 106614
rect 538142 106378 538226 106614
rect 538462 106378 547884 106614
rect 548120 106378 548204 106614
rect 548440 106378 548472 106614
rect -4476 106294 548472 106378
rect -4476 106058 -4444 106294
rect -4208 106058 -4124 106294
rect -3888 106058 15906 106294
rect 16142 106058 16226 106294
rect 16462 106058 33906 106294
rect 34142 106058 34226 106294
rect 34462 106058 51906 106294
rect 52142 106058 52226 106294
rect 52462 106058 69906 106294
rect 70142 106058 70226 106294
rect 70462 106058 87906 106294
rect 88142 106058 88226 106294
rect 88462 106058 105906 106294
rect 106142 106058 106226 106294
rect 106462 106058 123906 106294
rect 124142 106058 124226 106294
rect 124462 106058 141906 106294
rect 142142 106058 142226 106294
rect 142462 106058 159906 106294
rect 160142 106058 160226 106294
rect 160462 106058 177906 106294
rect 178142 106058 178226 106294
rect 178462 106058 195906 106294
rect 196142 106058 196226 106294
rect 196462 106058 213906 106294
rect 214142 106058 214226 106294
rect 214462 106058 231906 106294
rect 232142 106058 232226 106294
rect 232462 106058 249906 106294
rect 250142 106058 250226 106294
rect 250462 106058 267906 106294
rect 268142 106058 268226 106294
rect 268462 106058 285906 106294
rect 286142 106058 286226 106294
rect 286462 106058 303906 106294
rect 304142 106058 304226 106294
rect 304462 106058 321906 106294
rect 322142 106058 322226 106294
rect 322462 106058 339906 106294
rect 340142 106058 340226 106294
rect 340462 106058 357906 106294
rect 358142 106058 358226 106294
rect 358462 106058 375906 106294
rect 376142 106058 376226 106294
rect 376462 106058 393906 106294
rect 394142 106058 394226 106294
rect 394462 106058 411906 106294
rect 412142 106058 412226 106294
rect 412462 106058 429906 106294
rect 430142 106058 430226 106294
rect 430462 106058 447906 106294
rect 448142 106058 448226 106294
rect 448462 106058 465906 106294
rect 466142 106058 466226 106294
rect 466462 106058 483906 106294
rect 484142 106058 484226 106294
rect 484462 106058 501906 106294
rect 502142 106058 502226 106294
rect 502462 106058 519906 106294
rect 520142 106058 520226 106294
rect 520462 106058 537906 106294
rect 538142 106058 538226 106294
rect 538462 106058 547884 106294
rect 548120 106058 548204 106294
rect 548440 106058 548472 106294
rect -4476 106026 548472 106058
rect -4476 102894 548472 102926
rect -4476 102658 -3484 102894
rect -3248 102658 -3164 102894
rect -2928 102658 12186 102894
rect 12422 102658 12506 102894
rect 12742 102658 30186 102894
rect 30422 102658 30506 102894
rect 30742 102658 48186 102894
rect 48422 102658 48506 102894
rect 48742 102658 66186 102894
rect 66422 102658 66506 102894
rect 66742 102658 84186 102894
rect 84422 102658 84506 102894
rect 84742 102658 102186 102894
rect 102422 102658 102506 102894
rect 102742 102658 120186 102894
rect 120422 102658 120506 102894
rect 120742 102658 138186 102894
rect 138422 102658 138506 102894
rect 138742 102658 156186 102894
rect 156422 102658 156506 102894
rect 156742 102658 174186 102894
rect 174422 102658 174506 102894
rect 174742 102658 192186 102894
rect 192422 102658 192506 102894
rect 192742 102658 210186 102894
rect 210422 102658 210506 102894
rect 210742 102658 228186 102894
rect 228422 102658 228506 102894
rect 228742 102658 246186 102894
rect 246422 102658 246506 102894
rect 246742 102658 264186 102894
rect 264422 102658 264506 102894
rect 264742 102658 282186 102894
rect 282422 102658 282506 102894
rect 282742 102658 300186 102894
rect 300422 102658 300506 102894
rect 300742 102658 318186 102894
rect 318422 102658 318506 102894
rect 318742 102658 336186 102894
rect 336422 102658 336506 102894
rect 336742 102658 354186 102894
rect 354422 102658 354506 102894
rect 354742 102658 372186 102894
rect 372422 102658 372506 102894
rect 372742 102658 390186 102894
rect 390422 102658 390506 102894
rect 390742 102658 408186 102894
rect 408422 102658 408506 102894
rect 408742 102658 426186 102894
rect 426422 102658 426506 102894
rect 426742 102658 444186 102894
rect 444422 102658 444506 102894
rect 444742 102658 462186 102894
rect 462422 102658 462506 102894
rect 462742 102658 480186 102894
rect 480422 102658 480506 102894
rect 480742 102658 498186 102894
rect 498422 102658 498506 102894
rect 498742 102658 516186 102894
rect 516422 102658 516506 102894
rect 516742 102658 534186 102894
rect 534422 102658 534506 102894
rect 534742 102658 546924 102894
rect 547160 102658 547244 102894
rect 547480 102658 548472 102894
rect -4476 102574 548472 102658
rect -4476 102338 -3484 102574
rect -3248 102338 -3164 102574
rect -2928 102338 12186 102574
rect 12422 102338 12506 102574
rect 12742 102338 30186 102574
rect 30422 102338 30506 102574
rect 30742 102338 48186 102574
rect 48422 102338 48506 102574
rect 48742 102338 66186 102574
rect 66422 102338 66506 102574
rect 66742 102338 84186 102574
rect 84422 102338 84506 102574
rect 84742 102338 102186 102574
rect 102422 102338 102506 102574
rect 102742 102338 120186 102574
rect 120422 102338 120506 102574
rect 120742 102338 138186 102574
rect 138422 102338 138506 102574
rect 138742 102338 156186 102574
rect 156422 102338 156506 102574
rect 156742 102338 174186 102574
rect 174422 102338 174506 102574
rect 174742 102338 192186 102574
rect 192422 102338 192506 102574
rect 192742 102338 210186 102574
rect 210422 102338 210506 102574
rect 210742 102338 228186 102574
rect 228422 102338 228506 102574
rect 228742 102338 246186 102574
rect 246422 102338 246506 102574
rect 246742 102338 264186 102574
rect 264422 102338 264506 102574
rect 264742 102338 282186 102574
rect 282422 102338 282506 102574
rect 282742 102338 300186 102574
rect 300422 102338 300506 102574
rect 300742 102338 318186 102574
rect 318422 102338 318506 102574
rect 318742 102338 336186 102574
rect 336422 102338 336506 102574
rect 336742 102338 354186 102574
rect 354422 102338 354506 102574
rect 354742 102338 372186 102574
rect 372422 102338 372506 102574
rect 372742 102338 390186 102574
rect 390422 102338 390506 102574
rect 390742 102338 408186 102574
rect 408422 102338 408506 102574
rect 408742 102338 426186 102574
rect 426422 102338 426506 102574
rect 426742 102338 444186 102574
rect 444422 102338 444506 102574
rect 444742 102338 462186 102574
rect 462422 102338 462506 102574
rect 462742 102338 480186 102574
rect 480422 102338 480506 102574
rect 480742 102338 498186 102574
rect 498422 102338 498506 102574
rect 498742 102338 516186 102574
rect 516422 102338 516506 102574
rect 516742 102338 534186 102574
rect 534422 102338 534506 102574
rect 534742 102338 546924 102574
rect 547160 102338 547244 102574
rect 547480 102338 548472 102574
rect -4476 102306 548472 102338
rect -4476 99174 548472 99206
rect -4476 98938 -2524 99174
rect -2288 98938 -2204 99174
rect -1968 98938 8466 99174
rect 8702 98938 8786 99174
rect 9022 98938 26466 99174
rect 26702 98938 26786 99174
rect 27022 98938 44466 99174
rect 44702 98938 44786 99174
rect 45022 98938 62466 99174
rect 62702 98938 62786 99174
rect 63022 98938 80466 99174
rect 80702 98938 80786 99174
rect 81022 98938 98466 99174
rect 98702 98938 98786 99174
rect 99022 98938 116466 99174
rect 116702 98938 116786 99174
rect 117022 98938 134466 99174
rect 134702 98938 134786 99174
rect 135022 98938 152466 99174
rect 152702 98938 152786 99174
rect 153022 98938 170466 99174
rect 170702 98938 170786 99174
rect 171022 98938 188466 99174
rect 188702 98938 188786 99174
rect 189022 98938 206466 99174
rect 206702 98938 206786 99174
rect 207022 98938 224466 99174
rect 224702 98938 224786 99174
rect 225022 98938 242466 99174
rect 242702 98938 242786 99174
rect 243022 98938 260466 99174
rect 260702 98938 260786 99174
rect 261022 98938 278466 99174
rect 278702 98938 278786 99174
rect 279022 98938 296466 99174
rect 296702 98938 296786 99174
rect 297022 98938 314466 99174
rect 314702 98938 314786 99174
rect 315022 98938 332466 99174
rect 332702 98938 332786 99174
rect 333022 98938 350466 99174
rect 350702 98938 350786 99174
rect 351022 98938 368466 99174
rect 368702 98938 368786 99174
rect 369022 98938 386466 99174
rect 386702 98938 386786 99174
rect 387022 98938 404466 99174
rect 404702 98938 404786 99174
rect 405022 98938 422466 99174
rect 422702 98938 422786 99174
rect 423022 98938 440466 99174
rect 440702 98938 440786 99174
rect 441022 98938 458466 99174
rect 458702 98938 458786 99174
rect 459022 98938 476466 99174
rect 476702 98938 476786 99174
rect 477022 98938 494466 99174
rect 494702 98938 494786 99174
rect 495022 98938 512466 99174
rect 512702 98938 512786 99174
rect 513022 98938 530466 99174
rect 530702 98938 530786 99174
rect 531022 98938 545964 99174
rect 546200 98938 546284 99174
rect 546520 98938 548472 99174
rect -4476 98854 548472 98938
rect -4476 98618 -2524 98854
rect -2288 98618 -2204 98854
rect -1968 98618 8466 98854
rect 8702 98618 8786 98854
rect 9022 98618 26466 98854
rect 26702 98618 26786 98854
rect 27022 98618 44466 98854
rect 44702 98618 44786 98854
rect 45022 98618 62466 98854
rect 62702 98618 62786 98854
rect 63022 98618 80466 98854
rect 80702 98618 80786 98854
rect 81022 98618 98466 98854
rect 98702 98618 98786 98854
rect 99022 98618 116466 98854
rect 116702 98618 116786 98854
rect 117022 98618 134466 98854
rect 134702 98618 134786 98854
rect 135022 98618 152466 98854
rect 152702 98618 152786 98854
rect 153022 98618 170466 98854
rect 170702 98618 170786 98854
rect 171022 98618 188466 98854
rect 188702 98618 188786 98854
rect 189022 98618 206466 98854
rect 206702 98618 206786 98854
rect 207022 98618 224466 98854
rect 224702 98618 224786 98854
rect 225022 98618 242466 98854
rect 242702 98618 242786 98854
rect 243022 98618 260466 98854
rect 260702 98618 260786 98854
rect 261022 98618 278466 98854
rect 278702 98618 278786 98854
rect 279022 98618 296466 98854
rect 296702 98618 296786 98854
rect 297022 98618 314466 98854
rect 314702 98618 314786 98854
rect 315022 98618 332466 98854
rect 332702 98618 332786 98854
rect 333022 98618 350466 98854
rect 350702 98618 350786 98854
rect 351022 98618 368466 98854
rect 368702 98618 368786 98854
rect 369022 98618 386466 98854
rect 386702 98618 386786 98854
rect 387022 98618 404466 98854
rect 404702 98618 404786 98854
rect 405022 98618 422466 98854
rect 422702 98618 422786 98854
rect 423022 98618 440466 98854
rect 440702 98618 440786 98854
rect 441022 98618 458466 98854
rect 458702 98618 458786 98854
rect 459022 98618 476466 98854
rect 476702 98618 476786 98854
rect 477022 98618 494466 98854
rect 494702 98618 494786 98854
rect 495022 98618 512466 98854
rect 512702 98618 512786 98854
rect 513022 98618 530466 98854
rect 530702 98618 530786 98854
rect 531022 98618 545964 98854
rect 546200 98618 546284 98854
rect 546520 98618 548472 98854
rect -4476 98586 548472 98618
rect -4476 95454 548472 95486
rect -4476 95218 -1564 95454
rect -1328 95218 -1244 95454
rect -1008 95218 4746 95454
rect 4982 95218 5066 95454
rect 5302 95218 22746 95454
rect 22982 95218 23066 95454
rect 23302 95218 40746 95454
rect 40982 95218 41066 95454
rect 41302 95218 58746 95454
rect 58982 95218 59066 95454
rect 59302 95218 76746 95454
rect 76982 95218 77066 95454
rect 77302 95218 94746 95454
rect 94982 95218 95066 95454
rect 95302 95218 112746 95454
rect 112982 95218 113066 95454
rect 113302 95218 130746 95454
rect 130982 95218 131066 95454
rect 131302 95218 148746 95454
rect 148982 95218 149066 95454
rect 149302 95218 166746 95454
rect 166982 95218 167066 95454
rect 167302 95218 184746 95454
rect 184982 95218 185066 95454
rect 185302 95218 202746 95454
rect 202982 95218 203066 95454
rect 203302 95218 220746 95454
rect 220982 95218 221066 95454
rect 221302 95218 238746 95454
rect 238982 95218 239066 95454
rect 239302 95218 256746 95454
rect 256982 95218 257066 95454
rect 257302 95218 274746 95454
rect 274982 95218 275066 95454
rect 275302 95218 292746 95454
rect 292982 95218 293066 95454
rect 293302 95218 310746 95454
rect 310982 95218 311066 95454
rect 311302 95218 328746 95454
rect 328982 95218 329066 95454
rect 329302 95218 346746 95454
rect 346982 95218 347066 95454
rect 347302 95218 364746 95454
rect 364982 95218 365066 95454
rect 365302 95218 382746 95454
rect 382982 95218 383066 95454
rect 383302 95218 400746 95454
rect 400982 95218 401066 95454
rect 401302 95218 418746 95454
rect 418982 95218 419066 95454
rect 419302 95218 436746 95454
rect 436982 95218 437066 95454
rect 437302 95218 454746 95454
rect 454982 95218 455066 95454
rect 455302 95218 472746 95454
rect 472982 95218 473066 95454
rect 473302 95218 490746 95454
rect 490982 95218 491066 95454
rect 491302 95218 508746 95454
rect 508982 95218 509066 95454
rect 509302 95218 526746 95454
rect 526982 95218 527066 95454
rect 527302 95218 545004 95454
rect 545240 95218 545324 95454
rect 545560 95218 548472 95454
rect -4476 95134 548472 95218
rect -4476 94898 -1564 95134
rect -1328 94898 -1244 95134
rect -1008 94898 4746 95134
rect 4982 94898 5066 95134
rect 5302 94898 22746 95134
rect 22982 94898 23066 95134
rect 23302 94898 40746 95134
rect 40982 94898 41066 95134
rect 41302 94898 58746 95134
rect 58982 94898 59066 95134
rect 59302 94898 76746 95134
rect 76982 94898 77066 95134
rect 77302 94898 94746 95134
rect 94982 94898 95066 95134
rect 95302 94898 112746 95134
rect 112982 94898 113066 95134
rect 113302 94898 130746 95134
rect 130982 94898 131066 95134
rect 131302 94898 148746 95134
rect 148982 94898 149066 95134
rect 149302 94898 166746 95134
rect 166982 94898 167066 95134
rect 167302 94898 184746 95134
rect 184982 94898 185066 95134
rect 185302 94898 202746 95134
rect 202982 94898 203066 95134
rect 203302 94898 220746 95134
rect 220982 94898 221066 95134
rect 221302 94898 238746 95134
rect 238982 94898 239066 95134
rect 239302 94898 256746 95134
rect 256982 94898 257066 95134
rect 257302 94898 274746 95134
rect 274982 94898 275066 95134
rect 275302 94898 292746 95134
rect 292982 94898 293066 95134
rect 293302 94898 310746 95134
rect 310982 94898 311066 95134
rect 311302 94898 328746 95134
rect 328982 94898 329066 95134
rect 329302 94898 346746 95134
rect 346982 94898 347066 95134
rect 347302 94898 364746 95134
rect 364982 94898 365066 95134
rect 365302 94898 382746 95134
rect 382982 94898 383066 95134
rect 383302 94898 400746 95134
rect 400982 94898 401066 95134
rect 401302 94898 418746 95134
rect 418982 94898 419066 95134
rect 419302 94898 436746 95134
rect 436982 94898 437066 95134
rect 437302 94898 454746 95134
rect 454982 94898 455066 95134
rect 455302 94898 472746 95134
rect 472982 94898 473066 95134
rect 473302 94898 490746 95134
rect 490982 94898 491066 95134
rect 491302 94898 508746 95134
rect 508982 94898 509066 95134
rect 509302 94898 526746 95134
rect 526982 94898 527066 95134
rect 527302 94898 545004 95134
rect 545240 94898 545324 95134
rect 545560 94898 548472 95134
rect -4476 94866 548472 94898
rect -4476 88614 548472 88646
rect -4476 88378 -4444 88614
rect -4208 88378 -4124 88614
rect -3888 88378 15906 88614
rect 16142 88378 16226 88614
rect 16462 88378 33906 88614
rect 34142 88378 34226 88614
rect 34462 88378 51906 88614
rect 52142 88378 52226 88614
rect 52462 88378 69906 88614
rect 70142 88378 70226 88614
rect 70462 88378 87906 88614
rect 88142 88378 88226 88614
rect 88462 88378 105906 88614
rect 106142 88378 106226 88614
rect 106462 88378 123906 88614
rect 124142 88378 124226 88614
rect 124462 88378 141906 88614
rect 142142 88378 142226 88614
rect 142462 88378 159906 88614
rect 160142 88378 160226 88614
rect 160462 88378 177906 88614
rect 178142 88378 178226 88614
rect 178462 88378 195906 88614
rect 196142 88378 196226 88614
rect 196462 88378 213906 88614
rect 214142 88378 214226 88614
rect 214462 88378 231906 88614
rect 232142 88378 232226 88614
rect 232462 88378 249906 88614
rect 250142 88378 250226 88614
rect 250462 88378 267906 88614
rect 268142 88378 268226 88614
rect 268462 88378 285906 88614
rect 286142 88378 286226 88614
rect 286462 88378 303906 88614
rect 304142 88378 304226 88614
rect 304462 88378 321906 88614
rect 322142 88378 322226 88614
rect 322462 88378 339906 88614
rect 340142 88378 340226 88614
rect 340462 88378 357906 88614
rect 358142 88378 358226 88614
rect 358462 88378 375906 88614
rect 376142 88378 376226 88614
rect 376462 88378 393906 88614
rect 394142 88378 394226 88614
rect 394462 88378 411906 88614
rect 412142 88378 412226 88614
rect 412462 88378 429906 88614
rect 430142 88378 430226 88614
rect 430462 88378 447906 88614
rect 448142 88378 448226 88614
rect 448462 88378 465906 88614
rect 466142 88378 466226 88614
rect 466462 88378 483906 88614
rect 484142 88378 484226 88614
rect 484462 88378 501906 88614
rect 502142 88378 502226 88614
rect 502462 88378 519906 88614
rect 520142 88378 520226 88614
rect 520462 88378 537906 88614
rect 538142 88378 538226 88614
rect 538462 88378 547884 88614
rect 548120 88378 548204 88614
rect 548440 88378 548472 88614
rect -4476 88294 548472 88378
rect -4476 88058 -4444 88294
rect -4208 88058 -4124 88294
rect -3888 88058 15906 88294
rect 16142 88058 16226 88294
rect 16462 88058 33906 88294
rect 34142 88058 34226 88294
rect 34462 88058 51906 88294
rect 52142 88058 52226 88294
rect 52462 88058 69906 88294
rect 70142 88058 70226 88294
rect 70462 88058 87906 88294
rect 88142 88058 88226 88294
rect 88462 88058 105906 88294
rect 106142 88058 106226 88294
rect 106462 88058 123906 88294
rect 124142 88058 124226 88294
rect 124462 88058 141906 88294
rect 142142 88058 142226 88294
rect 142462 88058 159906 88294
rect 160142 88058 160226 88294
rect 160462 88058 177906 88294
rect 178142 88058 178226 88294
rect 178462 88058 195906 88294
rect 196142 88058 196226 88294
rect 196462 88058 213906 88294
rect 214142 88058 214226 88294
rect 214462 88058 231906 88294
rect 232142 88058 232226 88294
rect 232462 88058 249906 88294
rect 250142 88058 250226 88294
rect 250462 88058 267906 88294
rect 268142 88058 268226 88294
rect 268462 88058 285906 88294
rect 286142 88058 286226 88294
rect 286462 88058 303906 88294
rect 304142 88058 304226 88294
rect 304462 88058 321906 88294
rect 322142 88058 322226 88294
rect 322462 88058 339906 88294
rect 340142 88058 340226 88294
rect 340462 88058 357906 88294
rect 358142 88058 358226 88294
rect 358462 88058 375906 88294
rect 376142 88058 376226 88294
rect 376462 88058 393906 88294
rect 394142 88058 394226 88294
rect 394462 88058 411906 88294
rect 412142 88058 412226 88294
rect 412462 88058 429906 88294
rect 430142 88058 430226 88294
rect 430462 88058 447906 88294
rect 448142 88058 448226 88294
rect 448462 88058 465906 88294
rect 466142 88058 466226 88294
rect 466462 88058 483906 88294
rect 484142 88058 484226 88294
rect 484462 88058 501906 88294
rect 502142 88058 502226 88294
rect 502462 88058 519906 88294
rect 520142 88058 520226 88294
rect 520462 88058 537906 88294
rect 538142 88058 538226 88294
rect 538462 88058 547884 88294
rect 548120 88058 548204 88294
rect 548440 88058 548472 88294
rect -4476 88026 548472 88058
rect -4476 84894 548472 84926
rect -4476 84658 -3484 84894
rect -3248 84658 -3164 84894
rect -2928 84658 12186 84894
rect 12422 84658 12506 84894
rect 12742 84658 30186 84894
rect 30422 84658 30506 84894
rect 30742 84658 48186 84894
rect 48422 84658 48506 84894
rect 48742 84658 66186 84894
rect 66422 84658 66506 84894
rect 66742 84658 84186 84894
rect 84422 84658 84506 84894
rect 84742 84658 102186 84894
rect 102422 84658 102506 84894
rect 102742 84658 120186 84894
rect 120422 84658 120506 84894
rect 120742 84658 138186 84894
rect 138422 84658 138506 84894
rect 138742 84658 156186 84894
rect 156422 84658 156506 84894
rect 156742 84658 174186 84894
rect 174422 84658 174506 84894
rect 174742 84658 192186 84894
rect 192422 84658 192506 84894
rect 192742 84658 210186 84894
rect 210422 84658 210506 84894
rect 210742 84658 228186 84894
rect 228422 84658 228506 84894
rect 228742 84658 246186 84894
rect 246422 84658 246506 84894
rect 246742 84658 264186 84894
rect 264422 84658 264506 84894
rect 264742 84658 282186 84894
rect 282422 84658 282506 84894
rect 282742 84658 300186 84894
rect 300422 84658 300506 84894
rect 300742 84658 318186 84894
rect 318422 84658 318506 84894
rect 318742 84658 336186 84894
rect 336422 84658 336506 84894
rect 336742 84658 354186 84894
rect 354422 84658 354506 84894
rect 354742 84658 372186 84894
rect 372422 84658 372506 84894
rect 372742 84658 390186 84894
rect 390422 84658 390506 84894
rect 390742 84658 408186 84894
rect 408422 84658 408506 84894
rect 408742 84658 426186 84894
rect 426422 84658 426506 84894
rect 426742 84658 444186 84894
rect 444422 84658 444506 84894
rect 444742 84658 462186 84894
rect 462422 84658 462506 84894
rect 462742 84658 480186 84894
rect 480422 84658 480506 84894
rect 480742 84658 498186 84894
rect 498422 84658 498506 84894
rect 498742 84658 516186 84894
rect 516422 84658 516506 84894
rect 516742 84658 534186 84894
rect 534422 84658 534506 84894
rect 534742 84658 546924 84894
rect 547160 84658 547244 84894
rect 547480 84658 548472 84894
rect -4476 84574 548472 84658
rect -4476 84338 -3484 84574
rect -3248 84338 -3164 84574
rect -2928 84338 12186 84574
rect 12422 84338 12506 84574
rect 12742 84338 30186 84574
rect 30422 84338 30506 84574
rect 30742 84338 48186 84574
rect 48422 84338 48506 84574
rect 48742 84338 66186 84574
rect 66422 84338 66506 84574
rect 66742 84338 84186 84574
rect 84422 84338 84506 84574
rect 84742 84338 102186 84574
rect 102422 84338 102506 84574
rect 102742 84338 120186 84574
rect 120422 84338 120506 84574
rect 120742 84338 138186 84574
rect 138422 84338 138506 84574
rect 138742 84338 156186 84574
rect 156422 84338 156506 84574
rect 156742 84338 174186 84574
rect 174422 84338 174506 84574
rect 174742 84338 192186 84574
rect 192422 84338 192506 84574
rect 192742 84338 210186 84574
rect 210422 84338 210506 84574
rect 210742 84338 228186 84574
rect 228422 84338 228506 84574
rect 228742 84338 246186 84574
rect 246422 84338 246506 84574
rect 246742 84338 264186 84574
rect 264422 84338 264506 84574
rect 264742 84338 282186 84574
rect 282422 84338 282506 84574
rect 282742 84338 300186 84574
rect 300422 84338 300506 84574
rect 300742 84338 318186 84574
rect 318422 84338 318506 84574
rect 318742 84338 336186 84574
rect 336422 84338 336506 84574
rect 336742 84338 354186 84574
rect 354422 84338 354506 84574
rect 354742 84338 372186 84574
rect 372422 84338 372506 84574
rect 372742 84338 390186 84574
rect 390422 84338 390506 84574
rect 390742 84338 408186 84574
rect 408422 84338 408506 84574
rect 408742 84338 426186 84574
rect 426422 84338 426506 84574
rect 426742 84338 444186 84574
rect 444422 84338 444506 84574
rect 444742 84338 462186 84574
rect 462422 84338 462506 84574
rect 462742 84338 480186 84574
rect 480422 84338 480506 84574
rect 480742 84338 498186 84574
rect 498422 84338 498506 84574
rect 498742 84338 516186 84574
rect 516422 84338 516506 84574
rect 516742 84338 534186 84574
rect 534422 84338 534506 84574
rect 534742 84338 546924 84574
rect 547160 84338 547244 84574
rect 547480 84338 548472 84574
rect -4476 84306 548472 84338
rect -4476 81174 548472 81206
rect -4476 80938 -2524 81174
rect -2288 80938 -2204 81174
rect -1968 80938 8466 81174
rect 8702 80938 8786 81174
rect 9022 80938 26466 81174
rect 26702 80938 26786 81174
rect 27022 80938 44466 81174
rect 44702 80938 44786 81174
rect 45022 80938 62466 81174
rect 62702 80938 62786 81174
rect 63022 80938 80466 81174
rect 80702 80938 80786 81174
rect 81022 80938 98466 81174
rect 98702 80938 98786 81174
rect 99022 80938 116466 81174
rect 116702 80938 116786 81174
rect 117022 80938 134466 81174
rect 134702 80938 134786 81174
rect 135022 80938 152466 81174
rect 152702 80938 152786 81174
rect 153022 80938 170466 81174
rect 170702 80938 170786 81174
rect 171022 80938 188466 81174
rect 188702 80938 188786 81174
rect 189022 80938 206466 81174
rect 206702 80938 206786 81174
rect 207022 80938 224466 81174
rect 224702 80938 224786 81174
rect 225022 80938 242466 81174
rect 242702 80938 242786 81174
rect 243022 80938 260466 81174
rect 260702 80938 260786 81174
rect 261022 80938 278466 81174
rect 278702 80938 278786 81174
rect 279022 80938 296466 81174
rect 296702 80938 296786 81174
rect 297022 80938 314466 81174
rect 314702 80938 314786 81174
rect 315022 80938 332466 81174
rect 332702 80938 332786 81174
rect 333022 80938 350466 81174
rect 350702 80938 350786 81174
rect 351022 80938 368466 81174
rect 368702 80938 368786 81174
rect 369022 80938 386466 81174
rect 386702 80938 386786 81174
rect 387022 80938 404466 81174
rect 404702 80938 404786 81174
rect 405022 80938 422466 81174
rect 422702 80938 422786 81174
rect 423022 80938 440466 81174
rect 440702 80938 440786 81174
rect 441022 80938 458466 81174
rect 458702 80938 458786 81174
rect 459022 80938 476466 81174
rect 476702 80938 476786 81174
rect 477022 80938 494466 81174
rect 494702 80938 494786 81174
rect 495022 80938 512466 81174
rect 512702 80938 512786 81174
rect 513022 80938 530466 81174
rect 530702 80938 530786 81174
rect 531022 80938 545964 81174
rect 546200 80938 546284 81174
rect 546520 80938 548472 81174
rect -4476 80854 548472 80938
rect -4476 80618 -2524 80854
rect -2288 80618 -2204 80854
rect -1968 80618 8466 80854
rect 8702 80618 8786 80854
rect 9022 80618 26466 80854
rect 26702 80618 26786 80854
rect 27022 80618 44466 80854
rect 44702 80618 44786 80854
rect 45022 80618 62466 80854
rect 62702 80618 62786 80854
rect 63022 80618 80466 80854
rect 80702 80618 80786 80854
rect 81022 80618 98466 80854
rect 98702 80618 98786 80854
rect 99022 80618 116466 80854
rect 116702 80618 116786 80854
rect 117022 80618 134466 80854
rect 134702 80618 134786 80854
rect 135022 80618 152466 80854
rect 152702 80618 152786 80854
rect 153022 80618 170466 80854
rect 170702 80618 170786 80854
rect 171022 80618 188466 80854
rect 188702 80618 188786 80854
rect 189022 80618 206466 80854
rect 206702 80618 206786 80854
rect 207022 80618 224466 80854
rect 224702 80618 224786 80854
rect 225022 80618 242466 80854
rect 242702 80618 242786 80854
rect 243022 80618 260466 80854
rect 260702 80618 260786 80854
rect 261022 80618 278466 80854
rect 278702 80618 278786 80854
rect 279022 80618 296466 80854
rect 296702 80618 296786 80854
rect 297022 80618 314466 80854
rect 314702 80618 314786 80854
rect 315022 80618 332466 80854
rect 332702 80618 332786 80854
rect 333022 80618 350466 80854
rect 350702 80618 350786 80854
rect 351022 80618 368466 80854
rect 368702 80618 368786 80854
rect 369022 80618 386466 80854
rect 386702 80618 386786 80854
rect 387022 80618 404466 80854
rect 404702 80618 404786 80854
rect 405022 80618 422466 80854
rect 422702 80618 422786 80854
rect 423022 80618 440466 80854
rect 440702 80618 440786 80854
rect 441022 80618 458466 80854
rect 458702 80618 458786 80854
rect 459022 80618 476466 80854
rect 476702 80618 476786 80854
rect 477022 80618 494466 80854
rect 494702 80618 494786 80854
rect 495022 80618 512466 80854
rect 512702 80618 512786 80854
rect 513022 80618 530466 80854
rect 530702 80618 530786 80854
rect 531022 80618 545964 80854
rect 546200 80618 546284 80854
rect 546520 80618 548472 80854
rect -4476 80586 548472 80618
rect -4476 77454 548472 77486
rect -4476 77218 -1564 77454
rect -1328 77218 -1244 77454
rect -1008 77218 4746 77454
rect 4982 77218 5066 77454
rect 5302 77218 22746 77454
rect 22982 77218 23066 77454
rect 23302 77218 40746 77454
rect 40982 77218 41066 77454
rect 41302 77218 58746 77454
rect 58982 77218 59066 77454
rect 59302 77218 76746 77454
rect 76982 77218 77066 77454
rect 77302 77218 94746 77454
rect 94982 77218 95066 77454
rect 95302 77218 112746 77454
rect 112982 77218 113066 77454
rect 113302 77218 130746 77454
rect 130982 77218 131066 77454
rect 131302 77218 148746 77454
rect 148982 77218 149066 77454
rect 149302 77218 166746 77454
rect 166982 77218 167066 77454
rect 167302 77218 184746 77454
rect 184982 77218 185066 77454
rect 185302 77218 202746 77454
rect 202982 77218 203066 77454
rect 203302 77218 220746 77454
rect 220982 77218 221066 77454
rect 221302 77218 238746 77454
rect 238982 77218 239066 77454
rect 239302 77218 256746 77454
rect 256982 77218 257066 77454
rect 257302 77218 274746 77454
rect 274982 77218 275066 77454
rect 275302 77218 292746 77454
rect 292982 77218 293066 77454
rect 293302 77218 310746 77454
rect 310982 77218 311066 77454
rect 311302 77218 328746 77454
rect 328982 77218 329066 77454
rect 329302 77218 346746 77454
rect 346982 77218 347066 77454
rect 347302 77218 364746 77454
rect 364982 77218 365066 77454
rect 365302 77218 382746 77454
rect 382982 77218 383066 77454
rect 383302 77218 400746 77454
rect 400982 77218 401066 77454
rect 401302 77218 418746 77454
rect 418982 77218 419066 77454
rect 419302 77218 436746 77454
rect 436982 77218 437066 77454
rect 437302 77218 454746 77454
rect 454982 77218 455066 77454
rect 455302 77218 472746 77454
rect 472982 77218 473066 77454
rect 473302 77218 490746 77454
rect 490982 77218 491066 77454
rect 491302 77218 508746 77454
rect 508982 77218 509066 77454
rect 509302 77218 526746 77454
rect 526982 77218 527066 77454
rect 527302 77218 545004 77454
rect 545240 77218 545324 77454
rect 545560 77218 548472 77454
rect -4476 77134 548472 77218
rect -4476 76898 -1564 77134
rect -1328 76898 -1244 77134
rect -1008 76898 4746 77134
rect 4982 76898 5066 77134
rect 5302 76898 22746 77134
rect 22982 76898 23066 77134
rect 23302 76898 40746 77134
rect 40982 76898 41066 77134
rect 41302 76898 58746 77134
rect 58982 76898 59066 77134
rect 59302 76898 76746 77134
rect 76982 76898 77066 77134
rect 77302 76898 94746 77134
rect 94982 76898 95066 77134
rect 95302 76898 112746 77134
rect 112982 76898 113066 77134
rect 113302 76898 130746 77134
rect 130982 76898 131066 77134
rect 131302 76898 148746 77134
rect 148982 76898 149066 77134
rect 149302 76898 166746 77134
rect 166982 76898 167066 77134
rect 167302 76898 184746 77134
rect 184982 76898 185066 77134
rect 185302 76898 202746 77134
rect 202982 76898 203066 77134
rect 203302 76898 220746 77134
rect 220982 76898 221066 77134
rect 221302 76898 238746 77134
rect 238982 76898 239066 77134
rect 239302 76898 256746 77134
rect 256982 76898 257066 77134
rect 257302 76898 274746 77134
rect 274982 76898 275066 77134
rect 275302 76898 292746 77134
rect 292982 76898 293066 77134
rect 293302 76898 310746 77134
rect 310982 76898 311066 77134
rect 311302 76898 328746 77134
rect 328982 76898 329066 77134
rect 329302 76898 346746 77134
rect 346982 76898 347066 77134
rect 347302 76898 364746 77134
rect 364982 76898 365066 77134
rect 365302 76898 382746 77134
rect 382982 76898 383066 77134
rect 383302 76898 400746 77134
rect 400982 76898 401066 77134
rect 401302 76898 418746 77134
rect 418982 76898 419066 77134
rect 419302 76898 436746 77134
rect 436982 76898 437066 77134
rect 437302 76898 454746 77134
rect 454982 76898 455066 77134
rect 455302 76898 472746 77134
rect 472982 76898 473066 77134
rect 473302 76898 490746 77134
rect 490982 76898 491066 77134
rect 491302 76898 508746 77134
rect 508982 76898 509066 77134
rect 509302 76898 526746 77134
rect 526982 76898 527066 77134
rect 527302 76898 545004 77134
rect 545240 76898 545324 77134
rect 545560 76898 548472 77134
rect -4476 76866 548472 76898
rect -4476 70614 548472 70646
rect -4476 70378 -4444 70614
rect -4208 70378 -4124 70614
rect -3888 70378 15906 70614
rect 16142 70378 16226 70614
rect 16462 70378 33906 70614
rect 34142 70378 34226 70614
rect 34462 70378 51906 70614
rect 52142 70378 52226 70614
rect 52462 70378 69906 70614
rect 70142 70378 70226 70614
rect 70462 70378 87906 70614
rect 88142 70378 88226 70614
rect 88462 70378 105906 70614
rect 106142 70378 106226 70614
rect 106462 70378 123906 70614
rect 124142 70378 124226 70614
rect 124462 70378 141906 70614
rect 142142 70378 142226 70614
rect 142462 70378 159906 70614
rect 160142 70378 160226 70614
rect 160462 70378 177906 70614
rect 178142 70378 178226 70614
rect 178462 70378 195906 70614
rect 196142 70378 196226 70614
rect 196462 70378 213906 70614
rect 214142 70378 214226 70614
rect 214462 70378 231906 70614
rect 232142 70378 232226 70614
rect 232462 70378 249906 70614
rect 250142 70378 250226 70614
rect 250462 70378 267906 70614
rect 268142 70378 268226 70614
rect 268462 70378 285906 70614
rect 286142 70378 286226 70614
rect 286462 70378 303906 70614
rect 304142 70378 304226 70614
rect 304462 70378 321906 70614
rect 322142 70378 322226 70614
rect 322462 70378 339906 70614
rect 340142 70378 340226 70614
rect 340462 70378 357906 70614
rect 358142 70378 358226 70614
rect 358462 70378 375906 70614
rect 376142 70378 376226 70614
rect 376462 70378 393906 70614
rect 394142 70378 394226 70614
rect 394462 70378 411906 70614
rect 412142 70378 412226 70614
rect 412462 70378 429906 70614
rect 430142 70378 430226 70614
rect 430462 70378 447906 70614
rect 448142 70378 448226 70614
rect 448462 70378 465906 70614
rect 466142 70378 466226 70614
rect 466462 70378 483906 70614
rect 484142 70378 484226 70614
rect 484462 70378 501906 70614
rect 502142 70378 502226 70614
rect 502462 70378 519906 70614
rect 520142 70378 520226 70614
rect 520462 70378 537906 70614
rect 538142 70378 538226 70614
rect 538462 70378 547884 70614
rect 548120 70378 548204 70614
rect 548440 70378 548472 70614
rect -4476 70294 548472 70378
rect -4476 70058 -4444 70294
rect -4208 70058 -4124 70294
rect -3888 70058 15906 70294
rect 16142 70058 16226 70294
rect 16462 70058 33906 70294
rect 34142 70058 34226 70294
rect 34462 70058 51906 70294
rect 52142 70058 52226 70294
rect 52462 70058 69906 70294
rect 70142 70058 70226 70294
rect 70462 70058 87906 70294
rect 88142 70058 88226 70294
rect 88462 70058 105906 70294
rect 106142 70058 106226 70294
rect 106462 70058 123906 70294
rect 124142 70058 124226 70294
rect 124462 70058 141906 70294
rect 142142 70058 142226 70294
rect 142462 70058 159906 70294
rect 160142 70058 160226 70294
rect 160462 70058 177906 70294
rect 178142 70058 178226 70294
rect 178462 70058 195906 70294
rect 196142 70058 196226 70294
rect 196462 70058 213906 70294
rect 214142 70058 214226 70294
rect 214462 70058 231906 70294
rect 232142 70058 232226 70294
rect 232462 70058 249906 70294
rect 250142 70058 250226 70294
rect 250462 70058 267906 70294
rect 268142 70058 268226 70294
rect 268462 70058 285906 70294
rect 286142 70058 286226 70294
rect 286462 70058 303906 70294
rect 304142 70058 304226 70294
rect 304462 70058 321906 70294
rect 322142 70058 322226 70294
rect 322462 70058 339906 70294
rect 340142 70058 340226 70294
rect 340462 70058 357906 70294
rect 358142 70058 358226 70294
rect 358462 70058 375906 70294
rect 376142 70058 376226 70294
rect 376462 70058 393906 70294
rect 394142 70058 394226 70294
rect 394462 70058 411906 70294
rect 412142 70058 412226 70294
rect 412462 70058 429906 70294
rect 430142 70058 430226 70294
rect 430462 70058 447906 70294
rect 448142 70058 448226 70294
rect 448462 70058 465906 70294
rect 466142 70058 466226 70294
rect 466462 70058 483906 70294
rect 484142 70058 484226 70294
rect 484462 70058 501906 70294
rect 502142 70058 502226 70294
rect 502462 70058 519906 70294
rect 520142 70058 520226 70294
rect 520462 70058 537906 70294
rect 538142 70058 538226 70294
rect 538462 70058 547884 70294
rect 548120 70058 548204 70294
rect 548440 70058 548472 70294
rect -4476 70026 548472 70058
rect -4476 66894 548472 66926
rect -4476 66658 -3484 66894
rect -3248 66658 -3164 66894
rect -2928 66658 12186 66894
rect 12422 66658 12506 66894
rect 12742 66658 30186 66894
rect 30422 66658 30506 66894
rect 30742 66658 48186 66894
rect 48422 66658 48506 66894
rect 48742 66658 66186 66894
rect 66422 66658 66506 66894
rect 66742 66658 84186 66894
rect 84422 66658 84506 66894
rect 84742 66658 102186 66894
rect 102422 66658 102506 66894
rect 102742 66658 120186 66894
rect 120422 66658 120506 66894
rect 120742 66658 138186 66894
rect 138422 66658 138506 66894
rect 138742 66658 156186 66894
rect 156422 66658 156506 66894
rect 156742 66658 174186 66894
rect 174422 66658 174506 66894
rect 174742 66658 192186 66894
rect 192422 66658 192506 66894
rect 192742 66658 210186 66894
rect 210422 66658 210506 66894
rect 210742 66658 228186 66894
rect 228422 66658 228506 66894
rect 228742 66658 246186 66894
rect 246422 66658 246506 66894
rect 246742 66658 264186 66894
rect 264422 66658 264506 66894
rect 264742 66658 282186 66894
rect 282422 66658 282506 66894
rect 282742 66658 300186 66894
rect 300422 66658 300506 66894
rect 300742 66658 318186 66894
rect 318422 66658 318506 66894
rect 318742 66658 336186 66894
rect 336422 66658 336506 66894
rect 336742 66658 354186 66894
rect 354422 66658 354506 66894
rect 354742 66658 372186 66894
rect 372422 66658 372506 66894
rect 372742 66658 390186 66894
rect 390422 66658 390506 66894
rect 390742 66658 408186 66894
rect 408422 66658 408506 66894
rect 408742 66658 426186 66894
rect 426422 66658 426506 66894
rect 426742 66658 444186 66894
rect 444422 66658 444506 66894
rect 444742 66658 462186 66894
rect 462422 66658 462506 66894
rect 462742 66658 480186 66894
rect 480422 66658 480506 66894
rect 480742 66658 498186 66894
rect 498422 66658 498506 66894
rect 498742 66658 516186 66894
rect 516422 66658 516506 66894
rect 516742 66658 534186 66894
rect 534422 66658 534506 66894
rect 534742 66658 546924 66894
rect 547160 66658 547244 66894
rect 547480 66658 548472 66894
rect -4476 66574 548472 66658
rect -4476 66338 -3484 66574
rect -3248 66338 -3164 66574
rect -2928 66338 12186 66574
rect 12422 66338 12506 66574
rect 12742 66338 30186 66574
rect 30422 66338 30506 66574
rect 30742 66338 48186 66574
rect 48422 66338 48506 66574
rect 48742 66338 66186 66574
rect 66422 66338 66506 66574
rect 66742 66338 84186 66574
rect 84422 66338 84506 66574
rect 84742 66338 102186 66574
rect 102422 66338 102506 66574
rect 102742 66338 120186 66574
rect 120422 66338 120506 66574
rect 120742 66338 138186 66574
rect 138422 66338 138506 66574
rect 138742 66338 156186 66574
rect 156422 66338 156506 66574
rect 156742 66338 174186 66574
rect 174422 66338 174506 66574
rect 174742 66338 192186 66574
rect 192422 66338 192506 66574
rect 192742 66338 210186 66574
rect 210422 66338 210506 66574
rect 210742 66338 228186 66574
rect 228422 66338 228506 66574
rect 228742 66338 246186 66574
rect 246422 66338 246506 66574
rect 246742 66338 264186 66574
rect 264422 66338 264506 66574
rect 264742 66338 282186 66574
rect 282422 66338 282506 66574
rect 282742 66338 300186 66574
rect 300422 66338 300506 66574
rect 300742 66338 318186 66574
rect 318422 66338 318506 66574
rect 318742 66338 336186 66574
rect 336422 66338 336506 66574
rect 336742 66338 354186 66574
rect 354422 66338 354506 66574
rect 354742 66338 372186 66574
rect 372422 66338 372506 66574
rect 372742 66338 390186 66574
rect 390422 66338 390506 66574
rect 390742 66338 408186 66574
rect 408422 66338 408506 66574
rect 408742 66338 426186 66574
rect 426422 66338 426506 66574
rect 426742 66338 444186 66574
rect 444422 66338 444506 66574
rect 444742 66338 462186 66574
rect 462422 66338 462506 66574
rect 462742 66338 480186 66574
rect 480422 66338 480506 66574
rect 480742 66338 498186 66574
rect 498422 66338 498506 66574
rect 498742 66338 516186 66574
rect 516422 66338 516506 66574
rect 516742 66338 534186 66574
rect 534422 66338 534506 66574
rect 534742 66338 546924 66574
rect 547160 66338 547244 66574
rect 547480 66338 548472 66574
rect -4476 66306 548472 66338
rect -4476 63174 548472 63206
rect -4476 62938 -2524 63174
rect -2288 62938 -2204 63174
rect -1968 62938 8466 63174
rect 8702 62938 8786 63174
rect 9022 62938 26466 63174
rect 26702 62938 26786 63174
rect 27022 62938 44466 63174
rect 44702 62938 44786 63174
rect 45022 62938 62466 63174
rect 62702 62938 62786 63174
rect 63022 62938 80466 63174
rect 80702 62938 80786 63174
rect 81022 62938 98466 63174
rect 98702 62938 98786 63174
rect 99022 62938 116466 63174
rect 116702 62938 116786 63174
rect 117022 62938 134466 63174
rect 134702 62938 134786 63174
rect 135022 62938 152466 63174
rect 152702 62938 152786 63174
rect 153022 62938 170466 63174
rect 170702 62938 170786 63174
rect 171022 62938 188466 63174
rect 188702 62938 188786 63174
rect 189022 62938 206466 63174
rect 206702 62938 206786 63174
rect 207022 62938 224466 63174
rect 224702 62938 224786 63174
rect 225022 62938 242466 63174
rect 242702 62938 242786 63174
rect 243022 62938 260466 63174
rect 260702 62938 260786 63174
rect 261022 62938 278466 63174
rect 278702 62938 278786 63174
rect 279022 62938 296466 63174
rect 296702 62938 296786 63174
rect 297022 62938 314466 63174
rect 314702 62938 314786 63174
rect 315022 62938 332466 63174
rect 332702 62938 332786 63174
rect 333022 62938 350466 63174
rect 350702 62938 350786 63174
rect 351022 62938 368466 63174
rect 368702 62938 368786 63174
rect 369022 62938 386466 63174
rect 386702 62938 386786 63174
rect 387022 62938 404466 63174
rect 404702 62938 404786 63174
rect 405022 62938 422466 63174
rect 422702 62938 422786 63174
rect 423022 62938 440466 63174
rect 440702 62938 440786 63174
rect 441022 62938 458466 63174
rect 458702 62938 458786 63174
rect 459022 62938 476466 63174
rect 476702 62938 476786 63174
rect 477022 62938 494466 63174
rect 494702 62938 494786 63174
rect 495022 62938 512466 63174
rect 512702 62938 512786 63174
rect 513022 62938 530466 63174
rect 530702 62938 530786 63174
rect 531022 62938 545964 63174
rect 546200 62938 546284 63174
rect 546520 62938 548472 63174
rect -4476 62854 548472 62938
rect -4476 62618 -2524 62854
rect -2288 62618 -2204 62854
rect -1968 62618 8466 62854
rect 8702 62618 8786 62854
rect 9022 62618 26466 62854
rect 26702 62618 26786 62854
rect 27022 62618 44466 62854
rect 44702 62618 44786 62854
rect 45022 62618 62466 62854
rect 62702 62618 62786 62854
rect 63022 62618 80466 62854
rect 80702 62618 80786 62854
rect 81022 62618 98466 62854
rect 98702 62618 98786 62854
rect 99022 62618 116466 62854
rect 116702 62618 116786 62854
rect 117022 62618 134466 62854
rect 134702 62618 134786 62854
rect 135022 62618 152466 62854
rect 152702 62618 152786 62854
rect 153022 62618 170466 62854
rect 170702 62618 170786 62854
rect 171022 62618 188466 62854
rect 188702 62618 188786 62854
rect 189022 62618 206466 62854
rect 206702 62618 206786 62854
rect 207022 62618 224466 62854
rect 224702 62618 224786 62854
rect 225022 62618 242466 62854
rect 242702 62618 242786 62854
rect 243022 62618 260466 62854
rect 260702 62618 260786 62854
rect 261022 62618 278466 62854
rect 278702 62618 278786 62854
rect 279022 62618 296466 62854
rect 296702 62618 296786 62854
rect 297022 62618 314466 62854
rect 314702 62618 314786 62854
rect 315022 62618 332466 62854
rect 332702 62618 332786 62854
rect 333022 62618 350466 62854
rect 350702 62618 350786 62854
rect 351022 62618 368466 62854
rect 368702 62618 368786 62854
rect 369022 62618 386466 62854
rect 386702 62618 386786 62854
rect 387022 62618 404466 62854
rect 404702 62618 404786 62854
rect 405022 62618 422466 62854
rect 422702 62618 422786 62854
rect 423022 62618 440466 62854
rect 440702 62618 440786 62854
rect 441022 62618 458466 62854
rect 458702 62618 458786 62854
rect 459022 62618 476466 62854
rect 476702 62618 476786 62854
rect 477022 62618 494466 62854
rect 494702 62618 494786 62854
rect 495022 62618 512466 62854
rect 512702 62618 512786 62854
rect 513022 62618 530466 62854
rect 530702 62618 530786 62854
rect 531022 62618 545964 62854
rect 546200 62618 546284 62854
rect 546520 62618 548472 62854
rect -4476 62586 548472 62618
rect 116 60298 118012 60340
rect 116 60062 158 60298
rect 394 60062 117734 60298
rect 117970 60062 118012 60298
rect 116 60020 118012 60062
rect -4476 59454 548472 59486
rect -4476 59218 -1564 59454
rect -1328 59218 -1244 59454
rect -1008 59218 4746 59454
rect 4982 59218 5066 59454
rect 5302 59218 22746 59454
rect 22982 59218 23066 59454
rect 23302 59218 40746 59454
rect 40982 59218 41066 59454
rect 41302 59218 58746 59454
rect 58982 59218 59066 59454
rect 59302 59218 76746 59454
rect 76982 59218 77066 59454
rect 77302 59218 112746 59454
rect 112982 59218 113066 59454
rect 113302 59218 130746 59454
rect 130982 59218 131066 59454
rect 131302 59218 148746 59454
rect 148982 59218 149066 59454
rect 149302 59218 166746 59454
rect 166982 59218 167066 59454
rect 167302 59218 184746 59454
rect 184982 59218 185066 59454
rect 185302 59218 202746 59454
rect 202982 59218 203066 59454
rect 203302 59218 220746 59454
rect 220982 59218 221066 59454
rect 221302 59218 238746 59454
rect 238982 59218 239066 59454
rect 239302 59218 256746 59454
rect 256982 59218 257066 59454
rect 257302 59218 274746 59454
rect 274982 59218 275066 59454
rect 275302 59218 292746 59454
rect 292982 59218 293066 59454
rect 293302 59218 310746 59454
rect 310982 59218 311066 59454
rect 311302 59218 328746 59454
rect 328982 59218 329066 59454
rect 329302 59218 346746 59454
rect 346982 59218 347066 59454
rect 347302 59218 364746 59454
rect 364982 59218 365066 59454
rect 365302 59218 382746 59454
rect 382982 59218 383066 59454
rect 383302 59218 400746 59454
rect 400982 59218 401066 59454
rect 401302 59218 418746 59454
rect 418982 59218 419066 59454
rect 419302 59218 436746 59454
rect 436982 59218 437066 59454
rect 437302 59218 454746 59454
rect 454982 59218 455066 59454
rect 455302 59218 472746 59454
rect 472982 59218 473066 59454
rect 473302 59218 490746 59454
rect 490982 59218 491066 59454
rect 491302 59218 508746 59454
rect 508982 59218 509066 59454
rect 509302 59218 526746 59454
rect 526982 59218 527066 59454
rect 527302 59218 545004 59454
rect 545240 59218 545324 59454
rect 545560 59218 548472 59454
rect -4476 59134 548472 59218
rect -4476 58898 -1564 59134
rect -1328 58898 -1244 59134
rect -1008 58898 4746 59134
rect 4982 58898 5066 59134
rect 5302 58898 22746 59134
rect 22982 58898 23066 59134
rect 23302 58898 40746 59134
rect 40982 58898 41066 59134
rect 41302 58898 58746 59134
rect 58982 58898 59066 59134
rect 59302 58898 76746 59134
rect 76982 58898 77066 59134
rect 77302 58898 112746 59134
rect 112982 58898 113066 59134
rect 113302 58898 130746 59134
rect 130982 58898 131066 59134
rect 131302 58898 148746 59134
rect 148982 58898 149066 59134
rect 149302 58898 166746 59134
rect 166982 58898 167066 59134
rect 167302 58898 184746 59134
rect 184982 58898 185066 59134
rect 185302 58898 202746 59134
rect 202982 58898 203066 59134
rect 203302 58898 220746 59134
rect 220982 58898 221066 59134
rect 221302 58898 238746 59134
rect 238982 58898 239066 59134
rect 239302 58898 256746 59134
rect 256982 58898 257066 59134
rect 257302 58898 274746 59134
rect 274982 58898 275066 59134
rect 275302 58898 292746 59134
rect 292982 58898 293066 59134
rect 293302 58898 310746 59134
rect 310982 58898 311066 59134
rect 311302 58898 328746 59134
rect 328982 58898 329066 59134
rect 329302 58898 346746 59134
rect 346982 58898 347066 59134
rect 347302 58898 364746 59134
rect 364982 58898 365066 59134
rect 365302 58898 382746 59134
rect 382982 58898 383066 59134
rect 383302 58898 400746 59134
rect 400982 58898 401066 59134
rect 401302 58898 418746 59134
rect 418982 58898 419066 59134
rect 419302 58898 436746 59134
rect 436982 58898 437066 59134
rect 437302 58898 454746 59134
rect 454982 58898 455066 59134
rect 455302 58898 472746 59134
rect 472982 58898 473066 59134
rect 473302 58898 490746 59134
rect 490982 58898 491066 59134
rect 491302 58898 508746 59134
rect 508982 58898 509066 59134
rect 509302 58898 526746 59134
rect 526982 58898 527066 59134
rect 527302 58898 545004 59134
rect 545240 58898 545324 59134
rect 545560 58898 548472 59134
rect -4476 58866 548472 58898
rect -4476 52614 548472 52646
rect -4476 52378 -4444 52614
rect -4208 52378 -4124 52614
rect -3888 52378 15906 52614
rect 16142 52378 16226 52614
rect 16462 52378 33906 52614
rect 34142 52378 34226 52614
rect 34462 52378 51906 52614
rect 52142 52378 52226 52614
rect 52462 52378 69906 52614
rect 70142 52378 70226 52614
rect 70462 52378 87906 52614
rect 88142 52378 88226 52614
rect 88462 52378 141906 52614
rect 142142 52378 142226 52614
rect 142462 52378 159906 52614
rect 160142 52378 160226 52614
rect 160462 52378 177906 52614
rect 178142 52378 178226 52614
rect 178462 52378 195906 52614
rect 196142 52378 196226 52614
rect 196462 52378 213906 52614
rect 214142 52378 214226 52614
rect 214462 52378 231906 52614
rect 232142 52378 232226 52614
rect 232462 52378 249906 52614
rect 250142 52378 250226 52614
rect 250462 52378 267906 52614
rect 268142 52378 268226 52614
rect 268462 52378 285906 52614
rect 286142 52378 286226 52614
rect 286462 52378 303906 52614
rect 304142 52378 304226 52614
rect 304462 52378 321906 52614
rect 322142 52378 322226 52614
rect 322462 52378 339906 52614
rect 340142 52378 340226 52614
rect 340462 52378 357906 52614
rect 358142 52378 358226 52614
rect 358462 52378 375906 52614
rect 376142 52378 376226 52614
rect 376462 52378 393906 52614
rect 394142 52378 394226 52614
rect 394462 52378 411906 52614
rect 412142 52378 412226 52614
rect 412462 52378 429906 52614
rect 430142 52378 430226 52614
rect 430462 52378 447906 52614
rect 448142 52378 448226 52614
rect 448462 52378 465906 52614
rect 466142 52378 466226 52614
rect 466462 52378 483906 52614
rect 484142 52378 484226 52614
rect 484462 52378 501906 52614
rect 502142 52378 502226 52614
rect 502462 52378 519906 52614
rect 520142 52378 520226 52614
rect 520462 52378 537906 52614
rect 538142 52378 538226 52614
rect 538462 52378 547884 52614
rect 548120 52378 548204 52614
rect 548440 52378 548472 52614
rect -4476 52294 548472 52378
rect -4476 52058 -4444 52294
rect -4208 52058 -4124 52294
rect -3888 52058 15906 52294
rect 16142 52058 16226 52294
rect 16462 52058 33906 52294
rect 34142 52058 34226 52294
rect 34462 52058 51906 52294
rect 52142 52058 52226 52294
rect 52462 52058 69906 52294
rect 70142 52058 70226 52294
rect 70462 52058 87906 52294
rect 88142 52058 88226 52294
rect 88462 52058 141906 52294
rect 142142 52058 142226 52294
rect 142462 52058 159906 52294
rect 160142 52058 160226 52294
rect 160462 52058 177906 52294
rect 178142 52058 178226 52294
rect 178462 52058 195906 52294
rect 196142 52058 196226 52294
rect 196462 52058 213906 52294
rect 214142 52058 214226 52294
rect 214462 52058 231906 52294
rect 232142 52058 232226 52294
rect 232462 52058 249906 52294
rect 250142 52058 250226 52294
rect 250462 52058 267906 52294
rect 268142 52058 268226 52294
rect 268462 52058 285906 52294
rect 286142 52058 286226 52294
rect 286462 52058 303906 52294
rect 304142 52058 304226 52294
rect 304462 52058 321906 52294
rect 322142 52058 322226 52294
rect 322462 52058 339906 52294
rect 340142 52058 340226 52294
rect 340462 52058 357906 52294
rect 358142 52058 358226 52294
rect 358462 52058 375906 52294
rect 376142 52058 376226 52294
rect 376462 52058 393906 52294
rect 394142 52058 394226 52294
rect 394462 52058 411906 52294
rect 412142 52058 412226 52294
rect 412462 52058 429906 52294
rect 430142 52058 430226 52294
rect 430462 52058 447906 52294
rect 448142 52058 448226 52294
rect 448462 52058 465906 52294
rect 466142 52058 466226 52294
rect 466462 52058 483906 52294
rect 484142 52058 484226 52294
rect 484462 52058 501906 52294
rect 502142 52058 502226 52294
rect 502462 52058 519906 52294
rect 520142 52058 520226 52294
rect 520462 52058 537906 52294
rect 538142 52058 538226 52294
rect 538462 52058 547884 52294
rect 548120 52058 548204 52294
rect 548440 52058 548472 52294
rect -4476 52026 548472 52058
rect -4476 48894 548472 48926
rect -4476 48658 -3484 48894
rect -3248 48658 -3164 48894
rect -2928 48658 12186 48894
rect 12422 48658 12506 48894
rect 12742 48658 30186 48894
rect 30422 48658 30506 48894
rect 30742 48658 48186 48894
rect 48422 48658 48506 48894
rect 48742 48658 66186 48894
rect 66422 48658 66506 48894
rect 66742 48658 84186 48894
rect 84422 48658 84506 48894
rect 84742 48658 138186 48894
rect 138422 48658 138506 48894
rect 138742 48658 174186 48894
rect 174422 48658 174506 48894
rect 174742 48658 192186 48894
rect 192422 48658 192506 48894
rect 192742 48658 210186 48894
rect 210422 48658 210506 48894
rect 210742 48658 228186 48894
rect 228422 48658 228506 48894
rect 228742 48658 246186 48894
rect 246422 48658 246506 48894
rect 246742 48658 264186 48894
rect 264422 48658 264506 48894
rect 264742 48658 282186 48894
rect 282422 48658 282506 48894
rect 282742 48658 300186 48894
rect 300422 48658 300506 48894
rect 300742 48658 318186 48894
rect 318422 48658 318506 48894
rect 318742 48658 336186 48894
rect 336422 48658 336506 48894
rect 336742 48658 354186 48894
rect 354422 48658 354506 48894
rect 354742 48658 372186 48894
rect 372422 48658 372506 48894
rect 372742 48658 390186 48894
rect 390422 48658 390506 48894
rect 390742 48658 408186 48894
rect 408422 48658 408506 48894
rect 408742 48658 426186 48894
rect 426422 48658 426506 48894
rect 426742 48658 444186 48894
rect 444422 48658 444506 48894
rect 444742 48658 462186 48894
rect 462422 48658 462506 48894
rect 462742 48658 480186 48894
rect 480422 48658 480506 48894
rect 480742 48658 498186 48894
rect 498422 48658 498506 48894
rect 498742 48658 516186 48894
rect 516422 48658 516506 48894
rect 516742 48658 534186 48894
rect 534422 48658 534506 48894
rect 534742 48658 546924 48894
rect 547160 48658 547244 48894
rect 547480 48658 548472 48894
rect -4476 48574 548472 48658
rect -4476 48338 -3484 48574
rect -3248 48338 -3164 48574
rect -2928 48338 12186 48574
rect 12422 48338 12506 48574
rect 12742 48338 30186 48574
rect 30422 48338 30506 48574
rect 30742 48338 48186 48574
rect 48422 48338 48506 48574
rect 48742 48338 66186 48574
rect 66422 48338 66506 48574
rect 66742 48338 84186 48574
rect 84422 48338 84506 48574
rect 84742 48338 138186 48574
rect 138422 48338 138506 48574
rect 138742 48338 174186 48574
rect 174422 48338 174506 48574
rect 174742 48338 192186 48574
rect 192422 48338 192506 48574
rect 192742 48338 210186 48574
rect 210422 48338 210506 48574
rect 210742 48338 228186 48574
rect 228422 48338 228506 48574
rect 228742 48338 246186 48574
rect 246422 48338 246506 48574
rect 246742 48338 264186 48574
rect 264422 48338 264506 48574
rect 264742 48338 282186 48574
rect 282422 48338 282506 48574
rect 282742 48338 300186 48574
rect 300422 48338 300506 48574
rect 300742 48338 318186 48574
rect 318422 48338 318506 48574
rect 318742 48338 336186 48574
rect 336422 48338 336506 48574
rect 336742 48338 354186 48574
rect 354422 48338 354506 48574
rect 354742 48338 372186 48574
rect 372422 48338 372506 48574
rect 372742 48338 390186 48574
rect 390422 48338 390506 48574
rect 390742 48338 408186 48574
rect 408422 48338 408506 48574
rect 408742 48338 426186 48574
rect 426422 48338 426506 48574
rect 426742 48338 444186 48574
rect 444422 48338 444506 48574
rect 444742 48338 462186 48574
rect 462422 48338 462506 48574
rect 462742 48338 480186 48574
rect 480422 48338 480506 48574
rect 480742 48338 498186 48574
rect 498422 48338 498506 48574
rect 498742 48338 516186 48574
rect 516422 48338 516506 48574
rect 516742 48338 534186 48574
rect 534422 48338 534506 48574
rect 534742 48338 546924 48574
rect 547160 48338 547244 48574
rect 547480 48338 548472 48574
rect -4476 48306 548472 48338
rect -4476 45174 548472 45206
rect -4476 44938 -2524 45174
rect -2288 44938 -2204 45174
rect -1968 44938 8466 45174
rect 8702 44938 8786 45174
rect 9022 44938 26466 45174
rect 26702 44938 26786 45174
rect 27022 44938 44466 45174
rect 44702 44938 44786 45174
rect 45022 44938 62466 45174
rect 62702 44938 62786 45174
rect 63022 44938 80466 45174
rect 80702 44938 80786 45174
rect 81022 44938 95830 45174
rect 96066 44938 126550 45174
rect 126786 44938 134466 45174
rect 134702 44938 134786 45174
rect 135022 44938 152466 45174
rect 152702 44938 152786 45174
rect 153022 44938 157270 45174
rect 157506 44938 170466 45174
rect 170702 44938 170786 45174
rect 171022 44938 188466 45174
rect 188702 44938 188786 45174
rect 189022 44938 206466 45174
rect 206702 44938 206786 45174
rect 207022 44938 224466 45174
rect 224702 44938 224786 45174
rect 225022 44938 242466 45174
rect 242702 44938 242786 45174
rect 243022 44938 260466 45174
rect 260702 44938 260786 45174
rect 261022 44938 278466 45174
rect 278702 44938 278786 45174
rect 279022 44938 296466 45174
rect 296702 44938 296786 45174
rect 297022 44938 314466 45174
rect 314702 44938 314786 45174
rect 315022 44938 332466 45174
rect 332702 44938 332786 45174
rect 333022 44938 350466 45174
rect 350702 44938 350786 45174
rect 351022 44938 368466 45174
rect 368702 44938 368786 45174
rect 369022 44938 386466 45174
rect 386702 44938 386786 45174
rect 387022 44938 404466 45174
rect 404702 44938 404786 45174
rect 405022 44938 422466 45174
rect 422702 44938 422786 45174
rect 423022 44938 440466 45174
rect 440702 44938 440786 45174
rect 441022 44938 458466 45174
rect 458702 44938 458786 45174
rect 459022 44938 476466 45174
rect 476702 44938 476786 45174
rect 477022 44938 494466 45174
rect 494702 44938 494786 45174
rect 495022 44938 512466 45174
rect 512702 44938 512786 45174
rect 513022 44938 530466 45174
rect 530702 44938 530786 45174
rect 531022 44938 545964 45174
rect 546200 44938 546284 45174
rect 546520 44938 548472 45174
rect -4476 44854 548472 44938
rect -4476 44618 -2524 44854
rect -2288 44618 -2204 44854
rect -1968 44618 8466 44854
rect 8702 44618 8786 44854
rect 9022 44618 26466 44854
rect 26702 44618 26786 44854
rect 27022 44618 44466 44854
rect 44702 44618 44786 44854
rect 45022 44618 62466 44854
rect 62702 44618 62786 44854
rect 63022 44618 80466 44854
rect 80702 44618 80786 44854
rect 81022 44618 95830 44854
rect 96066 44618 126550 44854
rect 126786 44618 134466 44854
rect 134702 44618 134786 44854
rect 135022 44618 152466 44854
rect 152702 44618 152786 44854
rect 153022 44618 157270 44854
rect 157506 44618 170466 44854
rect 170702 44618 170786 44854
rect 171022 44618 188466 44854
rect 188702 44618 188786 44854
rect 189022 44618 206466 44854
rect 206702 44618 206786 44854
rect 207022 44618 224466 44854
rect 224702 44618 224786 44854
rect 225022 44618 242466 44854
rect 242702 44618 242786 44854
rect 243022 44618 260466 44854
rect 260702 44618 260786 44854
rect 261022 44618 278466 44854
rect 278702 44618 278786 44854
rect 279022 44618 296466 44854
rect 296702 44618 296786 44854
rect 297022 44618 314466 44854
rect 314702 44618 314786 44854
rect 315022 44618 332466 44854
rect 332702 44618 332786 44854
rect 333022 44618 350466 44854
rect 350702 44618 350786 44854
rect 351022 44618 368466 44854
rect 368702 44618 368786 44854
rect 369022 44618 386466 44854
rect 386702 44618 386786 44854
rect 387022 44618 404466 44854
rect 404702 44618 404786 44854
rect 405022 44618 422466 44854
rect 422702 44618 422786 44854
rect 423022 44618 440466 44854
rect 440702 44618 440786 44854
rect 441022 44618 458466 44854
rect 458702 44618 458786 44854
rect 459022 44618 476466 44854
rect 476702 44618 476786 44854
rect 477022 44618 494466 44854
rect 494702 44618 494786 44854
rect 495022 44618 512466 44854
rect 512702 44618 512786 44854
rect 513022 44618 530466 44854
rect 530702 44618 530786 44854
rect 531022 44618 545964 44854
rect 546200 44618 546284 44854
rect 546520 44618 548472 44854
rect -4476 44586 548472 44618
rect -4476 41454 548472 41486
rect -4476 41218 -1564 41454
rect -1328 41218 -1244 41454
rect -1008 41218 4746 41454
rect 4982 41218 5066 41454
rect 5302 41218 22746 41454
rect 22982 41218 23066 41454
rect 23302 41218 40746 41454
rect 40982 41218 41066 41454
rect 41302 41218 58746 41454
rect 58982 41218 59066 41454
rect 59302 41218 76746 41454
rect 76982 41218 77066 41454
rect 77302 41218 95170 41454
rect 95406 41218 125890 41454
rect 126126 41218 148746 41454
rect 148982 41218 149066 41454
rect 149302 41218 156610 41454
rect 156846 41218 166746 41454
rect 166982 41218 167066 41454
rect 167302 41218 184746 41454
rect 184982 41218 185066 41454
rect 185302 41218 202746 41454
rect 202982 41218 203066 41454
rect 203302 41218 220746 41454
rect 220982 41218 221066 41454
rect 221302 41218 238746 41454
rect 238982 41218 239066 41454
rect 239302 41218 256746 41454
rect 256982 41218 257066 41454
rect 257302 41218 274746 41454
rect 274982 41218 275066 41454
rect 275302 41218 292746 41454
rect 292982 41218 293066 41454
rect 293302 41218 310746 41454
rect 310982 41218 311066 41454
rect 311302 41218 328746 41454
rect 328982 41218 329066 41454
rect 329302 41218 346746 41454
rect 346982 41218 347066 41454
rect 347302 41218 364746 41454
rect 364982 41218 365066 41454
rect 365302 41218 382746 41454
rect 382982 41218 383066 41454
rect 383302 41218 400746 41454
rect 400982 41218 401066 41454
rect 401302 41218 418746 41454
rect 418982 41218 419066 41454
rect 419302 41218 436746 41454
rect 436982 41218 437066 41454
rect 437302 41218 454746 41454
rect 454982 41218 455066 41454
rect 455302 41218 472746 41454
rect 472982 41218 473066 41454
rect 473302 41218 490746 41454
rect 490982 41218 491066 41454
rect 491302 41218 508746 41454
rect 508982 41218 509066 41454
rect 509302 41218 526746 41454
rect 526982 41218 527066 41454
rect 527302 41218 545004 41454
rect 545240 41218 545324 41454
rect 545560 41218 548472 41454
rect -4476 41134 548472 41218
rect -4476 40898 -1564 41134
rect -1328 40898 -1244 41134
rect -1008 40898 4746 41134
rect 4982 40898 5066 41134
rect 5302 40898 22746 41134
rect 22982 40898 23066 41134
rect 23302 40898 40746 41134
rect 40982 40898 41066 41134
rect 41302 40898 58746 41134
rect 58982 40898 59066 41134
rect 59302 40898 76746 41134
rect 76982 40898 77066 41134
rect 77302 40898 95170 41134
rect 95406 40898 125890 41134
rect 126126 40898 148746 41134
rect 148982 40898 149066 41134
rect 149302 40898 156610 41134
rect 156846 40898 166746 41134
rect 166982 40898 167066 41134
rect 167302 40898 184746 41134
rect 184982 40898 185066 41134
rect 185302 40898 202746 41134
rect 202982 40898 203066 41134
rect 203302 40898 220746 41134
rect 220982 40898 221066 41134
rect 221302 40898 238746 41134
rect 238982 40898 239066 41134
rect 239302 40898 256746 41134
rect 256982 40898 257066 41134
rect 257302 40898 274746 41134
rect 274982 40898 275066 41134
rect 275302 40898 292746 41134
rect 292982 40898 293066 41134
rect 293302 40898 310746 41134
rect 310982 40898 311066 41134
rect 311302 40898 328746 41134
rect 328982 40898 329066 41134
rect 329302 40898 346746 41134
rect 346982 40898 347066 41134
rect 347302 40898 364746 41134
rect 364982 40898 365066 41134
rect 365302 40898 382746 41134
rect 382982 40898 383066 41134
rect 383302 40898 400746 41134
rect 400982 40898 401066 41134
rect 401302 40898 418746 41134
rect 418982 40898 419066 41134
rect 419302 40898 436746 41134
rect 436982 40898 437066 41134
rect 437302 40898 454746 41134
rect 454982 40898 455066 41134
rect 455302 40898 472746 41134
rect 472982 40898 473066 41134
rect 473302 40898 490746 41134
rect 490982 40898 491066 41134
rect 491302 40898 508746 41134
rect 508982 40898 509066 41134
rect 509302 40898 526746 41134
rect 526982 40898 527066 41134
rect 527302 40898 545004 41134
rect 545240 40898 545324 41134
rect 545560 40898 548472 41134
rect -4476 40866 548472 40898
rect -4476 34614 548472 34646
rect -4476 34378 -4444 34614
rect -4208 34378 -4124 34614
rect -3888 34378 15906 34614
rect 16142 34378 16226 34614
rect 16462 34378 33906 34614
rect 34142 34378 34226 34614
rect 34462 34378 51906 34614
rect 52142 34378 52226 34614
rect 52462 34378 69906 34614
rect 70142 34378 70226 34614
rect 70462 34378 87906 34614
rect 88142 34378 88226 34614
rect 88462 34378 141906 34614
rect 142142 34378 142226 34614
rect 142462 34378 159906 34614
rect 160142 34378 160226 34614
rect 160462 34378 177906 34614
rect 178142 34378 178226 34614
rect 178462 34378 195906 34614
rect 196142 34378 196226 34614
rect 196462 34378 213906 34614
rect 214142 34378 214226 34614
rect 214462 34378 231906 34614
rect 232142 34378 232226 34614
rect 232462 34378 249906 34614
rect 250142 34378 250226 34614
rect 250462 34378 267906 34614
rect 268142 34378 268226 34614
rect 268462 34378 285906 34614
rect 286142 34378 286226 34614
rect 286462 34378 303906 34614
rect 304142 34378 304226 34614
rect 304462 34378 321906 34614
rect 322142 34378 322226 34614
rect 322462 34378 339906 34614
rect 340142 34378 340226 34614
rect 340462 34378 357906 34614
rect 358142 34378 358226 34614
rect 358462 34378 375906 34614
rect 376142 34378 376226 34614
rect 376462 34378 393906 34614
rect 394142 34378 394226 34614
rect 394462 34378 411906 34614
rect 412142 34378 412226 34614
rect 412462 34378 429906 34614
rect 430142 34378 430226 34614
rect 430462 34378 447906 34614
rect 448142 34378 448226 34614
rect 448462 34378 465906 34614
rect 466142 34378 466226 34614
rect 466462 34378 483906 34614
rect 484142 34378 484226 34614
rect 484462 34378 501906 34614
rect 502142 34378 502226 34614
rect 502462 34378 519906 34614
rect 520142 34378 520226 34614
rect 520462 34378 537906 34614
rect 538142 34378 538226 34614
rect 538462 34378 547884 34614
rect 548120 34378 548204 34614
rect 548440 34378 548472 34614
rect -4476 34294 548472 34378
rect -4476 34058 -4444 34294
rect -4208 34058 -4124 34294
rect -3888 34058 15906 34294
rect 16142 34058 16226 34294
rect 16462 34058 33906 34294
rect 34142 34058 34226 34294
rect 34462 34058 51906 34294
rect 52142 34058 52226 34294
rect 52462 34058 69906 34294
rect 70142 34058 70226 34294
rect 70462 34058 87906 34294
rect 88142 34058 88226 34294
rect 88462 34058 141906 34294
rect 142142 34058 142226 34294
rect 142462 34058 159906 34294
rect 160142 34058 160226 34294
rect 160462 34058 177906 34294
rect 178142 34058 178226 34294
rect 178462 34058 195906 34294
rect 196142 34058 196226 34294
rect 196462 34058 213906 34294
rect 214142 34058 214226 34294
rect 214462 34058 231906 34294
rect 232142 34058 232226 34294
rect 232462 34058 249906 34294
rect 250142 34058 250226 34294
rect 250462 34058 267906 34294
rect 268142 34058 268226 34294
rect 268462 34058 285906 34294
rect 286142 34058 286226 34294
rect 286462 34058 303906 34294
rect 304142 34058 304226 34294
rect 304462 34058 321906 34294
rect 322142 34058 322226 34294
rect 322462 34058 339906 34294
rect 340142 34058 340226 34294
rect 340462 34058 357906 34294
rect 358142 34058 358226 34294
rect 358462 34058 375906 34294
rect 376142 34058 376226 34294
rect 376462 34058 393906 34294
rect 394142 34058 394226 34294
rect 394462 34058 411906 34294
rect 412142 34058 412226 34294
rect 412462 34058 429906 34294
rect 430142 34058 430226 34294
rect 430462 34058 447906 34294
rect 448142 34058 448226 34294
rect 448462 34058 465906 34294
rect 466142 34058 466226 34294
rect 466462 34058 483906 34294
rect 484142 34058 484226 34294
rect 484462 34058 501906 34294
rect 502142 34058 502226 34294
rect 502462 34058 519906 34294
rect 520142 34058 520226 34294
rect 520462 34058 537906 34294
rect 538142 34058 538226 34294
rect 538462 34058 547884 34294
rect 548120 34058 548204 34294
rect 548440 34058 548472 34294
rect -4476 34026 548472 34058
rect -4476 30894 101780 30926
rect -4476 30658 -3484 30894
rect -3248 30658 -3164 30894
rect -2928 30658 12186 30894
rect 12422 30658 12506 30894
rect 12742 30658 30186 30894
rect 30422 30658 30506 30894
rect 30742 30658 48186 30894
rect 48422 30658 48506 30894
rect 48742 30658 66186 30894
rect 66422 30658 66506 30894
rect 66742 30658 84186 30894
rect 84422 30658 84506 30894
rect 84742 30658 101780 30894
rect -4476 30574 101780 30658
rect -4476 30338 -3484 30574
rect -3248 30338 -3164 30574
rect -2928 30338 12186 30574
rect 12422 30338 12506 30574
rect 12742 30338 30186 30574
rect 30422 30338 30506 30574
rect 30742 30338 48186 30574
rect 48422 30338 48506 30574
rect 48742 30338 66186 30574
rect 66422 30338 66506 30574
rect 66742 30338 84186 30574
rect 84422 30338 84506 30574
rect 84742 30338 101780 30574
rect -4476 30306 101780 30338
rect 133972 30894 548472 30926
rect 133972 30658 138186 30894
rect 138422 30658 138506 30894
rect 138742 30658 174186 30894
rect 174422 30658 174506 30894
rect 174742 30658 192186 30894
rect 192422 30658 192506 30894
rect 192742 30658 210186 30894
rect 210422 30658 210506 30894
rect 210742 30658 228186 30894
rect 228422 30658 228506 30894
rect 228742 30658 246186 30894
rect 246422 30658 246506 30894
rect 246742 30658 264186 30894
rect 264422 30658 264506 30894
rect 264742 30658 282186 30894
rect 282422 30658 282506 30894
rect 282742 30658 300186 30894
rect 300422 30658 300506 30894
rect 300742 30658 318186 30894
rect 318422 30658 318506 30894
rect 318742 30658 336186 30894
rect 336422 30658 336506 30894
rect 336742 30658 354186 30894
rect 354422 30658 354506 30894
rect 354742 30658 372186 30894
rect 372422 30658 372506 30894
rect 372742 30658 390186 30894
rect 390422 30658 390506 30894
rect 390742 30658 408186 30894
rect 408422 30658 408506 30894
rect 408742 30658 426186 30894
rect 426422 30658 426506 30894
rect 426742 30658 444186 30894
rect 444422 30658 444506 30894
rect 444742 30658 462186 30894
rect 462422 30658 462506 30894
rect 462742 30658 480186 30894
rect 480422 30658 480506 30894
rect 480742 30658 498186 30894
rect 498422 30658 498506 30894
rect 498742 30658 516186 30894
rect 516422 30658 516506 30894
rect 516742 30658 534186 30894
rect 534422 30658 534506 30894
rect 534742 30658 546924 30894
rect 547160 30658 547244 30894
rect 547480 30658 548472 30894
rect 133972 30574 548472 30658
rect 133972 30338 138186 30574
rect 138422 30338 138506 30574
rect 138742 30338 174186 30574
rect 174422 30338 174506 30574
rect 174742 30338 192186 30574
rect 192422 30338 192506 30574
rect 192742 30338 210186 30574
rect 210422 30338 210506 30574
rect 210742 30338 228186 30574
rect 228422 30338 228506 30574
rect 228742 30338 246186 30574
rect 246422 30338 246506 30574
rect 246742 30338 264186 30574
rect 264422 30338 264506 30574
rect 264742 30338 282186 30574
rect 282422 30338 282506 30574
rect 282742 30338 300186 30574
rect 300422 30338 300506 30574
rect 300742 30338 318186 30574
rect 318422 30338 318506 30574
rect 318742 30338 336186 30574
rect 336422 30338 336506 30574
rect 336742 30338 354186 30574
rect 354422 30338 354506 30574
rect 354742 30338 372186 30574
rect 372422 30338 372506 30574
rect 372742 30338 390186 30574
rect 390422 30338 390506 30574
rect 390742 30338 408186 30574
rect 408422 30338 408506 30574
rect 408742 30338 426186 30574
rect 426422 30338 426506 30574
rect 426742 30338 444186 30574
rect 444422 30338 444506 30574
rect 444742 30338 462186 30574
rect 462422 30338 462506 30574
rect 462742 30338 480186 30574
rect 480422 30338 480506 30574
rect 480742 30338 498186 30574
rect 498422 30338 498506 30574
rect 498742 30338 516186 30574
rect 516422 30338 516506 30574
rect 516742 30338 534186 30574
rect 534422 30338 534506 30574
rect 534742 30338 546924 30574
rect 547160 30338 547244 30574
rect 547480 30338 548472 30574
rect 133972 30306 548472 30338
rect -4476 27174 101780 27206
rect -4476 26938 -2524 27174
rect -2288 26938 -2204 27174
rect -1968 26938 8466 27174
rect 8702 26938 8786 27174
rect 9022 26938 26466 27174
rect 26702 26938 26786 27174
rect 27022 26938 44466 27174
rect 44702 26938 44786 27174
rect 45022 26938 62466 27174
rect 62702 26938 62786 27174
rect 63022 26938 80466 27174
rect 80702 26938 80786 27174
rect 81022 26938 95830 27174
rect 96066 26938 101780 27174
rect -4476 26854 101780 26938
rect -4476 26618 -2524 26854
rect -2288 26618 -2204 26854
rect -1968 26618 8466 26854
rect 8702 26618 8786 26854
rect 9022 26618 26466 26854
rect 26702 26618 26786 26854
rect 27022 26618 44466 26854
rect 44702 26618 44786 26854
rect 45022 26618 62466 26854
rect 62702 26618 62786 26854
rect 63022 26618 80466 26854
rect 80702 26618 80786 26854
rect 81022 26618 95830 26854
rect 96066 26618 101780 26854
rect -4476 26586 101780 26618
rect 133972 27174 548472 27206
rect 133972 26938 134466 27174
rect 134702 26938 134786 27174
rect 135022 26938 152466 27174
rect 152702 26938 152786 27174
rect 153022 26938 157270 27174
rect 157506 26938 170466 27174
rect 170702 26938 170786 27174
rect 171022 26938 188466 27174
rect 188702 26938 188786 27174
rect 189022 26938 206466 27174
rect 206702 26938 206786 27174
rect 207022 26938 224466 27174
rect 224702 26938 224786 27174
rect 225022 26938 242466 27174
rect 242702 26938 242786 27174
rect 243022 26938 260466 27174
rect 260702 26938 260786 27174
rect 261022 26938 278466 27174
rect 278702 26938 278786 27174
rect 279022 26938 296466 27174
rect 296702 26938 296786 27174
rect 297022 26938 314466 27174
rect 314702 26938 314786 27174
rect 315022 26938 332466 27174
rect 332702 26938 332786 27174
rect 333022 26938 350466 27174
rect 350702 26938 350786 27174
rect 351022 26938 368466 27174
rect 368702 26938 368786 27174
rect 369022 26938 386466 27174
rect 386702 26938 386786 27174
rect 387022 26938 404466 27174
rect 404702 26938 404786 27174
rect 405022 26938 422466 27174
rect 422702 26938 422786 27174
rect 423022 26938 440466 27174
rect 440702 26938 440786 27174
rect 441022 26938 458466 27174
rect 458702 26938 458786 27174
rect 459022 26938 476466 27174
rect 476702 26938 476786 27174
rect 477022 26938 494466 27174
rect 494702 26938 494786 27174
rect 495022 26938 512466 27174
rect 512702 26938 512786 27174
rect 513022 26938 530466 27174
rect 530702 26938 530786 27174
rect 531022 26938 545964 27174
rect 546200 26938 546284 27174
rect 546520 26938 548472 27174
rect 133972 26854 548472 26938
rect 133972 26618 134466 26854
rect 134702 26618 134786 26854
rect 135022 26618 152466 26854
rect 152702 26618 152786 26854
rect 153022 26618 157270 26854
rect 157506 26618 170466 26854
rect 170702 26618 170786 26854
rect 171022 26618 188466 26854
rect 188702 26618 188786 26854
rect 189022 26618 206466 26854
rect 206702 26618 206786 26854
rect 207022 26618 224466 26854
rect 224702 26618 224786 26854
rect 225022 26618 242466 26854
rect 242702 26618 242786 26854
rect 243022 26618 260466 26854
rect 260702 26618 260786 26854
rect 261022 26618 278466 26854
rect 278702 26618 278786 26854
rect 279022 26618 296466 26854
rect 296702 26618 296786 26854
rect 297022 26618 314466 26854
rect 314702 26618 314786 26854
rect 315022 26618 332466 26854
rect 332702 26618 332786 26854
rect 333022 26618 350466 26854
rect 350702 26618 350786 26854
rect 351022 26618 368466 26854
rect 368702 26618 368786 26854
rect 369022 26618 386466 26854
rect 386702 26618 386786 26854
rect 387022 26618 404466 26854
rect 404702 26618 404786 26854
rect 405022 26618 422466 26854
rect 422702 26618 422786 26854
rect 423022 26618 440466 26854
rect 440702 26618 440786 26854
rect 441022 26618 458466 26854
rect 458702 26618 458786 26854
rect 459022 26618 476466 26854
rect 476702 26618 476786 26854
rect 477022 26618 494466 26854
rect 494702 26618 494786 26854
rect 495022 26618 512466 26854
rect 512702 26618 512786 26854
rect 513022 26618 530466 26854
rect 530702 26618 530786 26854
rect 531022 26618 545964 26854
rect 546200 26618 546284 26854
rect 546520 26618 548472 26854
rect 133972 26586 548472 26618
rect -4476 23454 101780 23486
rect -4476 23218 -1564 23454
rect -1328 23218 -1244 23454
rect -1008 23218 4746 23454
rect 4982 23218 5066 23454
rect 5302 23218 22746 23454
rect 22982 23218 23066 23454
rect 23302 23218 40746 23454
rect 40982 23218 41066 23454
rect 41302 23218 58746 23454
rect 58982 23218 59066 23454
rect 59302 23218 76746 23454
rect 76982 23218 77066 23454
rect 77302 23218 95170 23454
rect 95406 23218 101780 23454
rect -4476 23134 101780 23218
rect -4476 22898 -1564 23134
rect -1328 22898 -1244 23134
rect -1008 22898 4746 23134
rect 4982 22898 5066 23134
rect 5302 22898 22746 23134
rect 22982 22898 23066 23134
rect 23302 22898 40746 23134
rect 40982 22898 41066 23134
rect 41302 22898 58746 23134
rect 58982 22898 59066 23134
rect 59302 22898 76746 23134
rect 76982 22898 77066 23134
rect 77302 22898 95170 23134
rect 95406 22898 101780 23134
rect -4476 22866 101780 22898
rect 133972 23454 548472 23486
rect 133972 23218 148746 23454
rect 148982 23218 149066 23454
rect 149302 23218 156610 23454
rect 156846 23218 166746 23454
rect 166982 23218 167066 23454
rect 167302 23218 184746 23454
rect 184982 23218 185066 23454
rect 185302 23218 202746 23454
rect 202982 23218 203066 23454
rect 203302 23218 220746 23454
rect 220982 23218 221066 23454
rect 221302 23218 238746 23454
rect 238982 23218 239066 23454
rect 239302 23218 256746 23454
rect 256982 23218 257066 23454
rect 257302 23218 274746 23454
rect 274982 23218 275066 23454
rect 275302 23218 292746 23454
rect 292982 23218 293066 23454
rect 293302 23218 310746 23454
rect 310982 23218 311066 23454
rect 311302 23218 328746 23454
rect 328982 23218 329066 23454
rect 329302 23218 346746 23454
rect 346982 23218 347066 23454
rect 347302 23218 364746 23454
rect 364982 23218 365066 23454
rect 365302 23218 382746 23454
rect 382982 23218 383066 23454
rect 383302 23218 400746 23454
rect 400982 23218 401066 23454
rect 401302 23218 418746 23454
rect 418982 23218 419066 23454
rect 419302 23218 436746 23454
rect 436982 23218 437066 23454
rect 437302 23218 454746 23454
rect 454982 23218 455066 23454
rect 455302 23218 472746 23454
rect 472982 23218 473066 23454
rect 473302 23218 490746 23454
rect 490982 23218 491066 23454
rect 491302 23218 508746 23454
rect 508982 23218 509066 23454
rect 509302 23218 526746 23454
rect 526982 23218 527066 23454
rect 527302 23218 545004 23454
rect 545240 23218 545324 23454
rect 545560 23218 548472 23454
rect 133972 23134 548472 23218
rect 133972 22898 148746 23134
rect 148982 22898 149066 23134
rect 149302 22898 156610 23134
rect 156846 22898 166746 23134
rect 166982 22898 167066 23134
rect 167302 22898 184746 23134
rect 184982 22898 185066 23134
rect 185302 22898 202746 23134
rect 202982 22898 203066 23134
rect 203302 22898 220746 23134
rect 220982 22898 221066 23134
rect 221302 22898 238746 23134
rect 238982 22898 239066 23134
rect 239302 22898 256746 23134
rect 256982 22898 257066 23134
rect 257302 22898 274746 23134
rect 274982 22898 275066 23134
rect 275302 22898 292746 23134
rect 292982 22898 293066 23134
rect 293302 22898 310746 23134
rect 310982 22898 311066 23134
rect 311302 22898 328746 23134
rect 328982 22898 329066 23134
rect 329302 22898 346746 23134
rect 346982 22898 347066 23134
rect 347302 22898 364746 23134
rect 364982 22898 365066 23134
rect 365302 22898 382746 23134
rect 382982 22898 383066 23134
rect 383302 22898 400746 23134
rect 400982 22898 401066 23134
rect 401302 22898 418746 23134
rect 418982 22898 419066 23134
rect 419302 22898 436746 23134
rect 436982 22898 437066 23134
rect 437302 22898 454746 23134
rect 454982 22898 455066 23134
rect 455302 22898 472746 23134
rect 472982 22898 473066 23134
rect 473302 22898 490746 23134
rect 490982 22898 491066 23134
rect 491302 22898 508746 23134
rect 508982 22898 509066 23134
rect 509302 22898 526746 23134
rect 526982 22898 527066 23134
rect 527302 22898 545004 23134
rect 545240 22898 545324 23134
rect 545560 22898 548472 23134
rect 133972 22866 548472 22898
rect -4476 16614 548472 16646
rect -4476 16378 -4444 16614
rect -4208 16378 -4124 16614
rect -3888 16378 15906 16614
rect 16142 16378 16226 16614
rect 16462 16378 33906 16614
rect 34142 16378 34226 16614
rect 34462 16378 51906 16614
rect 52142 16378 52226 16614
rect 52462 16378 69906 16614
rect 70142 16378 70226 16614
rect 70462 16378 87906 16614
rect 88142 16378 88226 16614
rect 88462 16378 105906 16614
rect 106142 16378 106226 16614
rect 106462 16378 123906 16614
rect 124142 16378 124226 16614
rect 124462 16378 141906 16614
rect 142142 16378 142226 16614
rect 142462 16378 159906 16614
rect 160142 16378 160226 16614
rect 160462 16378 177906 16614
rect 178142 16378 178226 16614
rect 178462 16378 195906 16614
rect 196142 16378 196226 16614
rect 196462 16378 213906 16614
rect 214142 16378 214226 16614
rect 214462 16378 231906 16614
rect 232142 16378 232226 16614
rect 232462 16378 249906 16614
rect 250142 16378 250226 16614
rect 250462 16378 267906 16614
rect 268142 16378 268226 16614
rect 268462 16378 285906 16614
rect 286142 16378 286226 16614
rect 286462 16378 303906 16614
rect 304142 16378 304226 16614
rect 304462 16378 321906 16614
rect 322142 16378 322226 16614
rect 322462 16378 339906 16614
rect 340142 16378 340226 16614
rect 340462 16378 357906 16614
rect 358142 16378 358226 16614
rect 358462 16378 375906 16614
rect 376142 16378 376226 16614
rect 376462 16378 393906 16614
rect 394142 16378 394226 16614
rect 394462 16378 411906 16614
rect 412142 16378 412226 16614
rect 412462 16378 429906 16614
rect 430142 16378 430226 16614
rect 430462 16378 447906 16614
rect 448142 16378 448226 16614
rect 448462 16378 465906 16614
rect 466142 16378 466226 16614
rect 466462 16378 483906 16614
rect 484142 16378 484226 16614
rect 484462 16378 501906 16614
rect 502142 16378 502226 16614
rect 502462 16378 519906 16614
rect 520142 16378 520226 16614
rect 520462 16378 537906 16614
rect 538142 16378 538226 16614
rect 538462 16378 547884 16614
rect 548120 16378 548204 16614
rect 548440 16378 548472 16614
rect -4476 16294 548472 16378
rect -4476 16058 -4444 16294
rect -4208 16058 -4124 16294
rect -3888 16058 15906 16294
rect 16142 16058 16226 16294
rect 16462 16058 33906 16294
rect 34142 16058 34226 16294
rect 34462 16058 51906 16294
rect 52142 16058 52226 16294
rect 52462 16058 69906 16294
rect 70142 16058 70226 16294
rect 70462 16058 87906 16294
rect 88142 16058 88226 16294
rect 88462 16058 105906 16294
rect 106142 16058 106226 16294
rect 106462 16058 123906 16294
rect 124142 16058 124226 16294
rect 124462 16058 141906 16294
rect 142142 16058 142226 16294
rect 142462 16058 159906 16294
rect 160142 16058 160226 16294
rect 160462 16058 177906 16294
rect 178142 16058 178226 16294
rect 178462 16058 195906 16294
rect 196142 16058 196226 16294
rect 196462 16058 213906 16294
rect 214142 16058 214226 16294
rect 214462 16058 231906 16294
rect 232142 16058 232226 16294
rect 232462 16058 249906 16294
rect 250142 16058 250226 16294
rect 250462 16058 267906 16294
rect 268142 16058 268226 16294
rect 268462 16058 285906 16294
rect 286142 16058 286226 16294
rect 286462 16058 303906 16294
rect 304142 16058 304226 16294
rect 304462 16058 321906 16294
rect 322142 16058 322226 16294
rect 322462 16058 339906 16294
rect 340142 16058 340226 16294
rect 340462 16058 357906 16294
rect 358142 16058 358226 16294
rect 358462 16058 375906 16294
rect 376142 16058 376226 16294
rect 376462 16058 393906 16294
rect 394142 16058 394226 16294
rect 394462 16058 411906 16294
rect 412142 16058 412226 16294
rect 412462 16058 429906 16294
rect 430142 16058 430226 16294
rect 430462 16058 447906 16294
rect 448142 16058 448226 16294
rect 448462 16058 465906 16294
rect 466142 16058 466226 16294
rect 466462 16058 483906 16294
rect 484142 16058 484226 16294
rect 484462 16058 501906 16294
rect 502142 16058 502226 16294
rect 502462 16058 519906 16294
rect 520142 16058 520226 16294
rect 520462 16058 537906 16294
rect 538142 16058 538226 16294
rect 538462 16058 547884 16294
rect 548120 16058 548204 16294
rect 548440 16058 548472 16294
rect -4476 16026 548472 16058
rect -4476 12894 548472 12926
rect -4476 12658 -3484 12894
rect -3248 12658 -3164 12894
rect -2928 12658 12186 12894
rect 12422 12658 12506 12894
rect 12742 12658 30186 12894
rect 30422 12658 30506 12894
rect 30742 12658 48186 12894
rect 48422 12658 48506 12894
rect 48742 12658 66186 12894
rect 66422 12658 66506 12894
rect 66742 12658 84186 12894
rect 84422 12658 84506 12894
rect 84742 12658 102186 12894
rect 102422 12658 102506 12894
rect 102742 12658 120186 12894
rect 120422 12658 120506 12894
rect 120742 12658 138186 12894
rect 138422 12658 138506 12894
rect 138742 12658 156186 12894
rect 156422 12658 156506 12894
rect 156742 12658 174186 12894
rect 174422 12658 174506 12894
rect 174742 12658 192186 12894
rect 192422 12658 192506 12894
rect 192742 12658 210186 12894
rect 210422 12658 210506 12894
rect 210742 12658 228186 12894
rect 228422 12658 228506 12894
rect 228742 12658 246186 12894
rect 246422 12658 246506 12894
rect 246742 12658 264186 12894
rect 264422 12658 264506 12894
rect 264742 12658 282186 12894
rect 282422 12658 282506 12894
rect 282742 12658 300186 12894
rect 300422 12658 300506 12894
rect 300742 12658 318186 12894
rect 318422 12658 318506 12894
rect 318742 12658 336186 12894
rect 336422 12658 336506 12894
rect 336742 12658 354186 12894
rect 354422 12658 354506 12894
rect 354742 12658 372186 12894
rect 372422 12658 372506 12894
rect 372742 12658 390186 12894
rect 390422 12658 390506 12894
rect 390742 12658 408186 12894
rect 408422 12658 408506 12894
rect 408742 12658 426186 12894
rect 426422 12658 426506 12894
rect 426742 12658 444186 12894
rect 444422 12658 444506 12894
rect 444742 12658 462186 12894
rect 462422 12658 462506 12894
rect 462742 12658 480186 12894
rect 480422 12658 480506 12894
rect 480742 12658 498186 12894
rect 498422 12658 498506 12894
rect 498742 12658 516186 12894
rect 516422 12658 516506 12894
rect 516742 12658 534186 12894
rect 534422 12658 534506 12894
rect 534742 12658 546924 12894
rect 547160 12658 547244 12894
rect 547480 12658 548472 12894
rect -4476 12574 548472 12658
rect -4476 12338 -3484 12574
rect -3248 12338 -3164 12574
rect -2928 12338 12186 12574
rect 12422 12338 12506 12574
rect 12742 12338 30186 12574
rect 30422 12338 30506 12574
rect 30742 12338 48186 12574
rect 48422 12338 48506 12574
rect 48742 12338 66186 12574
rect 66422 12338 66506 12574
rect 66742 12338 84186 12574
rect 84422 12338 84506 12574
rect 84742 12338 102186 12574
rect 102422 12338 102506 12574
rect 102742 12338 120186 12574
rect 120422 12338 120506 12574
rect 120742 12338 138186 12574
rect 138422 12338 138506 12574
rect 138742 12338 156186 12574
rect 156422 12338 156506 12574
rect 156742 12338 174186 12574
rect 174422 12338 174506 12574
rect 174742 12338 192186 12574
rect 192422 12338 192506 12574
rect 192742 12338 210186 12574
rect 210422 12338 210506 12574
rect 210742 12338 228186 12574
rect 228422 12338 228506 12574
rect 228742 12338 246186 12574
rect 246422 12338 246506 12574
rect 246742 12338 264186 12574
rect 264422 12338 264506 12574
rect 264742 12338 282186 12574
rect 282422 12338 282506 12574
rect 282742 12338 300186 12574
rect 300422 12338 300506 12574
rect 300742 12338 318186 12574
rect 318422 12338 318506 12574
rect 318742 12338 336186 12574
rect 336422 12338 336506 12574
rect 336742 12338 354186 12574
rect 354422 12338 354506 12574
rect 354742 12338 372186 12574
rect 372422 12338 372506 12574
rect 372742 12338 390186 12574
rect 390422 12338 390506 12574
rect 390742 12338 408186 12574
rect 408422 12338 408506 12574
rect 408742 12338 426186 12574
rect 426422 12338 426506 12574
rect 426742 12338 444186 12574
rect 444422 12338 444506 12574
rect 444742 12338 462186 12574
rect 462422 12338 462506 12574
rect 462742 12338 480186 12574
rect 480422 12338 480506 12574
rect 480742 12338 498186 12574
rect 498422 12338 498506 12574
rect 498742 12338 516186 12574
rect 516422 12338 516506 12574
rect 516742 12338 534186 12574
rect 534422 12338 534506 12574
rect 534742 12338 546924 12574
rect 547160 12338 547244 12574
rect 547480 12338 548472 12574
rect -4476 12306 548472 12338
rect -4476 9174 548472 9206
rect -4476 8938 -2524 9174
rect -2288 8938 -2204 9174
rect -1968 8938 8466 9174
rect 8702 8938 8786 9174
rect 9022 8938 26466 9174
rect 26702 8938 26786 9174
rect 27022 8938 44466 9174
rect 44702 8938 44786 9174
rect 45022 8938 62466 9174
rect 62702 8938 62786 9174
rect 63022 8938 80466 9174
rect 80702 8938 80786 9174
rect 81022 8938 98466 9174
rect 98702 8938 98786 9174
rect 99022 8938 116466 9174
rect 116702 8938 116786 9174
rect 117022 8938 134466 9174
rect 134702 8938 134786 9174
rect 135022 8938 152466 9174
rect 152702 8938 152786 9174
rect 153022 8938 170466 9174
rect 170702 8938 170786 9174
rect 171022 8938 188466 9174
rect 188702 8938 188786 9174
rect 189022 8938 206466 9174
rect 206702 8938 206786 9174
rect 207022 8938 224466 9174
rect 224702 8938 224786 9174
rect 225022 8938 242466 9174
rect 242702 8938 242786 9174
rect 243022 8938 260466 9174
rect 260702 8938 260786 9174
rect 261022 8938 278466 9174
rect 278702 8938 278786 9174
rect 279022 8938 296466 9174
rect 296702 8938 296786 9174
rect 297022 8938 314466 9174
rect 314702 8938 314786 9174
rect 315022 8938 332466 9174
rect 332702 8938 332786 9174
rect 333022 8938 350466 9174
rect 350702 8938 350786 9174
rect 351022 8938 368466 9174
rect 368702 8938 368786 9174
rect 369022 8938 386466 9174
rect 386702 8938 386786 9174
rect 387022 8938 404466 9174
rect 404702 8938 404786 9174
rect 405022 8938 422466 9174
rect 422702 8938 422786 9174
rect 423022 8938 440466 9174
rect 440702 8938 440786 9174
rect 441022 8938 458466 9174
rect 458702 8938 458786 9174
rect 459022 8938 476466 9174
rect 476702 8938 476786 9174
rect 477022 8938 494466 9174
rect 494702 8938 494786 9174
rect 495022 8938 512466 9174
rect 512702 8938 512786 9174
rect 513022 8938 530466 9174
rect 530702 8938 530786 9174
rect 531022 8938 545964 9174
rect 546200 8938 546284 9174
rect 546520 8938 548472 9174
rect -4476 8854 548472 8938
rect -4476 8618 -2524 8854
rect -2288 8618 -2204 8854
rect -1968 8618 8466 8854
rect 8702 8618 8786 8854
rect 9022 8618 26466 8854
rect 26702 8618 26786 8854
rect 27022 8618 44466 8854
rect 44702 8618 44786 8854
rect 45022 8618 62466 8854
rect 62702 8618 62786 8854
rect 63022 8618 80466 8854
rect 80702 8618 80786 8854
rect 81022 8618 98466 8854
rect 98702 8618 98786 8854
rect 99022 8618 116466 8854
rect 116702 8618 116786 8854
rect 117022 8618 134466 8854
rect 134702 8618 134786 8854
rect 135022 8618 152466 8854
rect 152702 8618 152786 8854
rect 153022 8618 170466 8854
rect 170702 8618 170786 8854
rect 171022 8618 188466 8854
rect 188702 8618 188786 8854
rect 189022 8618 206466 8854
rect 206702 8618 206786 8854
rect 207022 8618 224466 8854
rect 224702 8618 224786 8854
rect 225022 8618 242466 8854
rect 242702 8618 242786 8854
rect 243022 8618 260466 8854
rect 260702 8618 260786 8854
rect 261022 8618 278466 8854
rect 278702 8618 278786 8854
rect 279022 8618 296466 8854
rect 296702 8618 296786 8854
rect 297022 8618 314466 8854
rect 314702 8618 314786 8854
rect 315022 8618 332466 8854
rect 332702 8618 332786 8854
rect 333022 8618 350466 8854
rect 350702 8618 350786 8854
rect 351022 8618 368466 8854
rect 368702 8618 368786 8854
rect 369022 8618 386466 8854
rect 386702 8618 386786 8854
rect 387022 8618 404466 8854
rect 404702 8618 404786 8854
rect 405022 8618 422466 8854
rect 422702 8618 422786 8854
rect 423022 8618 440466 8854
rect 440702 8618 440786 8854
rect 441022 8618 458466 8854
rect 458702 8618 458786 8854
rect 459022 8618 476466 8854
rect 476702 8618 476786 8854
rect 477022 8618 494466 8854
rect 494702 8618 494786 8854
rect 495022 8618 512466 8854
rect 512702 8618 512786 8854
rect 513022 8618 530466 8854
rect 530702 8618 530786 8854
rect 531022 8618 545964 8854
rect 546200 8618 546284 8854
rect 546520 8618 548472 8854
rect -4476 8586 548472 8618
rect -4476 5454 548472 5486
rect -4476 5218 -1564 5454
rect -1328 5218 -1244 5454
rect -1008 5218 4746 5454
rect 4982 5218 5066 5454
rect 5302 5218 22746 5454
rect 22982 5218 23066 5454
rect 23302 5218 40746 5454
rect 40982 5218 41066 5454
rect 41302 5218 58746 5454
rect 58982 5218 59066 5454
rect 59302 5218 76746 5454
rect 76982 5218 77066 5454
rect 77302 5218 94746 5454
rect 94982 5218 95066 5454
rect 95302 5218 112746 5454
rect 112982 5218 113066 5454
rect 113302 5218 130746 5454
rect 130982 5218 131066 5454
rect 131302 5218 148746 5454
rect 148982 5218 149066 5454
rect 149302 5218 166746 5454
rect 166982 5218 167066 5454
rect 167302 5218 184746 5454
rect 184982 5218 185066 5454
rect 185302 5218 202746 5454
rect 202982 5218 203066 5454
rect 203302 5218 220746 5454
rect 220982 5218 221066 5454
rect 221302 5218 238746 5454
rect 238982 5218 239066 5454
rect 239302 5218 256746 5454
rect 256982 5218 257066 5454
rect 257302 5218 274746 5454
rect 274982 5218 275066 5454
rect 275302 5218 292746 5454
rect 292982 5218 293066 5454
rect 293302 5218 310746 5454
rect 310982 5218 311066 5454
rect 311302 5218 328746 5454
rect 328982 5218 329066 5454
rect 329302 5218 346746 5454
rect 346982 5218 347066 5454
rect 347302 5218 364746 5454
rect 364982 5218 365066 5454
rect 365302 5218 382746 5454
rect 382982 5218 383066 5454
rect 383302 5218 400746 5454
rect 400982 5218 401066 5454
rect 401302 5218 418746 5454
rect 418982 5218 419066 5454
rect 419302 5218 436746 5454
rect 436982 5218 437066 5454
rect 437302 5218 454746 5454
rect 454982 5218 455066 5454
rect 455302 5218 472746 5454
rect 472982 5218 473066 5454
rect 473302 5218 490746 5454
rect 490982 5218 491066 5454
rect 491302 5218 508746 5454
rect 508982 5218 509066 5454
rect 509302 5218 526746 5454
rect 526982 5218 527066 5454
rect 527302 5218 545004 5454
rect 545240 5218 545324 5454
rect 545560 5218 548472 5454
rect -4476 5134 548472 5218
rect -4476 4898 -1564 5134
rect -1328 4898 -1244 5134
rect -1008 4898 4746 5134
rect 4982 4898 5066 5134
rect 5302 4898 22746 5134
rect 22982 4898 23066 5134
rect 23302 4898 40746 5134
rect 40982 4898 41066 5134
rect 41302 4898 58746 5134
rect 58982 4898 59066 5134
rect 59302 4898 76746 5134
rect 76982 4898 77066 5134
rect 77302 4898 94746 5134
rect 94982 4898 95066 5134
rect 95302 4898 112746 5134
rect 112982 4898 113066 5134
rect 113302 4898 130746 5134
rect 130982 4898 131066 5134
rect 131302 4898 148746 5134
rect 148982 4898 149066 5134
rect 149302 4898 166746 5134
rect 166982 4898 167066 5134
rect 167302 4898 184746 5134
rect 184982 4898 185066 5134
rect 185302 4898 202746 5134
rect 202982 4898 203066 5134
rect 203302 4898 220746 5134
rect 220982 4898 221066 5134
rect 221302 4898 238746 5134
rect 238982 4898 239066 5134
rect 239302 4898 256746 5134
rect 256982 4898 257066 5134
rect 257302 4898 274746 5134
rect 274982 4898 275066 5134
rect 275302 4898 292746 5134
rect 292982 4898 293066 5134
rect 293302 4898 310746 5134
rect 310982 4898 311066 5134
rect 311302 4898 328746 5134
rect 328982 4898 329066 5134
rect 329302 4898 346746 5134
rect 346982 4898 347066 5134
rect 347302 4898 364746 5134
rect 364982 4898 365066 5134
rect 365302 4898 382746 5134
rect 382982 4898 383066 5134
rect 383302 4898 400746 5134
rect 400982 4898 401066 5134
rect 401302 4898 418746 5134
rect 418982 4898 419066 5134
rect 419302 4898 436746 5134
rect 436982 4898 437066 5134
rect 437302 4898 454746 5134
rect 454982 4898 455066 5134
rect 455302 4898 472746 5134
rect 472982 4898 473066 5134
rect 473302 4898 490746 5134
rect 490982 4898 491066 5134
rect 491302 4898 508746 5134
rect 508982 4898 509066 5134
rect 509302 4898 526746 5134
rect 526982 4898 527066 5134
rect 527302 4898 545004 5134
rect 545240 4898 545324 5134
rect 545560 4898 548472 5134
rect -4476 4866 548472 4898
rect 100212 1138 108444 1180
rect 100212 902 100254 1138
rect 100490 902 108166 1138
rect 108402 902 108444 1138
rect 100212 860 108444 902
rect 108860 1138 137700 1180
rect 108860 902 108902 1138
rect 109138 902 137422 1138
rect 137658 902 137700 1138
rect 108860 860 137700 902
rect 137748 458 152052 500
rect 137748 222 137790 458
rect 138026 222 151774 458
rect 152010 222 152052 458
rect 137748 180 152052 222
rect -1596 -856 545592 -824
rect -1596 -1092 -1564 -856
rect -1328 -1092 -1244 -856
rect -1008 -1092 58746 -856
rect 58982 -1092 59066 -856
rect 59302 -1092 76746 -856
rect 76982 -1092 77066 -856
rect 77302 -1092 94746 -856
rect 94982 -1092 95066 -856
rect 95302 -1092 112746 -856
rect 112982 -1092 113066 -856
rect 113302 -1092 130746 -856
rect 130982 -1092 131066 -856
rect 131302 -1092 148746 -856
rect 148982 -1092 149066 -856
rect 149302 -1092 166746 -856
rect 166982 -1092 167066 -856
rect 167302 -1092 184746 -856
rect 184982 -1092 185066 -856
rect 185302 -1092 202746 -856
rect 202982 -1092 203066 -856
rect 203302 -1092 220746 -856
rect 220982 -1092 221066 -856
rect 221302 -1092 238746 -856
rect 238982 -1092 239066 -856
rect 239302 -1092 256746 -856
rect 256982 -1092 257066 -856
rect 257302 -1092 274746 -856
rect 274982 -1092 275066 -856
rect 275302 -1092 292746 -856
rect 292982 -1092 293066 -856
rect 293302 -1092 310746 -856
rect 310982 -1092 311066 -856
rect 311302 -1092 328746 -856
rect 328982 -1092 329066 -856
rect 329302 -1092 346746 -856
rect 346982 -1092 347066 -856
rect 347302 -1092 364746 -856
rect 364982 -1092 365066 -856
rect 365302 -1092 382746 -856
rect 382982 -1092 383066 -856
rect 383302 -1092 400746 -856
rect 400982 -1092 401066 -856
rect 401302 -1092 418746 -856
rect 418982 -1092 419066 -856
rect 419302 -1092 436746 -856
rect 436982 -1092 437066 -856
rect 437302 -1092 454746 -856
rect 454982 -1092 455066 -856
rect 455302 -1092 472746 -856
rect 472982 -1092 473066 -856
rect 473302 -1092 490746 -856
rect 490982 -1092 491066 -856
rect 491302 -1092 545004 -856
rect 545240 -1092 545324 -856
rect 545560 -1092 545592 -856
rect -1596 -1176 545592 -1092
rect -1596 -1412 -1564 -1176
rect -1328 -1412 -1244 -1176
rect -1008 -1412 58746 -1176
rect 58982 -1412 59066 -1176
rect 59302 -1412 76746 -1176
rect 76982 -1412 77066 -1176
rect 77302 -1412 94746 -1176
rect 94982 -1412 95066 -1176
rect 95302 -1412 112746 -1176
rect 112982 -1412 113066 -1176
rect 113302 -1412 130746 -1176
rect 130982 -1412 131066 -1176
rect 131302 -1412 148746 -1176
rect 148982 -1412 149066 -1176
rect 149302 -1412 166746 -1176
rect 166982 -1412 167066 -1176
rect 167302 -1412 184746 -1176
rect 184982 -1412 185066 -1176
rect 185302 -1412 202746 -1176
rect 202982 -1412 203066 -1176
rect 203302 -1412 220746 -1176
rect 220982 -1412 221066 -1176
rect 221302 -1412 238746 -1176
rect 238982 -1412 239066 -1176
rect 239302 -1412 256746 -1176
rect 256982 -1412 257066 -1176
rect 257302 -1412 274746 -1176
rect 274982 -1412 275066 -1176
rect 275302 -1412 292746 -1176
rect 292982 -1412 293066 -1176
rect 293302 -1412 310746 -1176
rect 310982 -1412 311066 -1176
rect 311302 -1412 328746 -1176
rect 328982 -1412 329066 -1176
rect 329302 -1412 346746 -1176
rect 346982 -1412 347066 -1176
rect 347302 -1412 364746 -1176
rect 364982 -1412 365066 -1176
rect 365302 -1412 382746 -1176
rect 382982 -1412 383066 -1176
rect 383302 -1412 400746 -1176
rect 400982 -1412 401066 -1176
rect 401302 -1412 418746 -1176
rect 418982 -1412 419066 -1176
rect 419302 -1412 436746 -1176
rect 436982 -1412 437066 -1176
rect 437302 -1412 454746 -1176
rect 454982 -1412 455066 -1176
rect 455302 -1412 472746 -1176
rect 472982 -1412 473066 -1176
rect 473302 -1412 490746 -1176
rect 490982 -1412 491066 -1176
rect 491302 -1412 545004 -1176
rect 545240 -1412 545324 -1176
rect 545560 -1412 545592 -1176
rect -1596 -1444 545592 -1412
rect -2556 -1816 546552 -1784
rect -2556 -2052 -2524 -1816
rect -2288 -2052 -2204 -1816
rect -1968 -2052 62466 -1816
rect 62702 -2052 62786 -1816
rect 63022 -2052 80466 -1816
rect 80702 -2052 80786 -1816
rect 81022 -2052 98466 -1816
rect 98702 -2052 98786 -1816
rect 99022 -2052 116466 -1816
rect 116702 -2052 116786 -1816
rect 117022 -2052 134466 -1816
rect 134702 -2052 134786 -1816
rect 135022 -2052 152466 -1816
rect 152702 -2052 152786 -1816
rect 153022 -2052 170466 -1816
rect 170702 -2052 170786 -1816
rect 171022 -2052 188466 -1816
rect 188702 -2052 188786 -1816
rect 189022 -2052 206466 -1816
rect 206702 -2052 206786 -1816
rect 207022 -2052 224466 -1816
rect 224702 -2052 224786 -1816
rect 225022 -2052 242466 -1816
rect 242702 -2052 242786 -1816
rect 243022 -2052 260466 -1816
rect 260702 -2052 260786 -1816
rect 261022 -2052 278466 -1816
rect 278702 -2052 278786 -1816
rect 279022 -2052 296466 -1816
rect 296702 -2052 296786 -1816
rect 297022 -2052 314466 -1816
rect 314702 -2052 314786 -1816
rect 315022 -2052 332466 -1816
rect 332702 -2052 332786 -1816
rect 333022 -2052 350466 -1816
rect 350702 -2052 350786 -1816
rect 351022 -2052 368466 -1816
rect 368702 -2052 368786 -1816
rect 369022 -2052 386466 -1816
rect 386702 -2052 386786 -1816
rect 387022 -2052 404466 -1816
rect 404702 -2052 404786 -1816
rect 405022 -2052 422466 -1816
rect 422702 -2052 422786 -1816
rect 423022 -2052 440466 -1816
rect 440702 -2052 440786 -1816
rect 441022 -2052 458466 -1816
rect 458702 -2052 458786 -1816
rect 459022 -2052 476466 -1816
rect 476702 -2052 476786 -1816
rect 477022 -2052 494466 -1816
rect 494702 -2052 494786 -1816
rect 495022 -2052 545964 -1816
rect 546200 -2052 546284 -1816
rect 546520 -2052 546552 -1816
rect -2556 -2136 546552 -2052
rect -2556 -2372 -2524 -2136
rect -2288 -2372 -2204 -2136
rect -1968 -2372 62466 -2136
rect 62702 -2372 62786 -2136
rect 63022 -2372 80466 -2136
rect 80702 -2372 80786 -2136
rect 81022 -2372 98466 -2136
rect 98702 -2372 98786 -2136
rect 99022 -2372 116466 -2136
rect 116702 -2372 116786 -2136
rect 117022 -2372 134466 -2136
rect 134702 -2372 134786 -2136
rect 135022 -2372 152466 -2136
rect 152702 -2372 152786 -2136
rect 153022 -2372 170466 -2136
rect 170702 -2372 170786 -2136
rect 171022 -2372 188466 -2136
rect 188702 -2372 188786 -2136
rect 189022 -2372 206466 -2136
rect 206702 -2372 206786 -2136
rect 207022 -2372 224466 -2136
rect 224702 -2372 224786 -2136
rect 225022 -2372 242466 -2136
rect 242702 -2372 242786 -2136
rect 243022 -2372 260466 -2136
rect 260702 -2372 260786 -2136
rect 261022 -2372 278466 -2136
rect 278702 -2372 278786 -2136
rect 279022 -2372 296466 -2136
rect 296702 -2372 296786 -2136
rect 297022 -2372 314466 -2136
rect 314702 -2372 314786 -2136
rect 315022 -2372 332466 -2136
rect 332702 -2372 332786 -2136
rect 333022 -2372 350466 -2136
rect 350702 -2372 350786 -2136
rect 351022 -2372 368466 -2136
rect 368702 -2372 368786 -2136
rect 369022 -2372 386466 -2136
rect 386702 -2372 386786 -2136
rect 387022 -2372 404466 -2136
rect 404702 -2372 404786 -2136
rect 405022 -2372 422466 -2136
rect 422702 -2372 422786 -2136
rect 423022 -2372 440466 -2136
rect 440702 -2372 440786 -2136
rect 441022 -2372 458466 -2136
rect 458702 -2372 458786 -2136
rect 459022 -2372 476466 -2136
rect 476702 -2372 476786 -2136
rect 477022 -2372 494466 -2136
rect 494702 -2372 494786 -2136
rect 495022 -2372 545964 -2136
rect 546200 -2372 546284 -2136
rect 546520 -2372 546552 -2136
rect -2556 -2404 546552 -2372
rect -3516 -2776 547512 -2744
rect -3516 -3012 -3484 -2776
rect -3248 -3012 -3164 -2776
rect -2928 -3012 48186 -2776
rect 48422 -3012 48506 -2776
rect 48742 -3012 66186 -2776
rect 66422 -3012 66506 -2776
rect 66742 -3012 84186 -2776
rect 84422 -3012 84506 -2776
rect 84742 -3012 102186 -2776
rect 102422 -3012 102506 -2776
rect 102742 -3012 120186 -2776
rect 120422 -3012 120506 -2776
rect 120742 -3012 138186 -2776
rect 138422 -3012 138506 -2776
rect 138742 -3012 156186 -2776
rect 156422 -3012 156506 -2776
rect 156742 -3012 174186 -2776
rect 174422 -3012 174506 -2776
rect 174742 -3012 192186 -2776
rect 192422 -3012 192506 -2776
rect 192742 -3012 210186 -2776
rect 210422 -3012 210506 -2776
rect 210742 -3012 228186 -2776
rect 228422 -3012 228506 -2776
rect 228742 -3012 246186 -2776
rect 246422 -3012 246506 -2776
rect 246742 -3012 264186 -2776
rect 264422 -3012 264506 -2776
rect 264742 -3012 282186 -2776
rect 282422 -3012 282506 -2776
rect 282742 -3012 300186 -2776
rect 300422 -3012 300506 -2776
rect 300742 -3012 318186 -2776
rect 318422 -3012 318506 -2776
rect 318742 -3012 336186 -2776
rect 336422 -3012 336506 -2776
rect 336742 -3012 354186 -2776
rect 354422 -3012 354506 -2776
rect 354742 -3012 372186 -2776
rect 372422 -3012 372506 -2776
rect 372742 -3012 390186 -2776
rect 390422 -3012 390506 -2776
rect 390742 -3012 408186 -2776
rect 408422 -3012 408506 -2776
rect 408742 -3012 426186 -2776
rect 426422 -3012 426506 -2776
rect 426742 -3012 444186 -2776
rect 444422 -3012 444506 -2776
rect 444742 -3012 462186 -2776
rect 462422 -3012 462506 -2776
rect 462742 -3012 480186 -2776
rect 480422 -3012 480506 -2776
rect 480742 -3012 498186 -2776
rect 498422 -3012 498506 -2776
rect 498742 -3012 546924 -2776
rect 547160 -3012 547244 -2776
rect 547480 -3012 547512 -2776
rect -3516 -3096 547512 -3012
rect -3516 -3332 -3484 -3096
rect -3248 -3332 -3164 -3096
rect -2928 -3332 48186 -3096
rect 48422 -3332 48506 -3096
rect 48742 -3332 66186 -3096
rect 66422 -3332 66506 -3096
rect 66742 -3332 84186 -3096
rect 84422 -3332 84506 -3096
rect 84742 -3332 102186 -3096
rect 102422 -3332 102506 -3096
rect 102742 -3332 120186 -3096
rect 120422 -3332 120506 -3096
rect 120742 -3332 138186 -3096
rect 138422 -3332 138506 -3096
rect 138742 -3332 156186 -3096
rect 156422 -3332 156506 -3096
rect 156742 -3332 174186 -3096
rect 174422 -3332 174506 -3096
rect 174742 -3332 192186 -3096
rect 192422 -3332 192506 -3096
rect 192742 -3332 210186 -3096
rect 210422 -3332 210506 -3096
rect 210742 -3332 228186 -3096
rect 228422 -3332 228506 -3096
rect 228742 -3332 246186 -3096
rect 246422 -3332 246506 -3096
rect 246742 -3332 264186 -3096
rect 264422 -3332 264506 -3096
rect 264742 -3332 282186 -3096
rect 282422 -3332 282506 -3096
rect 282742 -3332 300186 -3096
rect 300422 -3332 300506 -3096
rect 300742 -3332 318186 -3096
rect 318422 -3332 318506 -3096
rect 318742 -3332 336186 -3096
rect 336422 -3332 336506 -3096
rect 336742 -3332 354186 -3096
rect 354422 -3332 354506 -3096
rect 354742 -3332 372186 -3096
rect 372422 -3332 372506 -3096
rect 372742 -3332 390186 -3096
rect 390422 -3332 390506 -3096
rect 390742 -3332 408186 -3096
rect 408422 -3332 408506 -3096
rect 408742 -3332 426186 -3096
rect 426422 -3332 426506 -3096
rect 426742 -3332 444186 -3096
rect 444422 -3332 444506 -3096
rect 444742 -3332 462186 -3096
rect 462422 -3332 462506 -3096
rect 462742 -3332 480186 -3096
rect 480422 -3332 480506 -3096
rect 480742 -3332 498186 -3096
rect 498422 -3332 498506 -3096
rect 498742 -3332 546924 -3096
rect 547160 -3332 547244 -3096
rect 547480 -3332 547512 -3096
rect -3516 -3364 547512 -3332
rect -4476 -3736 548472 -3704
rect -4476 -3972 -4444 -3736
rect -4208 -3972 -4124 -3736
rect -3888 -3972 51906 -3736
rect 52142 -3972 52226 -3736
rect 52462 -3972 69906 -3736
rect 70142 -3972 70226 -3736
rect 70462 -3972 87906 -3736
rect 88142 -3972 88226 -3736
rect 88462 -3972 105906 -3736
rect 106142 -3972 106226 -3736
rect 106462 -3972 123906 -3736
rect 124142 -3972 124226 -3736
rect 124462 -3972 141906 -3736
rect 142142 -3972 142226 -3736
rect 142462 -3972 159906 -3736
rect 160142 -3972 160226 -3736
rect 160462 -3972 177906 -3736
rect 178142 -3972 178226 -3736
rect 178462 -3972 195906 -3736
rect 196142 -3972 196226 -3736
rect 196462 -3972 213906 -3736
rect 214142 -3972 214226 -3736
rect 214462 -3972 231906 -3736
rect 232142 -3972 232226 -3736
rect 232462 -3972 249906 -3736
rect 250142 -3972 250226 -3736
rect 250462 -3972 267906 -3736
rect 268142 -3972 268226 -3736
rect 268462 -3972 285906 -3736
rect 286142 -3972 286226 -3736
rect 286462 -3972 303906 -3736
rect 304142 -3972 304226 -3736
rect 304462 -3972 321906 -3736
rect 322142 -3972 322226 -3736
rect 322462 -3972 339906 -3736
rect 340142 -3972 340226 -3736
rect 340462 -3972 357906 -3736
rect 358142 -3972 358226 -3736
rect 358462 -3972 375906 -3736
rect 376142 -3972 376226 -3736
rect 376462 -3972 393906 -3736
rect 394142 -3972 394226 -3736
rect 394462 -3972 411906 -3736
rect 412142 -3972 412226 -3736
rect 412462 -3972 429906 -3736
rect 430142 -3972 430226 -3736
rect 430462 -3972 447906 -3736
rect 448142 -3972 448226 -3736
rect 448462 -3972 465906 -3736
rect 466142 -3972 466226 -3736
rect 466462 -3972 483906 -3736
rect 484142 -3972 484226 -3736
rect 484462 -3972 547884 -3736
rect 548120 -3972 548204 -3736
rect 548440 -3972 548472 -3736
rect -4476 -4056 548472 -3972
rect -4476 -4292 -4444 -4056
rect -4208 -4292 -4124 -4056
rect -3888 -4292 51906 -4056
rect 52142 -4292 52226 -4056
rect 52462 -4292 69906 -4056
rect 70142 -4292 70226 -4056
rect 70462 -4292 87906 -4056
rect 88142 -4292 88226 -4056
rect 88462 -4292 105906 -4056
rect 106142 -4292 106226 -4056
rect 106462 -4292 123906 -4056
rect 124142 -4292 124226 -4056
rect 124462 -4292 141906 -4056
rect 142142 -4292 142226 -4056
rect 142462 -4292 159906 -4056
rect 160142 -4292 160226 -4056
rect 160462 -4292 177906 -4056
rect 178142 -4292 178226 -4056
rect 178462 -4292 195906 -4056
rect 196142 -4292 196226 -4056
rect 196462 -4292 213906 -4056
rect 214142 -4292 214226 -4056
rect 214462 -4292 231906 -4056
rect 232142 -4292 232226 -4056
rect 232462 -4292 249906 -4056
rect 250142 -4292 250226 -4056
rect 250462 -4292 267906 -4056
rect 268142 -4292 268226 -4056
rect 268462 -4292 285906 -4056
rect 286142 -4292 286226 -4056
rect 286462 -4292 303906 -4056
rect 304142 -4292 304226 -4056
rect 304462 -4292 321906 -4056
rect 322142 -4292 322226 -4056
rect 322462 -4292 339906 -4056
rect 340142 -4292 340226 -4056
rect 340462 -4292 357906 -4056
rect 358142 -4292 358226 -4056
rect 358462 -4292 375906 -4056
rect 376142 -4292 376226 -4056
rect 376462 -4292 393906 -4056
rect 394142 -4292 394226 -4056
rect 394462 -4292 411906 -4056
rect 412142 -4292 412226 -4056
rect 412462 -4292 429906 -4056
rect 430142 -4292 430226 -4056
rect 430462 -4292 447906 -4056
rect 448142 -4292 448226 -4056
rect 448462 -4292 465906 -4056
rect 466142 -4292 466226 -4056
rect 466462 -4292 483906 -4056
rect 484142 -4292 484226 -4056
rect 484462 -4292 547884 -4056
rect 548120 -4292 548204 -4056
rect 548440 -4292 548472 -4056
rect -4476 -4324 548472 -4292
use ahb_counter  frigate_prj
timestamp 0
transform 1 0 90000 0 1 20000
box 0 0 1 1
<< labels >>
flabel metal2 s 51622 -400 51678 800 0 FreeSans 224 90 0 0 HADDR[0]
port 0 nsew signal input
flabel metal2 s 67262 -400 67318 800 0 FreeSans 224 90 0 0 HADDR[10]
port 1 nsew signal input
flabel metal2 s 68826 -400 68882 800 0 FreeSans 224 90 0 0 HADDR[11]
port 2 nsew signal input
flabel metal2 s 70390 -400 70446 800 0 FreeSans 224 90 0 0 HADDR[12]
port 3 nsew signal input
flabel metal2 s 71954 -400 72010 800 0 FreeSans 224 90 0 0 HADDR[13]
port 4 nsew signal input
flabel metal2 s 73518 -400 73574 800 0 FreeSans 224 90 0 0 HADDR[14]
port 5 nsew signal input
flabel metal2 s 75082 -400 75138 800 0 FreeSans 224 90 0 0 HADDR[15]
port 6 nsew signal input
flabel metal2 s 76646 -400 76702 800 0 FreeSans 224 90 0 0 HADDR[16]
port 7 nsew signal input
flabel metal2 s 78210 -400 78266 800 0 FreeSans 224 90 0 0 HADDR[17]
port 8 nsew signal input
flabel metal2 s 79774 -400 79830 800 0 FreeSans 224 90 0 0 HADDR[18]
port 9 nsew signal input
flabel metal2 s 81338 -400 81394 800 0 FreeSans 224 90 0 0 HADDR[19]
port 10 nsew signal input
flabel metal2 s 53186 -400 53242 800 0 FreeSans 224 90 0 0 HADDR[1]
port 11 nsew signal input
flabel metal2 s 82902 -400 82958 800 0 FreeSans 224 90 0 0 HADDR[20]
port 12 nsew signal input
flabel metal2 s 84466 -400 84522 800 0 FreeSans 224 90 0 0 HADDR[21]
port 13 nsew signal input
flabel metal2 s 86030 -400 86086 800 0 FreeSans 224 90 0 0 HADDR[22]
port 14 nsew signal input
flabel metal2 s 87594 -400 87650 800 0 FreeSans 224 90 0 0 HADDR[23]
port 15 nsew signal input
flabel metal2 s 89158 -400 89214 800 0 FreeSans 224 90 0 0 HADDR[24]
port 16 nsew signal input
flabel metal2 s 90722 -400 90778 800 0 FreeSans 224 90 0 0 HADDR[25]
port 17 nsew signal input
flabel metal2 s 92286 -400 92342 800 0 FreeSans 224 90 0 0 HADDR[26]
port 18 nsew signal input
flabel metal2 s 93850 -400 93906 800 0 FreeSans 224 90 0 0 HADDR[27]
port 19 nsew signal input
flabel metal2 s 95414 -400 95470 800 0 FreeSans 224 90 0 0 HADDR[28]
port 20 nsew signal input
flabel metal2 s 96978 -400 97034 800 0 FreeSans 224 90 0 0 HADDR[29]
port 21 nsew signal input
flabel metal2 s 54750 -400 54806 800 0 FreeSans 224 90 0 0 HADDR[2]
port 22 nsew signal input
flabel metal2 s 98542 -400 98598 800 0 FreeSans 224 90 0 0 HADDR[30]
port 23 nsew signal input
flabel metal2 s 100106 -400 100162 800 0 FreeSans 224 90 0 0 HADDR[31]
port 24 nsew signal input
flabel metal2 s 56314 -400 56370 800 0 FreeSans 224 90 0 0 HADDR[3]
port 25 nsew signal input
flabel metal2 s 57878 -400 57934 800 0 FreeSans 224 90 0 0 HADDR[4]
port 26 nsew signal input
flabel metal2 s 59442 -400 59498 800 0 FreeSans 224 90 0 0 HADDR[5]
port 27 nsew signal input
flabel metal2 s 61006 -400 61062 800 0 FreeSans 224 90 0 0 HADDR[6]
port 28 nsew signal input
flabel metal2 s 62570 -400 62626 800 0 FreeSans 224 90 0 0 HADDR[7]
port 29 nsew signal input
flabel metal2 s 64134 -400 64190 800 0 FreeSans 224 90 0 0 HADDR[8]
port 30 nsew signal input
flabel metal2 s 65698 -400 65754 800 0 FreeSans 224 90 0 0 HADDR[9]
port 31 nsew signal input
flabel metal2 s 46930 -400 46986 800 0 FreeSans 224 90 0 0 HCLK
port 32 nsew signal input
flabel metal2 s 162666 -400 162722 800 0 FreeSans 224 90 0 0 HRDATA[0]
port 33 nsew signal output
flabel metal2 s 178306 -400 178362 800 0 FreeSans 224 90 0 0 HRDATA[10]
port 34 nsew signal output
flabel metal2 s 179870 -400 179926 800 0 FreeSans 224 90 0 0 HRDATA[11]
port 35 nsew signal output
flabel metal2 s 181434 -400 181490 800 0 FreeSans 224 90 0 0 HRDATA[12]
port 36 nsew signal output
flabel metal2 s 182998 -400 183054 800 0 FreeSans 224 90 0 0 HRDATA[13]
port 37 nsew signal output
flabel metal2 s 184562 -400 184618 800 0 FreeSans 224 90 0 0 HRDATA[14]
port 38 nsew signal output
flabel metal2 s 186126 -400 186182 800 0 FreeSans 224 90 0 0 HRDATA[15]
port 39 nsew signal output
flabel metal2 s 187690 -400 187746 800 0 FreeSans 224 90 0 0 HRDATA[16]
port 40 nsew signal output
flabel metal2 s 189254 -400 189310 800 0 FreeSans 224 90 0 0 HRDATA[17]
port 41 nsew signal output
flabel metal2 s 190818 -400 190874 800 0 FreeSans 224 90 0 0 HRDATA[18]
port 42 nsew signal output
flabel metal2 s 192382 -400 192438 800 0 FreeSans 224 90 0 0 HRDATA[19]
port 43 nsew signal output
flabel metal2 s 164230 -400 164286 800 0 FreeSans 224 90 0 0 HRDATA[1]
port 44 nsew signal output
flabel metal2 s 193946 -400 194002 800 0 FreeSans 224 90 0 0 HRDATA[20]
port 45 nsew signal output
flabel metal2 s 195510 -400 195566 800 0 FreeSans 224 90 0 0 HRDATA[21]
port 46 nsew signal output
flabel metal2 s 197074 -400 197130 800 0 FreeSans 224 90 0 0 HRDATA[22]
port 47 nsew signal output
flabel metal2 s 198638 -400 198694 800 0 FreeSans 224 90 0 0 HRDATA[23]
port 48 nsew signal output
flabel metal2 s 200202 -400 200258 800 0 FreeSans 224 90 0 0 HRDATA[24]
port 49 nsew signal output
flabel metal2 s 201766 -400 201822 800 0 FreeSans 224 90 0 0 HRDATA[25]
port 50 nsew signal output
flabel metal2 s 203330 -400 203386 800 0 FreeSans 224 90 0 0 HRDATA[26]
port 51 nsew signal output
flabel metal2 s 204894 -400 204950 800 0 FreeSans 224 90 0 0 HRDATA[27]
port 52 nsew signal output
flabel metal2 s 206458 -400 206514 800 0 FreeSans 224 90 0 0 HRDATA[28]
port 53 nsew signal output
flabel metal2 s 208022 -400 208078 800 0 FreeSans 224 90 0 0 HRDATA[29]
port 54 nsew signal output
flabel metal2 s 165794 -400 165850 800 0 FreeSans 224 90 0 0 HRDATA[2]
port 55 nsew signal output
flabel metal2 s 209586 -400 209642 800 0 FreeSans 224 90 0 0 HRDATA[30]
port 56 nsew signal output
flabel metal2 s 211150 -400 211206 800 0 FreeSans 224 90 0 0 HRDATA[31]
port 57 nsew signal output
flabel metal2 s 167358 -400 167414 800 0 FreeSans 224 90 0 0 HRDATA[3]
port 58 nsew signal output
flabel metal2 s 168922 -400 168978 800 0 FreeSans 224 90 0 0 HRDATA[4]
port 59 nsew signal output
flabel metal2 s 170486 -400 170542 800 0 FreeSans 224 90 0 0 HRDATA[5]
port 60 nsew signal output
flabel metal2 s 172050 -400 172106 800 0 FreeSans 224 90 0 0 HRDATA[6]
port 61 nsew signal output
flabel metal2 s 173614 -400 173670 800 0 FreeSans 224 90 0 0 HRDATA[7]
port 62 nsew signal output
flabel metal2 s 175178 -400 175234 800 0 FreeSans 224 90 0 0 HRDATA[8]
port 63 nsew signal output
flabel metal2 s 176742 -400 176798 800 0 FreeSans 224 90 0 0 HRDATA[9]
port 64 nsew signal output
flabel metal2 s 151718 -400 151774 800 0 FreeSans 224 90 0 0 HREADY
port 65 nsew signal input
flabel metal2 s 212714 -400 212770 800 0 FreeSans 224 90 0 0 HREADYOUT
port 66 nsew signal output
flabel metal2 s 48494 -400 48550 800 0 FreeSans 224 90 0 0 HRESETn
port 67 nsew signal input
flabel metal2 s 50058 -400 50114 800 0 FreeSans 224 90 0 0 HSEL
port 68 nsew signal input
flabel metal2 s 157974 -400 158030 800 0 FreeSans 224 90 0 0 HSIZE[0]
port 69 nsew signal input
flabel metal2 s 159538 -400 159594 800 0 FreeSans 224 90 0 0 HSIZE[1]
port 70 nsew signal input
flabel metal2 s 161102 -400 161158 800 0 FreeSans 224 90 0 0 HSIZE[2]
port 71 nsew signal input
flabel metal2 s 154846 -400 154902 800 0 FreeSans 224 90 0 0 HTRANS[0]
port 72 nsew signal input
flabel metal2 s 156410 -400 156466 800 0 FreeSans 224 90 0 0 HTRANS[1]
port 73 nsew signal input
flabel metal2 s 101670 -400 101726 800 0 FreeSans 224 90 0 0 HWDATA[0]
port 74 nsew signal input
flabel metal2 s 117310 -400 117366 800 0 FreeSans 224 90 0 0 HWDATA[10]
port 75 nsew signal input
flabel metal2 s 118874 -400 118930 800 0 FreeSans 224 90 0 0 HWDATA[11]
port 76 nsew signal input
flabel metal2 s 120438 -400 120494 800 0 FreeSans 224 90 0 0 HWDATA[12]
port 77 nsew signal input
flabel metal2 s 122002 -400 122058 800 0 FreeSans 224 90 0 0 HWDATA[13]
port 78 nsew signal input
flabel metal2 s 123566 -400 123622 800 0 FreeSans 224 90 0 0 HWDATA[14]
port 79 nsew signal input
flabel metal2 s 125130 -400 125186 800 0 FreeSans 224 90 0 0 HWDATA[15]
port 80 nsew signal input
flabel metal2 s 126694 -400 126750 800 0 FreeSans 224 90 0 0 HWDATA[16]
port 81 nsew signal input
flabel metal2 s 128258 -400 128314 800 0 FreeSans 224 90 0 0 HWDATA[17]
port 82 nsew signal input
flabel metal2 s 129822 -400 129878 800 0 FreeSans 224 90 0 0 HWDATA[18]
port 83 nsew signal input
flabel metal2 s 131386 -400 131442 800 0 FreeSans 224 90 0 0 HWDATA[19]
port 84 nsew signal input
flabel metal2 s 103234 -400 103290 800 0 FreeSans 224 90 0 0 HWDATA[1]
port 85 nsew signal input
flabel metal2 s 132950 -400 133006 800 0 FreeSans 224 90 0 0 HWDATA[20]
port 86 nsew signal input
flabel metal2 s 134514 -400 134570 800 0 FreeSans 224 90 0 0 HWDATA[21]
port 87 nsew signal input
flabel metal2 s 136078 -400 136134 800 0 FreeSans 224 90 0 0 HWDATA[22]
port 88 nsew signal input
flabel metal2 s 137642 -400 137698 800 0 FreeSans 224 90 0 0 HWDATA[23]
port 89 nsew signal input
flabel metal2 s 139206 -400 139262 800 0 FreeSans 224 90 0 0 HWDATA[24]
port 90 nsew signal input
flabel metal2 s 140770 -400 140826 800 0 FreeSans 224 90 0 0 HWDATA[25]
port 91 nsew signal input
flabel metal2 s 142334 -400 142390 800 0 FreeSans 224 90 0 0 HWDATA[26]
port 92 nsew signal input
flabel metal2 s 143898 -400 143954 800 0 FreeSans 224 90 0 0 HWDATA[27]
port 93 nsew signal input
flabel metal2 s 145462 -400 145518 800 0 FreeSans 224 90 0 0 HWDATA[28]
port 94 nsew signal input
flabel metal2 s 147026 -400 147082 800 0 FreeSans 224 90 0 0 HWDATA[29]
port 95 nsew signal input
flabel metal2 s 104798 -400 104854 800 0 FreeSans 224 90 0 0 HWDATA[2]
port 96 nsew signal input
flabel metal2 s 148590 -400 148646 800 0 FreeSans 224 90 0 0 HWDATA[30]
port 97 nsew signal input
flabel metal2 s 150154 -400 150210 800 0 FreeSans 224 90 0 0 HWDATA[31]
port 98 nsew signal input
flabel metal2 s 106362 -400 106418 800 0 FreeSans 224 90 0 0 HWDATA[3]
port 99 nsew signal input
flabel metal2 s 107926 -400 107982 800 0 FreeSans 224 90 0 0 HWDATA[4]
port 100 nsew signal input
flabel metal2 s 109490 -400 109546 800 0 FreeSans 224 90 0 0 HWDATA[5]
port 101 nsew signal input
flabel metal2 s 111054 -400 111110 800 0 FreeSans 224 90 0 0 HWDATA[6]
port 102 nsew signal input
flabel metal2 s 112618 -400 112674 800 0 FreeSans 224 90 0 0 HWDATA[7]
port 103 nsew signal input
flabel metal2 s 114182 -400 114238 800 0 FreeSans 224 90 0 0 HWDATA[8]
port 104 nsew signal input
flabel metal2 s 115746 -400 115802 800 0 FreeSans 224 90 0 0 HWDATA[9]
port 105 nsew signal input
flabel metal2 s 153282 -400 153338 800 0 FreeSans 224 90 0 0 HWRITE
port 106 nsew signal input
flabel metal4 s 339625 459700 339753 460000 0 FreeSans 960 90 0 0 adc0
port 107 nsew signal bidirectional
flabel metal4 s 340137 459700 340265 460000 0 FreeSans 960 90 0 0 adc1
port 108 nsew signal bidirectional
flabel metal4 s 340649 459700 340777 460000 0 FreeSans 960 90 0 0 comp_n
port 109 nsew signal bidirectional
flabel metal4 s 341161 459700 341289 460000 0 FreeSans 960 90 0 0 comp_p
port 110 nsew signal bidirectional
flabel metal4 s 336553 459700 336681 460000 0 FreeSans 960 90 0 0 dac0
port 111 nsew signal bidirectional
flabel metal4 s 337065 459700 337193 460000 0 FreeSans 960 90 0 0 dac1
port 112 nsew signal bidirectional
flabel metal3 s 543200 19418 544400 19538 0 FreeSans 480 0 0 0 gpio0_in[0]
port 113 nsew signal input
flabel metal3 s 543200 33290 544400 33410 0 FreeSans 480 0 0 0 gpio0_in[1]
port 114 nsew signal input
flabel metal3 s 543200 47162 544400 47282 0 FreeSans 480 0 0 0 gpio0_in[2]
port 115 nsew signal input
flabel metal3 s 543200 61034 544400 61154 0 FreeSans 480 0 0 0 gpio0_in[3]
port 116 nsew signal input
flabel metal3 s 543200 74906 544400 75026 0 FreeSans 480 0 0 0 gpio0_in[4]
port 117 nsew signal input
flabel metal3 s 543200 88778 544400 88898 0 FreeSans 480 0 0 0 gpio0_in[5]
port 118 nsew signal input
flabel metal3 s 543200 102650 544400 102770 0 FreeSans 480 0 0 0 gpio0_in[6]
port 119 nsew signal input
flabel metal3 s 543200 116522 544400 116642 0 FreeSans 480 0 0 0 gpio0_in[7]
port 120 nsew signal input
flabel metal3 s 543200 28666 544400 28786 0 FreeSans 480 0 0 0 gpio0_oeb[0]
port 121 nsew signal output
flabel metal3 s 543200 42538 544400 42658 0 FreeSans 480 0 0 0 gpio0_oeb[1]
port 122 nsew signal output
flabel metal3 s 543200 56410 544400 56530 0 FreeSans 480 0 0 0 gpio0_oeb[2]
port 123 nsew signal output
flabel metal3 s 543200 70282 544400 70402 0 FreeSans 480 0 0 0 gpio0_oeb[3]
port 124 nsew signal output
flabel metal3 s 543200 84154 544400 84274 0 FreeSans 480 0 0 0 gpio0_oeb[4]
port 125 nsew signal output
flabel metal3 s 543200 98026 544400 98146 0 FreeSans 480 0 0 0 gpio0_oeb[5]
port 126 nsew signal output
flabel metal3 s 543200 111898 544400 112018 0 FreeSans 480 0 0 0 gpio0_oeb[6]
port 127 nsew signal output
flabel metal3 s 543200 125770 544400 125890 0 FreeSans 480 0 0 0 gpio0_oeb[7]
port 128 nsew signal output
flabel metal3 s 543200 24042 544400 24162 0 FreeSans 480 0 0 0 gpio0_out[0]
port 129 nsew signal output
flabel metal3 s 543200 37914 544400 38034 0 FreeSans 480 0 0 0 gpio0_out[1]
port 130 nsew signal output
flabel metal3 s 543200 51786 544400 51906 0 FreeSans 480 0 0 0 gpio0_out[2]
port 131 nsew signal output
flabel metal3 s 543200 65658 544400 65778 0 FreeSans 480 0 0 0 gpio0_out[3]
port 132 nsew signal output
flabel metal3 s 543200 79530 544400 79650 0 FreeSans 480 0 0 0 gpio0_out[4]
port 133 nsew signal output
flabel metal3 s 543200 93402 544400 93522 0 FreeSans 480 0 0 0 gpio0_out[5]
port 134 nsew signal output
flabel metal3 s 543200 107274 544400 107394 0 FreeSans 480 0 0 0 gpio0_out[6]
port 135 nsew signal output
flabel metal3 s 543200 121146 544400 121266 0 FreeSans 480 0 0 0 gpio0_out[7]
port 136 nsew signal output
flabel metal3 s 543200 178984 544400 179104 0 FreeSans 480 0 0 0 gpio1_in[0]
port 137 nsew signal input
flabel metal3 s 543200 192856 544400 192976 0 FreeSans 480 0 0 0 gpio1_in[1]
port 138 nsew signal input
flabel metal3 s 543200 206728 544400 206848 0 FreeSans 480 0 0 0 gpio1_in[2]
port 139 nsew signal input
flabel metal3 s 543200 220600 544400 220720 0 FreeSans 480 0 0 0 gpio1_in[3]
port 140 nsew signal input
flabel metal3 s 543200 234472 544400 234592 0 FreeSans 480 0 0 0 gpio1_in[4]
port 141 nsew signal input
flabel metal3 s 543200 248344 544400 248464 0 FreeSans 480 0 0 0 gpio1_in[5]
port 142 nsew signal input
flabel metal3 s 543200 262216 544400 262336 0 FreeSans 480 0 0 0 gpio1_in[6]
port 143 nsew signal input
flabel metal3 s 543200 276088 544400 276208 0 FreeSans 480 0 0 0 gpio1_in[7]
port 144 nsew signal input
flabel metal3 s 543200 188232 544400 188352 0 FreeSans 480 0 0 0 gpio1_oeb[0]
port 145 nsew signal output
flabel metal3 s 543200 202104 544400 202224 0 FreeSans 480 0 0 0 gpio1_oeb[1]
port 146 nsew signal output
flabel metal3 s 543200 215976 544400 216096 0 FreeSans 480 0 0 0 gpio1_oeb[2]
port 147 nsew signal output
flabel metal3 s 543200 229848 544400 229968 0 FreeSans 480 0 0 0 gpio1_oeb[3]
port 148 nsew signal output
flabel metal3 s 543200 243720 544400 243840 0 FreeSans 480 0 0 0 gpio1_oeb[4]
port 149 nsew signal output
flabel metal3 s 543200 257592 544400 257712 0 FreeSans 480 0 0 0 gpio1_oeb[5]
port 150 nsew signal output
flabel metal3 s 543200 271464 544400 271584 0 FreeSans 480 0 0 0 gpio1_oeb[6]
port 151 nsew signal output
flabel metal3 s 543200 285336 544400 285456 0 FreeSans 480 0 0 0 gpio1_oeb[7]
port 152 nsew signal output
flabel metal3 s 543200 183608 544400 183728 0 FreeSans 480 0 0 0 gpio1_out[0]
port 153 nsew signal output
flabel metal3 s 543200 197480 544400 197600 0 FreeSans 480 0 0 0 gpio1_out[1]
port 154 nsew signal output
flabel metal3 s 543200 211352 544400 211472 0 FreeSans 480 0 0 0 gpio1_out[2]
port 155 nsew signal output
flabel metal3 s 543200 225224 544400 225344 0 FreeSans 480 0 0 0 gpio1_out[3]
port 156 nsew signal output
flabel metal3 s 543200 239096 544400 239216 0 FreeSans 480 0 0 0 gpio1_out[4]
port 157 nsew signal output
flabel metal3 s 543200 252968 544400 253088 0 FreeSans 480 0 0 0 gpio1_out[5]
port 158 nsew signal output
flabel metal3 s 543200 266840 544400 266960 0 FreeSans 480 0 0 0 gpio1_out[6]
port 159 nsew signal output
flabel metal3 s 543200 280712 544400 280832 0 FreeSans 480 0 0 0 gpio1_out[7]
port 160 nsew signal output
flabel metal3 s 543200 289960 544400 290080 0 FreeSans 480 0 0 0 gpio2_in[0]
port 161 nsew signal input
flabel metal3 s 543200 303832 544400 303952 0 FreeSans 480 0 0 0 gpio2_in[1]
port 162 nsew signal input
flabel metal3 s 543200 317704 544400 317824 0 FreeSans 480 0 0 0 gpio2_in[2]
port 163 nsew signal input
flabel metal3 s 543200 331576 544400 331696 0 FreeSans 480 0 0 0 gpio2_in[3]
port 164 nsew signal input
flabel metal3 s 543200 405560 544400 405680 0 FreeSans 480 0 0 0 gpio2_in[4]
port 165 nsew signal input
flabel metal3 s 543200 419432 544400 419552 0 FreeSans 480 0 0 0 gpio2_in[5]
port 166 nsew signal input
flabel metal3 s 543200 433304 544400 433424 0 FreeSans 480 0 0 0 gpio2_in[6]
port 167 nsew signal input
flabel metal3 s 543200 447176 544400 447296 0 FreeSans 480 0 0 0 gpio2_in[7]
port 168 nsew signal input
flabel metal3 s 543200 299208 544400 299328 0 FreeSans 480 0 0 0 gpio2_oeb[0]
port 169 nsew signal output
flabel metal3 s 543200 313080 544400 313200 0 FreeSans 480 0 0 0 gpio2_oeb[1]
port 170 nsew signal output
flabel metal3 s 543200 326952 544400 327072 0 FreeSans 480 0 0 0 gpio2_oeb[2]
port 171 nsew signal output
flabel metal3 s 543200 340824 544400 340944 0 FreeSans 480 0 0 0 gpio2_oeb[3]
port 172 nsew signal output
flabel metal3 s 543200 414808 544400 414928 0 FreeSans 480 0 0 0 gpio2_oeb[4]
port 173 nsew signal output
flabel metal3 s 543200 428680 544400 428800 0 FreeSans 480 0 0 0 gpio2_oeb[5]
port 174 nsew signal output
flabel metal3 s 543200 442552 544400 442672 0 FreeSans 480 0 0 0 gpio2_oeb[6]
port 175 nsew signal output
flabel metal3 s 543200 456424 544400 456544 0 FreeSans 480 0 0 0 gpio2_oeb[7]
port 176 nsew signal output
flabel metal3 s 543200 294584 544400 294704 0 FreeSans 480 0 0 0 gpio2_out[0]
port 177 nsew signal output
flabel metal3 s 543200 308456 544400 308576 0 FreeSans 480 0 0 0 gpio2_out[1]
port 178 nsew signal output
flabel metal3 s 543200 322328 544400 322448 0 FreeSans 480 0 0 0 gpio2_out[2]
port 179 nsew signal output
flabel metal3 s 543200 336200 544400 336320 0 FreeSans 480 0 0 0 gpio2_out[3]
port 180 nsew signal output
flabel metal3 s 543200 410184 544400 410304 0 FreeSans 480 0 0 0 gpio2_out[4]
port 181 nsew signal output
flabel metal3 s 543200 424056 544400 424176 0 FreeSans 480 0 0 0 gpio2_out[5]
port 182 nsew signal output
flabel metal3 s 543200 437928 544400 438048 0 FreeSans 480 0 0 0 gpio2_out[6]
port 183 nsew signal output
flabel metal3 s 543200 451800 544400 451920 0 FreeSans 480 0 0 0 gpio2_out[7]
port 184 nsew signal output
flabel metal4 s 350377 459700 350505 460000 0 FreeSans 960 90 0 0 gpio3_0_analog
port 185 nsew signal bidirectional
flabel metal4 s 349865 459700 349993 460000 0 FreeSans 960 90 0 0 gpio3_1_analog
port 186 nsew signal bidirectional
flabel metal4 s 349353 459700 349481 460000 0 FreeSans 960 90 0 0 gpio3_2_analog
port 187 nsew signal bidirectional
flabel metal4 s 348841 459700 348969 460000 0 FreeSans 960 90 0 0 gpio3_3_analog
port 188 nsew signal bidirectional
flabel metal4 s 348329 459700 348457 460000 0 FreeSans 960 90 0 0 gpio3_4_analog
port 189 nsew signal bidirectional
flabel metal4 s 347817 459700 347945 460000 0 FreeSans 960 90 0 0 gpio3_5_analog
port 190 nsew signal bidirectional
flabel metal4 s 347305 459700 347433 460000 0 FreeSans 960 90 0 0 gpio3_6_analog
port 191 nsew signal bidirectional
flabel metal4 s 346793 459700 346921 460000 0 FreeSans 960 90 0 0 gpio3_7_analog
port 192 nsew signal bidirectional
flabel metal2 s 531410 459200 531466 460400 0 FreeSans 224 90 0 0 gpio3_in[0]
port 193 nsew signal input
flabel metal2 s 525890 459200 525946 460400 0 FreeSans 224 90 0 0 gpio3_in[1]
port 194 nsew signal input
flabel metal2 s 520370 459200 520426 460400 0 FreeSans 224 90 0 0 gpio3_in[2]
port 195 nsew signal input
flabel metal2 s 514850 459200 514906 460400 0 FreeSans 224 90 0 0 gpio3_in[3]
port 196 nsew signal input
flabel metal2 s 509330 459200 509386 460400 0 FreeSans 224 90 0 0 gpio3_in[4]
port 197 nsew signal input
flabel metal2 s 503810 459200 503866 460400 0 FreeSans 224 90 0 0 gpio3_in[5]
port 198 nsew signal input
flabel metal2 s 498290 459200 498346 460400 0 FreeSans 224 90 0 0 gpio3_in[6]
port 199 nsew signal input
flabel metal2 s 492770 459200 492826 460400 0 FreeSans 224 90 0 0 gpio3_in[7]
port 200 nsew signal input
flabel metal2 s 527730 459200 527786 460400 0 FreeSans 224 90 0 0 gpio3_oeb[0]
port 201 nsew signal output
flabel metal2 s 522210 459200 522266 460400 0 FreeSans 224 90 0 0 gpio3_oeb[1]
port 202 nsew signal output
flabel metal2 s 516690 459200 516746 460400 0 FreeSans 224 90 0 0 gpio3_oeb[2]
port 203 nsew signal output
flabel metal2 s 511170 459200 511226 460400 0 FreeSans 224 90 0 0 gpio3_oeb[3]
port 204 nsew signal output
flabel metal2 s 505650 459200 505706 460400 0 FreeSans 224 90 0 0 gpio3_oeb[4]
port 205 nsew signal output
flabel metal2 s 500130 459200 500186 460400 0 FreeSans 224 90 0 0 gpio3_oeb[5]
port 206 nsew signal output
flabel metal2 s 494610 459200 494666 460400 0 FreeSans 224 90 0 0 gpio3_oeb[6]
port 207 nsew signal output
flabel metal2 s 489090 459200 489146 460400 0 FreeSans 224 90 0 0 gpio3_oeb[7]
port 208 nsew signal output
flabel metal2 s 529570 459200 529626 460400 0 FreeSans 224 90 0 0 gpio3_out[0]
port 209 nsew signal output
flabel metal2 s 524050 459200 524106 460400 0 FreeSans 224 90 0 0 gpio3_out[1]
port 210 nsew signal output
flabel metal2 s 518530 459200 518586 460400 0 FreeSans 224 90 0 0 gpio3_out[2]
port 211 nsew signal output
flabel metal2 s 513010 459200 513066 460400 0 FreeSans 224 90 0 0 gpio3_out[3]
port 212 nsew signal output
flabel metal2 s 507490 459200 507546 460400 0 FreeSans 224 90 0 0 gpio3_out[4]
port 213 nsew signal output
flabel metal2 s 501970 459200 502026 460400 0 FreeSans 224 90 0 0 gpio3_out[5]
port 214 nsew signal output
flabel metal2 s 496450 459200 496506 460400 0 FreeSans 224 90 0 0 gpio3_out[6]
port 215 nsew signal output
flabel metal2 s 490930 459200 490986 460400 0 FreeSans 224 90 0 0 gpio3_out[7]
port 216 nsew signal output
flabel metal4 s 346281 459700 346409 460000 0 FreeSans 960 90 0 0 gpio4_0_analog
port 217 nsew signal bidirectional
flabel metal4 s 345769 459700 345897 460000 0 FreeSans 960 90 0 0 gpio4_1_analog
port 218 nsew signal bidirectional
flabel metal4 s 345257 459700 345385 460000 0 FreeSans 960 90 0 0 gpio4_2_analog
port 219 nsew signal bidirectional
flabel metal4 s 344745 459700 344873 460000 0 FreeSans 960 90 0 0 gpio4_3_analog
port 220 nsew signal bidirectional
flabel metal4 s 344233 459700 344361 460000 0 FreeSans 960 90 0 0 gpio4_4_analog
port 221 nsew signal bidirectional
flabel metal4 s 343721 459700 343849 460000 0 FreeSans 960 90 0 0 gpio4_5_analog
port 222 nsew signal bidirectional
flabel metal4 s 343209 459700 343337 460000 0 FreeSans 960 90 0 0 gpio4_6_analog
port 223 nsew signal bidirectional
flabel metal4 s 342697 459700 342825 460000 0 FreeSans 960 90 0 0 gpio4_7_analog
port 224 nsew signal bidirectional
flabel metal2 s 54850 459200 54906 460400 0 FreeSans 224 90 0 0 gpio4_in[0]
port 225 nsew signal input
flabel metal2 s 49330 459200 49386 460400 0 FreeSans 224 90 0 0 gpio4_in[1]
port 226 nsew signal input
flabel metal2 s 43810 459200 43866 460400 0 FreeSans 224 90 0 0 gpio4_in[2]
port 227 nsew signal input
flabel metal2 s 38290 459200 38346 460400 0 FreeSans 224 90 0 0 gpio4_in[3]
port 228 nsew signal input
flabel metal2 s 32770 459200 32826 460400 0 FreeSans 224 90 0 0 gpio4_in[4]
port 229 nsew signal input
flabel metal2 s 27250 459200 27306 460400 0 FreeSans 224 90 0 0 gpio4_in[5]
port 230 nsew signal input
flabel metal2 s 21730 459200 21786 460400 0 FreeSans 224 90 0 0 gpio4_in[6]
port 231 nsew signal input
flabel metal2 s 16210 459200 16266 460400 0 FreeSans 224 90 0 0 gpio4_in[7]
port 232 nsew signal input
flabel metal2 s 51170 459200 51226 460400 0 FreeSans 224 90 0 0 gpio4_oeb[0]
port 233 nsew signal output
flabel metal2 s 45650 459200 45706 460400 0 FreeSans 224 90 0 0 gpio4_oeb[1]
port 234 nsew signal output
flabel metal2 s 40130 459200 40186 460400 0 FreeSans 224 90 0 0 gpio4_oeb[2]
port 235 nsew signal output
flabel metal2 s 34610 459200 34666 460400 0 FreeSans 224 90 0 0 gpio4_oeb[3]
port 236 nsew signal output
flabel metal2 s 29090 459200 29146 460400 0 FreeSans 224 90 0 0 gpio4_oeb[4]
port 237 nsew signal output
flabel metal2 s 23570 459200 23626 460400 0 FreeSans 224 90 0 0 gpio4_oeb[5]
port 238 nsew signal output
flabel metal2 s 18050 459200 18106 460400 0 FreeSans 224 90 0 0 gpio4_oeb[6]
port 239 nsew signal output
flabel metal2 s 12530 459200 12586 460400 0 FreeSans 224 90 0 0 gpio4_oeb[7]
port 240 nsew signal output
flabel metal2 s 53010 459200 53066 460400 0 FreeSans 224 90 0 0 gpio4_out[0]
port 241 nsew signal output
flabel metal2 s 47490 459200 47546 460400 0 FreeSans 224 90 0 0 gpio4_out[1]
port 242 nsew signal output
flabel metal2 s 41970 459200 42026 460400 0 FreeSans 224 90 0 0 gpio4_out[2]
port 243 nsew signal output
flabel metal2 s 36450 459200 36506 460400 0 FreeSans 224 90 0 0 gpio4_out[3]
port 244 nsew signal output
flabel metal2 s 30930 459200 30986 460400 0 FreeSans 224 90 0 0 gpio4_out[4]
port 245 nsew signal output
flabel metal2 s 25410 459200 25466 460400 0 FreeSans 224 90 0 0 gpio4_out[5]
port 246 nsew signal output
flabel metal2 s 19890 459200 19946 460400 0 FreeSans 224 90 0 0 gpio4_out[6]
port 247 nsew signal output
flabel metal2 s 14370 459200 14426 460400 0 FreeSans 224 90 0 0 gpio4_out[7]
port 248 nsew signal output
flabel metal3 s -400 456824 800 456944 0 FreeSans 480 0 0 0 gpio5_in[0]
port 249 nsew signal input
flabel metal3 s -400 442952 800 443072 0 FreeSans 480 0 0 0 gpio5_in[1]
port 250 nsew signal input
flabel metal3 s -400 429080 800 429200 0 FreeSans 480 0 0 0 gpio5_in[2]
port 251 nsew signal input
flabel metal3 s -400 415208 800 415328 0 FreeSans 480 0 0 0 gpio5_in[3]
port 252 nsew signal input
flabel metal3 s -400 340824 800 340944 0 FreeSans 480 0 0 0 gpio5_in[4]
port 253 nsew signal input
flabel metal3 s -400 326952 800 327072 0 FreeSans 480 0 0 0 gpio5_in[5]
port 254 nsew signal input
flabel metal3 s -400 313080 800 313200 0 FreeSans 480 0 0 0 gpio5_in[6]
port 255 nsew signal input
flabel metal3 s -400 299208 800 299328 0 FreeSans 480 0 0 0 gpio5_in[7]
port 256 nsew signal input
flabel metal3 s -400 447576 800 447696 0 FreeSans 480 0 0 0 gpio5_oeb[0]
port 257 nsew signal output
flabel metal3 s -400 433704 800 433824 0 FreeSans 480 0 0 0 gpio5_oeb[1]
port 258 nsew signal output
flabel metal3 s -400 419832 800 419952 0 FreeSans 480 0 0 0 gpio5_oeb[2]
port 259 nsew signal output
flabel metal3 s -400 405960 800 406080 0 FreeSans 480 0 0 0 gpio5_oeb[3]
port 260 nsew signal output
flabel metal3 s -400 331576 800 331696 0 FreeSans 480 0 0 0 gpio5_oeb[4]
port 261 nsew signal output
flabel metal3 s -400 317704 800 317824 0 FreeSans 480 0 0 0 gpio5_oeb[5]
port 262 nsew signal output
flabel metal3 s -400 303832 800 303952 0 FreeSans 480 0 0 0 gpio5_oeb[6]
port 263 nsew signal output
flabel metal3 s -400 289960 800 290080 0 FreeSans 480 0 0 0 gpio5_oeb[7]
port 264 nsew signal output
flabel metal3 s -400 452200 800 452320 0 FreeSans 480 0 0 0 gpio5_out[0]
port 265 nsew signal output
flabel metal3 s -400 438328 800 438448 0 FreeSans 480 0 0 0 gpio5_out[1]
port 266 nsew signal output
flabel metal3 s -400 424456 800 424576 0 FreeSans 480 0 0 0 gpio5_out[2]
port 267 nsew signal output
flabel metal3 s -400 410584 800 410704 0 FreeSans 480 0 0 0 gpio5_out[3]
port 268 nsew signal output
flabel metal3 s -400 336200 800 336320 0 FreeSans 480 0 0 0 gpio5_out[4]
port 269 nsew signal output
flabel metal3 s -400 322328 800 322448 0 FreeSans 480 0 0 0 gpio5_out[5]
port 270 nsew signal output
flabel metal3 s -400 308456 800 308576 0 FreeSans 480 0 0 0 gpio5_out[6]
port 271 nsew signal output
flabel metal3 s -400 294584 800 294704 0 FreeSans 480 0 0 0 gpio5_out[7]
port 272 nsew signal output
flabel metal3 s -400 285336 800 285456 0 FreeSans 480 0 0 0 gpio6_in[0]
port 273 nsew signal input
flabel metal3 s -400 271464 800 271584 0 FreeSans 480 0 0 0 gpio6_in[1]
port 274 nsew signal input
flabel metal3 s -400 257592 800 257712 0 FreeSans 480 0 0 0 gpio6_in[2]
port 275 nsew signal input
flabel metal3 s -400 243720 800 243840 0 FreeSans 480 0 0 0 gpio6_in[3]
port 276 nsew signal input
flabel metal3 s -400 229848 800 229968 0 FreeSans 480 0 0 0 gpio6_in[4]
port 277 nsew signal input
flabel metal3 s -400 215976 800 216096 0 FreeSans 480 0 0 0 gpio6_in[5]
port 278 nsew signal input
flabel metal3 s -400 202104 800 202224 0 FreeSans 480 0 0 0 gpio6_in[6]
port 279 nsew signal input
flabel metal3 s -400 188232 800 188352 0 FreeSans 480 0 0 0 gpio6_in[7]
port 280 nsew signal input
flabel metal3 s -400 276088 800 276208 0 FreeSans 480 0 0 0 gpio6_oeb[0]
port 281 nsew signal output
flabel metal3 s -400 262216 800 262336 0 FreeSans 480 0 0 0 gpio6_oeb[1]
port 282 nsew signal output
flabel metal3 s -400 248344 800 248464 0 FreeSans 480 0 0 0 gpio6_oeb[2]
port 283 nsew signal output
flabel metal3 s -400 234472 800 234592 0 FreeSans 480 0 0 0 gpio6_oeb[3]
port 284 nsew signal output
flabel metal3 s -400 220600 800 220720 0 FreeSans 480 0 0 0 gpio6_oeb[4]
port 285 nsew signal output
flabel metal3 s -400 206728 800 206848 0 FreeSans 480 0 0 0 gpio6_oeb[5]
port 286 nsew signal output
flabel metal3 s -400 192856 800 192976 0 FreeSans 480 0 0 0 gpio6_oeb[6]
port 287 nsew signal output
flabel metal3 s -400 178984 800 179104 0 FreeSans 480 0 0 0 gpio6_oeb[7]
port 288 nsew signal output
flabel metal3 s -400 280712 800 280832 0 FreeSans 480 0 0 0 gpio6_out[0]
port 289 nsew signal output
flabel metal3 s -400 266840 800 266960 0 FreeSans 480 0 0 0 gpio6_out[1]
port 290 nsew signal output
flabel metal3 s -400 252968 800 253088 0 FreeSans 480 0 0 0 gpio6_out[2]
port 291 nsew signal output
flabel metal3 s -400 239096 800 239216 0 FreeSans 480 0 0 0 gpio6_out[3]
port 292 nsew signal output
flabel metal3 s -400 225224 800 225344 0 FreeSans 480 0 0 0 gpio6_out[4]
port 293 nsew signal output
flabel metal3 s -400 211352 800 211472 0 FreeSans 480 0 0 0 gpio6_out[5]
port 294 nsew signal output
flabel metal3 s -400 197480 800 197600 0 FreeSans 480 0 0 0 gpio6_out[6]
port 295 nsew signal output
flabel metal3 s -400 183608 800 183728 0 FreeSans 480 0 0 0 gpio6_out[7]
port 296 nsew signal output
flabel metal3 s -400 174064 800 174184 0 FreeSans 480 0 0 0 gpio7_in[0]
port 297 nsew signal input
flabel metal3 s -400 160192 800 160312 0 FreeSans 480 0 0 0 gpio7_in[1]
port 298 nsew signal input
flabel metal3 s -400 146320 800 146440 0 FreeSans 480 0 0 0 gpio7_in[2]
port 299 nsew signal input
flabel metal3 s -400 114248 800 114368 0 FreeSans 480 0 0 0 gpio7_in[3]
port 300 nsew signal input
flabel metal3 s -400 100376 800 100496 0 FreeSans 480 0 0 0 gpio7_in[4]
port 301 nsew signal input
flabel metal3 s -400 86504 800 86624 0 FreeSans 480 0 0 0 gpio7_in[5]
port 302 nsew signal input
flabel metal3 s -400 72632 800 72752 0 FreeSans 480 0 0 0 gpio7_in[6]
port 303 nsew signal input
flabel metal3 s -400 58760 800 58880 0 FreeSans 480 0 0 0 gpio7_in[7]
port 304 nsew signal input
flabel metal3 s -400 164816 800 164936 0 FreeSans 480 0 0 0 gpio7_oeb[0]
port 305 nsew signal output
flabel metal3 s -400 150944 800 151064 0 FreeSans 480 0 0 0 gpio7_oeb[1]
port 306 nsew signal output
flabel metal3 s -400 118872 800 118992 0 FreeSans 480 0 0 0 gpio7_oeb[2]
port 307 nsew signal output
flabel metal3 s -400 105000 800 105120 0 FreeSans 480 0 0 0 gpio7_oeb[3]
port 308 nsew signal output
flabel metal3 s -400 91128 800 91248 0 FreeSans 480 0 0 0 gpio7_oeb[4]
port 309 nsew signal output
flabel metal3 s -400 77256 800 77376 0 FreeSans 480 0 0 0 gpio7_oeb[5]
port 310 nsew signal output
flabel metal3 s -400 63384 800 63504 0 FreeSans 480 0 0 0 gpio7_oeb[6]
port 311 nsew signal output
flabel metal3 s -400 49512 800 49632 0 FreeSans 480 0 0 0 gpio7_oeb[7]
port 312 nsew signal output
flabel metal3 s -400 169440 800 169560 0 FreeSans 480 0 0 0 gpio7_out[0]
port 313 nsew signal output
flabel metal3 s -400 155568 800 155688 0 FreeSans 480 0 0 0 gpio7_out[1]
port 314 nsew signal output
flabel metal3 s -400 123496 800 123616 0 FreeSans 480 0 0 0 gpio7_out[2]
port 315 nsew signal output
flabel metal3 s -400 109624 800 109744 0 FreeSans 480 0 0 0 gpio7_out[3]
port 316 nsew signal output
flabel metal3 s -400 95752 800 95872 0 FreeSans 480 0 0 0 gpio7_out[4]
port 317 nsew signal output
flabel metal3 s -400 81880 800 82000 0 FreeSans 480 0 0 0 gpio7_out[5]
port 318 nsew signal output
flabel metal3 s -400 68008 800 68128 0 FreeSans 480 0 0 0 gpio7_out[6]
port 319 nsew signal output
flabel metal3 s -400 54136 800 54256 0 FreeSans 480 0 0 0 gpio7_out[7]
port 320 nsew signal output
flabel metal4 s 339113 459700 339241 460000 0 FreeSans 960 90 0 0 ibias100
port 321 nsew signal bidirectional
flabel metal4 s 338601 459700 338729 460000 0 FreeSans 960 90 0 0 ibias50
port 322 nsew signal bidirectional
flabel metal4 s 335017 459700 335145 460000 0 FreeSans 960 90 0 0 left_vref
port 323 nsew signal bidirectional
flabel metal4 s 335529 459700 335657 460000 0 FreeSans 960 90 0 0 right_vref
port 324 nsew signal bidirectional
flabel metal2 s 489194 -400 489250 800 0 FreeSans 224 90 0 0 sio_in[0]
port 325 nsew signal input
flabel metal2 s 493886 -400 493942 800 0 FreeSans 224 90 0 0 sio_in[1]
port 326 nsew signal input
flabel metal2 s 492322 -400 492378 800 0 FreeSans 224 90 0 0 sio_oeb[0]
port 327 nsew signal output
flabel metal2 s 497014 -400 497070 800 0 FreeSans 224 90 0 0 sio_oeb[1]
port 328 nsew signal output
flabel metal2 s 490758 -400 490814 800 0 FreeSans 224 90 0 0 sio_out[0]
port 329 nsew signal output
flabel metal2 s 495450 -400 495506 800 0 FreeSans 224 90 0 0 sio_out[1]
port 330 nsew signal output
flabel metal4 s 336041 459700 336169 460000 0 FreeSans 960 90 0 0 tempsense
port 331 nsew signal bidirectional
flabel metal4 s 341673 459700 341801 460000 0 FreeSans 960 90 0 0 ulpcomp_n
port 332 nsew signal bidirectional
flabel metal4 s 342185 459700 342313 460000 0 FreeSans 960 90 0 0 ulpcomp_p
port 333 nsew signal bidirectional
flabel metal2 s 214278 -400 214334 800 0 FreeSans 224 90 0 0 user_irq[0]
port 334 nsew signal output
flabel metal2 s 229918 -400 229974 800 0 FreeSans 224 90 0 0 user_irq[10]
port 335 nsew signal output
flabel metal2 s 231482 -400 231538 800 0 FreeSans 224 90 0 0 user_irq[11]
port 336 nsew signal output
flabel metal2 s 233046 -400 233102 800 0 FreeSans 224 90 0 0 user_irq[12]
port 337 nsew signal output
flabel metal2 s 234610 -400 234666 800 0 FreeSans 224 90 0 0 user_irq[13]
port 338 nsew signal output
flabel metal2 s 236174 -400 236230 800 0 FreeSans 224 90 0 0 user_irq[14]
port 339 nsew signal output
flabel metal2 s 237738 -400 237794 800 0 FreeSans 224 90 0 0 user_irq[15]
port 340 nsew signal output
flabel metal2 s 215842 -400 215898 800 0 FreeSans 224 90 0 0 user_irq[1]
port 341 nsew signal output
flabel metal2 s 217406 -400 217462 800 0 FreeSans 224 90 0 0 user_irq[2]
port 342 nsew signal output
flabel metal2 s 218970 -400 219026 800 0 FreeSans 224 90 0 0 user_irq[3]
port 343 nsew signal output
flabel metal2 s 220534 -400 220590 800 0 FreeSans 224 90 0 0 user_irq[4]
port 344 nsew signal output
flabel metal2 s 222098 -400 222154 800 0 FreeSans 224 90 0 0 user_irq[5]
port 345 nsew signal output
flabel metal2 s 223662 -400 223718 800 0 FreeSans 224 90 0 0 user_irq[6]
port 346 nsew signal output
flabel metal2 s 225226 -400 225282 800 0 FreeSans 224 90 0 0 user_irq[7]
port 347 nsew signal output
flabel metal2 s 226790 -400 226846 800 0 FreeSans 224 90 0 0 user_irq[8]
port 348 nsew signal output
flabel metal2 s 228354 -400 228410 800 0 FreeSans 224 90 0 0 user_irq[9]
port 349 nsew signal output
flabel metal4 s 338089 459700 338217 460000 0 FreeSans 960 90 0 0 vbgsc
port 350 nsew signal bidirectional
flabel metal4 s 337577 459700 337705 460000 0 FreeSans 960 90 0 0 vbgtc
port 351 nsew signal bidirectional
flabel metal4 s -1596 -1444 -976 461124 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -1596 -1444 545592 -824 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -1596 460504 545592 461124 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 544972 -1444 545592 461124 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 4714 880 5334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 22714 880 23334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 40714 880 41334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 58714 -4324 59334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 76714 -4324 77334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 94714 -4324 95334 19988 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 94714 59724 95334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 112714 -4324 113334 17955 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 112714 58629 113334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 130714 -4324 131334 17955 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 130714 58629 131334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 148714 -4324 149334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 166714 -4324 167334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 184714 -4324 185334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 202714 -4324 203334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 220714 -4324 221334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 238714 -4324 239334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 256714 -4324 257334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 274714 -4324 275334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 292714 -4324 293334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 310714 -4324 311334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 328714 -4324 329334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 346714 -4324 347334 458520 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 364714 -4324 365334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 382714 -4324 383334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 400714 -4324 401334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 418714 -4324 419334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 436714 -4324 437334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 454714 -4324 455334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 472714 -4324 473334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 490714 -4324 491334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 508714 880 509334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s 526714 880 527334 464004 0 FreeSans 3840 90 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 4866 548472 5486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 22866 101780 23486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 40866 548472 41486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 58866 548472 59486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 76866 548472 77486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 94866 548472 95486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 112866 548472 113486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 130866 548472 131486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 148866 548472 149486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 166866 548472 167486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 184866 548472 185486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 202866 548472 203486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 220866 548472 221486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 238866 548472 239486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 256866 548472 257486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 274866 548472 275486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 292866 548472 293486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 310866 548472 311486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 328866 548472 329486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 346866 548472 347486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 364866 548472 365486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 382866 548472 383486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 400866 548472 401486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 418866 548472 419486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 436866 548472 437486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s -4476 454866 548472 455486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal5 s 133972 22866 548472 23486 0 FreeSans 2560 0 0 0 vccd1
port 352 nsew power bidirectional
flabel metal4 s -3516 -3364 -2896 463044 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -3516 -3364 547512 -2744 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -3516 462424 547512 463044 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 546892 -3364 547512 463044 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 12154 880 12774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 30154 880 30774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 48154 -4324 48774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 66154 -4324 66774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 84154 -4324 84774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 102154 -4324 102774 17955 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 102154 58629 102774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 120154 -4324 120774 17955 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 120154 58629 120774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 138154 -4324 138774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 156154 -4324 156774 19988 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 156154 59724 156774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 174154 -4324 174774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 192154 -4324 192774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 210154 -4324 210774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 228154 -4324 228774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 246154 -4324 246774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 264154 -4324 264774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 282154 -4324 282774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 300154 -4324 300774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 318154 -4324 318774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 336154 -4324 336774 458520 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 354154 -4324 354774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 372154 -4324 372774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 390154 -4324 390774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 408154 -4324 408774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 426154 -4324 426774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 444154 -4324 444774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 462154 -4324 462774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 480154 -4324 480774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 498154 -4324 498774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 516154 880 516774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal4 s 534154 880 534774 464004 0 FreeSans 3840 90 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 12306 548472 12926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 30306 101780 30926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 48306 548472 48926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 66306 548472 66926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 84306 548472 84926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 102306 548472 102926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 120306 548472 120926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 138306 548472 138926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 156306 548472 156926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 174306 548472 174926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 192306 548472 192926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 210306 548472 210926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 228306 548472 228926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 246306 548472 246926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 264306 548472 264926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 282306 548472 282926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 300306 548472 300926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 318306 548472 318926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 336306 548472 336926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 354306 548472 354926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 372306 548472 372926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 390306 548472 390926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 408306 548472 408926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 426306 548472 426926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s -4476 444306 548472 444926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal5 s 133972 30306 548472 30926 0 FreeSans 2560 0 0 0 vccd2
port 353 nsew power bidirectional
flabel metal3 s 543356 344572 544000 349352 0 FreeSans 3840 90 0 0 vdda1
port 354 nsew power input
flabel metal3 s 543356 354551 544000 359331 0 FreeSans 3840 90 0 0 vdda1
port 355 nsew power input
flabel metal4 s 500302 0 505082 638 0 FreeSans 3840 0 0 0 vdda1
port 356 nsew power input
flabel metal4 s 510281 0 515061 638 0 FreeSans 3840 0 0 0 vdda1
port 357 nsew power input
flabel metal3 s 0 357308 644 362088 0 FreeSans 3840 90 0 0 vdda2
port 358 nsew power input
flabel metal3 s 0 347329 644 352109 0 FreeSans 3840 90 0 0 vdda2
port 359 nsew power input
flabel metal4 s 28939 0 33719 638 0 FreeSans 3840 0 0 0 vdda2
port 360 nsew power input
flabel metal4 s 38918 0 43698 638 0 FreeSans 3840 0 0 0 vdda2
port 361 nsew power input
flabel metal4 s 334505 459700 334633 460000 0 FreeSans 960 90 0 0 vinref
port 362 nsew signal bidirectional
flabel metal4 s 333993 459700 334121 460000 0 FreeSans 960 90 0 0 voutref
port 363 nsew signal bidirectional
flabel metal3 s 543356 378550 544000 383330 0 FreeSans 3840 90 0 0 vssa1
port 364 nsew ground input
flabel metal3 s 543356 368571 544000 373351 0 FreeSans 3840 90 0 0 vssa1
port 365 nsew ground input
flabel metal4 s 534281 0 539061 638 0 FreeSans 3840 0 0 0 vssa1
port 366 nsew ground input
flabel metal4 s 524302 0 529082 638 0 FreeSans 3840 0 0 0 vssa1
port 367 nsew ground input
flabel metal3 s 0 380308 644 385088 0 FreeSans 3840 90 0 0 vssa2
port 368 nsew ground input
flabel metal3 s 0 370329 644 375109 0 FreeSans 3840 90 0 0 vssa2
port 369 nsew ground input
flabel metal4 s 14918 0 19698 638 0 FreeSans 3840 0 0 0 vssa2
port 370 nsew ground input
flabel metal4 s 4939 0 9719 638 0 FreeSans 3840 0 0 0 vssa2
port 371 nsew ground input
flabel metal4 s -2556 -2404 -1936 462084 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -2556 -2404 546552 -1784 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -2556 461464 546552 462084 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 545932 -2404 546552 462084 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 8434 880 9054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 26434 880 27054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 44434 880 45054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 62434 -4324 63054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 80434 -4324 81054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 98434 -4324 99054 17955 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 98434 58629 99054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 116434 -4324 117054 17955 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 116434 58629 117054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 134434 -4324 135054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 152434 -4324 153054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 170434 -4324 171054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 188434 -4324 189054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 206434 -4324 207054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 224434 -4324 225054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 242434 -4324 243054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 260434 -4324 261054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 278434 -4324 279054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 296434 -4324 297054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 314434 -4324 315054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 332434 -4324 333054 458520 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 350434 -4324 351054 458520 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 368434 -4324 369054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 386434 -4324 387054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 404434 -4324 405054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 422434 -4324 423054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 440434 -4324 441054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 458434 -4324 459054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 476434 -4324 477054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 494434 -4324 495054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 512434 880 513054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s 530434 880 531054 464004 0 FreeSans 3840 90 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 8586 548472 9206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 26586 101780 27206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 44586 548472 45206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 62586 548472 63206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 80586 548472 81206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 98586 548472 99206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 116586 548472 117206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 134586 548472 135206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 152586 548472 153206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 170586 548472 171206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 188586 548472 189206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 206586 548472 207206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 224586 548472 225206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 242586 548472 243206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 260586 548472 261206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 278586 548472 279206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 296586 548472 297206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 314586 548472 315206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 332586 548472 333206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 350586 548472 351206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 368586 548472 369206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 386586 548472 387206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 404586 548472 405206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 422586 548472 423206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s -4476 440586 548472 441206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal5 s 133972 26586 548472 27206 0 FreeSans 2560 0 0 0 vssd1
port 372 nsew ground bidirectional
flabel metal4 s -4476 -4324 -3856 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 -4324 548472 -3704 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 463384 548472 464004 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 547852 -4324 548472 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 15874 880 16494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 33874 880 34494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 51874 -4324 52494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 69874 -4324 70494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 87874 -4324 88494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 105874 -4324 106494 17955 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 105874 58629 106494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 123874 -4324 124494 17955 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 123874 58629 124494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 141874 -4324 142494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 159874 -4324 160494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 177874 -4324 178494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 195874 -4324 196494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 213874 -4324 214494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 231874 -4324 232494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 249874 -4324 250494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 267874 -4324 268494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 285874 -4324 286494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 303874 -4324 304494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 321874 -4324 322494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 339874 -4324 340494 458520 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 357874 -4324 358494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 375874 -4324 376494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 393874 -4324 394494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 411874 -4324 412494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 429874 -4324 430494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 447874 -4324 448494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 465874 -4324 466494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 483874 -4324 484494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 501874 880 502494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 519874 880 520494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal4 s 537874 880 538494 464004 0 FreeSans 3840 90 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 16026 548472 16646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 34026 548472 34646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 52026 548472 52646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 70026 548472 70646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 88026 548472 88646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 106026 548472 106646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 124026 548472 124646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 142026 548472 142646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 160026 548472 160646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 178026 548472 178646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 196026 548472 196646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 214026 548472 214646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 232026 548472 232646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 250026 548472 250646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 268026 548472 268646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 286026 548472 286646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 304026 548472 304646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 322026 548472 322646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 340026 548472 340646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 358026 548472 358646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 376026 548472 376646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 394026 548472 394646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 412026 548472 412646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 430026 548472 430646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
flabel metal5 s -4476 448026 548472 448646 0 FreeSans 2560 0 0 0 vssd2
port 373 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 544000 460000
<< end >>
